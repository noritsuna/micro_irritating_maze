magic
tech gf180mcuD
magscale 1 10
timestamp 1698784607
<< metal2 >>
rect 11032 595672 11256 597000
rect 33096 595672 33320 597000
rect 55160 595672 55384 597000
rect 11004 595560 11256 595672
rect 33068 595560 33320 595672
rect 55132 595560 55384 595672
rect 77224 595560 77448 597000
rect 99288 595672 99512 597000
rect 121352 595672 121576 597000
rect 143416 595672 143640 597000
rect 165480 595672 165704 597000
rect 187544 595672 187768 597000
rect 209608 595672 209832 597000
rect 231672 595672 231896 597000
rect 253736 595672 253960 597000
rect 275800 595672 276024 597000
rect 297864 595672 298088 597000
rect 319928 595672 320152 597000
rect 341992 595672 342216 597000
rect 364056 595672 364280 597000
rect 386120 595672 386344 597000
rect 99260 595560 99512 595672
rect 121324 595560 121576 595672
rect 143388 595560 143640 595672
rect 165452 595560 165704 595672
rect 187516 595560 187768 595672
rect 209580 595560 209832 595672
rect 231644 595560 231896 595672
rect 253708 595560 253960 595672
rect 275772 595560 276024 595672
rect 297836 595560 298088 595672
rect 319900 595560 320152 595672
rect 341964 595560 342216 595672
rect 364028 595560 364280 595672
rect 386092 595560 386344 595672
rect 408184 595560 408408 597000
rect 430248 595672 430472 597000
rect 452312 595672 452536 597000
rect 474376 595672 474600 597000
rect 496440 595672 496664 597000
rect 518504 595672 518728 597000
rect 540568 595672 540792 597000
rect 562632 595672 562856 597000
rect 584696 595672 584920 597000
rect 430220 595560 430472 595672
rect 452284 595560 452536 595672
rect 474348 595560 474600 595672
rect 496412 595560 496664 595672
rect 518476 595560 518728 595672
rect 540540 595560 540792 595672
rect 562604 595560 562856 595672
rect 584668 595560 584920 595672
rect 9996 590548 10052 590558
rect 1596 583828 1652 583838
rect 1484 86548 1540 86558
rect 1484 36708 1540 86492
rect 1596 38500 1652 583772
rect 8316 91588 8372 91598
rect 8204 89908 8260 89918
rect 1596 38434 1652 38444
rect 3276 86660 3332 86670
rect 1484 36642 1540 36652
rect 3276 34020 3332 86604
rect 4956 84980 5012 84990
rect 4844 83188 4900 83198
rect 4844 42980 4900 83132
rect 4844 42914 4900 42924
rect 4956 37604 5012 84924
rect 7980 84868 8036 84878
rect 4956 37538 5012 37548
rect 6636 73220 6692 73230
rect 3276 33954 3332 33964
rect 6636 29540 6692 73164
rect 7980 49252 8036 84812
rect 7980 49186 8036 49196
rect 8092 74900 8148 74910
rect 8092 31332 8148 74844
rect 8204 43876 8260 89852
rect 8204 43810 8260 43820
rect 8316 41188 8372 91532
rect 9772 76468 9828 76478
rect 9660 73444 9716 73454
rect 9660 65604 9716 73388
rect 9772 69636 9828 76412
rect 9772 69570 9828 69580
rect 9884 73332 9940 73342
rect 9660 65538 9716 65548
rect 9884 57204 9940 73276
rect 9884 57138 9940 57148
rect 9996 51940 10052 590492
rect 9996 51874 10052 51884
rect 8316 41122 8372 41132
rect 8092 31266 8148 31276
rect 6636 29474 6692 29484
rect 11004 28644 11060 595560
rect 22652 469700 22708 469710
rect 12124 103348 12180 103358
rect 12012 101668 12068 101678
rect 11676 96628 11732 96638
rect 11564 88228 11620 88238
rect 11452 73108 11508 73118
rect 11452 30436 11508 73052
rect 11564 46564 11620 88172
rect 11676 50148 11732 96572
rect 11676 50082 11732 50092
rect 11564 46498 11620 46508
rect 12012 39956 12068 101612
rect 12124 46340 12180 103292
rect 12236 98308 12292 98318
rect 12236 48132 12292 98252
rect 22652 73444 22708 469644
rect 22652 73378 22708 73388
rect 33068 73220 33124 595560
rect 34412 535780 34468 535790
rect 34412 73332 34468 535724
rect 46172 377188 46228 377198
rect 46172 76468 46228 377132
rect 46172 76402 46228 76412
rect 34412 73266 34468 73276
rect 33068 73154 33124 73164
rect 55132 73108 55188 595560
rect 77308 74900 77364 595560
rect 99260 590212 99316 595560
rect 99260 590146 99316 590156
rect 121324 590212 121380 595560
rect 121324 590146 121380 590156
rect 143388 86660 143444 595560
rect 165452 590212 165508 595560
rect 165452 590146 165508 590156
rect 187516 590212 187572 595560
rect 187516 590146 187572 590156
rect 143388 86594 143444 86604
rect 209580 86548 209636 595560
rect 209580 86482 209636 86492
rect 231644 84980 231700 595560
rect 253708 583828 253764 595560
rect 253708 583762 253764 583772
rect 275772 101668 275828 595560
rect 297836 590212 297892 595560
rect 297836 590146 297892 590156
rect 275772 101602 275828 101612
rect 319900 91588 319956 595560
rect 341964 590212 342020 595560
rect 341964 590146 342020 590156
rect 319900 91522 319956 91532
rect 231644 84914 231700 84924
rect 364028 83188 364084 595560
rect 386092 89908 386148 595560
rect 408268 590660 408324 595560
rect 408268 590594 408324 590604
rect 430220 103348 430276 595560
rect 430220 103282 430276 103292
rect 386092 89842 386148 89852
rect 452284 88228 452340 595560
rect 474348 98308 474404 595560
rect 496412 578788 496468 595560
rect 496412 578722 496468 578732
rect 474348 98242 474404 98252
rect 452284 88162 452340 88172
rect 518476 84868 518532 595560
rect 540540 96628 540596 595560
rect 562604 582148 562660 595560
rect 584668 590548 584724 595560
rect 584668 590482 584724 590492
rect 562604 582082 562660 582092
rect 540540 96562 540596 96572
rect 518476 84802 518532 84812
rect 364028 83122 364084 83132
rect 129388 82516 129444 82526
rect 125580 82404 125636 82414
rect 123676 80836 123732 80846
rect 123564 79044 123620 79054
rect 77308 74834 77364 74844
rect 123452 75684 123508 75694
rect 55132 73042 55188 73052
rect 12236 48066 12292 48076
rect 12124 46274 12180 46284
rect 12012 39890 12068 39900
rect 11452 30370 11508 30380
rect 11004 28578 11060 28588
rect 123452 6244 123508 75628
rect 123564 11060 123620 78988
rect 123564 10994 123620 11004
rect 123452 6178 123508 6188
rect 123564 6916 123620 6926
rect 40012 3780 40068 3790
rect 40012 3714 40068 3724
rect 40908 3780 40964 3790
rect 40908 3714 40964 3724
rect 41356 3780 41412 3790
rect 41356 3714 41412 3724
rect 43148 3780 43204 3790
rect 43148 3714 43204 3724
rect 44268 3780 44324 3790
rect 44268 3714 44324 3724
rect 44716 3780 44772 3790
rect 44716 3714 44772 3724
rect 44940 3780 44996 3790
rect 44940 3714 44996 3724
rect 45612 3780 45668 3790
rect 45612 3714 45668 3724
rect 46284 3780 46340 3790
rect 46284 3714 46340 3724
rect 46732 3780 46788 3790
rect 46732 3714 46788 3724
rect 47628 3780 47684 3790
rect 47628 3714 47684 3724
rect 48300 3780 48356 3790
rect 48300 3714 48356 3724
rect 48524 3780 48580 3790
rect 48524 3714 48580 3724
rect 48972 3780 49028 3790
rect 48972 3714 49028 3724
rect 49196 3780 49252 3790
rect 49196 3714 49252 3724
rect 49868 3780 49924 3790
rect 49868 3714 49924 3724
rect 50316 3780 50372 3790
rect 50316 3714 50372 3724
rect 50540 3780 50596 3790
rect 50540 3714 50596 3724
rect 50988 3780 51044 3790
rect 50988 3714 51044 3724
rect 51212 3780 51268 3790
rect 51212 3714 51268 3724
rect 51884 3780 51940 3790
rect 51884 3714 51940 3724
rect 52332 3780 52388 3790
rect 52332 3714 52388 3724
rect 53228 3780 53284 3790
rect 53228 3714 53284 3724
rect 53676 3780 53732 3790
rect 53676 3714 53732 3724
rect 53900 3780 53956 3790
rect 53900 3714 53956 3724
rect 54124 3780 54180 3790
rect 54124 3714 54180 3724
rect 54348 3780 54404 3790
rect 54348 3714 54404 3724
rect 55020 3780 55076 3790
rect 55020 3714 55076 3724
rect 55692 3780 55748 3790
rect 55692 3714 55748 3724
rect 55916 3780 55972 3790
rect 55916 3714 55972 3724
rect 57036 3780 57092 3790
rect 57036 3714 57092 3724
rect 57260 3780 57316 3790
rect 57260 3714 57316 3724
rect 57708 3780 57764 3790
rect 57708 3714 57764 3724
rect 57932 3780 57988 3790
rect 57932 3714 57988 3724
rect 58604 3780 58660 3790
rect 58604 3714 58660 3724
rect 58828 3780 58884 3790
rect 58828 3714 58884 3724
rect 59276 3780 59332 3790
rect 59276 3714 59332 3724
rect 59500 3780 59556 3790
rect 59500 3714 59556 3724
rect 59724 3780 59780 3790
rect 59724 3714 59780 3724
rect 60172 3780 60228 3790
rect 60172 3714 60228 3724
rect 60396 3780 60452 3790
rect 60396 3714 60452 3724
rect 60844 3780 60900 3790
rect 60844 3714 60900 3724
rect 61068 3780 61124 3790
rect 61068 3714 61124 3724
rect 61292 3780 61348 3790
rect 61292 3714 61348 3724
rect 61964 3780 62020 3790
rect 61964 3714 62020 3724
rect 63084 3780 63140 3790
rect 63084 3714 63140 3724
rect 63980 3780 64036 3790
rect 63980 3714 64036 3724
rect 64204 3780 64260 3790
rect 64204 3714 64260 3724
rect 64428 3780 64484 3790
rect 64428 3714 64484 3724
rect 64652 3780 64708 3790
rect 64652 3714 64708 3724
rect 65324 3780 65380 3790
rect 65324 3714 65380 3724
rect 65996 3780 66052 3790
rect 65996 3714 66052 3724
rect 66220 3780 66276 3790
rect 66220 3714 66276 3724
rect 67116 3780 67172 3790
rect 67116 3714 67172 3724
rect 67788 3780 67844 3790
rect 67788 3714 67844 3724
rect 68684 3780 68740 3790
rect 68684 3714 68740 3724
rect 68908 3780 68964 3790
rect 68908 3714 68964 3724
rect 69132 3780 69188 3790
rect 69132 3714 69188 3724
rect 69356 3780 69412 3790
rect 69356 3714 69412 3724
rect 69804 3780 69860 3790
rect 69804 3714 69860 3724
rect 70476 3780 70532 3790
rect 70476 3714 70532 3724
rect 71596 3780 71652 3790
rect 71596 3714 71652 3724
rect 71820 3780 71876 3790
rect 71820 3714 71876 3724
rect 72268 3780 72324 3790
rect 72268 3714 72324 3724
rect 72492 3780 72548 3790
rect 72492 3714 72548 3724
rect 72716 3780 72772 3790
rect 72716 3714 72772 3724
rect 72940 3780 72996 3790
rect 72940 3714 72996 3724
rect 73612 3780 73668 3790
rect 73612 3714 73668 3724
rect 73836 3780 73892 3790
rect 73836 3714 73892 3724
rect 74508 3780 74564 3790
rect 74508 3714 74564 3724
rect 74956 3780 75012 3790
rect 74956 3714 75012 3724
rect 75404 3780 75460 3790
rect 75404 3714 75460 3724
rect 75852 3780 75908 3790
rect 75852 3714 75908 3724
rect 76076 3780 76132 3790
rect 76076 3714 76132 3724
rect 77196 3780 77252 3790
rect 77196 3714 77252 3724
rect 77644 3780 77700 3790
rect 77644 3714 77700 3724
rect 77868 3780 77924 3790
rect 77868 3714 77924 3724
rect 79212 3780 79268 3790
rect 79212 3714 79268 3724
rect 79884 3780 79940 3790
rect 79884 3714 79940 3724
rect 80108 3780 80164 3790
rect 80108 3714 80164 3724
rect 80780 3780 80836 3790
rect 80780 3714 80836 3724
rect 81228 3780 81284 3790
rect 81228 3714 81284 3724
rect 81900 3780 81956 3790
rect 81900 3714 81956 3724
rect 82572 3780 82628 3790
rect 82572 3714 82628 3724
rect 82796 3780 82852 3790
rect 82796 3714 82852 3724
rect 83244 3780 83300 3790
rect 83244 3714 83300 3724
rect 83692 3780 83748 3790
rect 83692 3714 83748 3724
rect 84140 3780 84196 3790
rect 84140 3714 84196 3724
rect 84588 3780 84644 3790
rect 84588 3714 84644 3724
rect 85260 3780 85316 3790
rect 85260 3714 85316 3724
rect 85932 3780 85988 3790
rect 85932 3714 85988 3724
rect 86156 3780 86212 3790
rect 86156 3714 86212 3724
rect 86604 3780 86660 3790
rect 86604 3714 86660 3724
rect 86828 3780 86884 3790
rect 86828 3714 86884 3724
rect 87276 3780 87332 3790
rect 87276 3714 87332 3724
rect 87500 3780 87556 3790
rect 87500 3714 87556 3724
rect 87948 3780 88004 3790
rect 87948 3714 88004 3724
rect 88620 3780 88676 3790
rect 88620 3714 88676 3724
rect 88844 3780 88900 3790
rect 88844 3714 88900 3724
rect 89068 3780 89124 3790
rect 89068 3714 89124 3724
rect 89292 3780 89348 3790
rect 89292 3714 89348 3724
rect 89516 3780 89572 3790
rect 89516 3714 89572 3724
rect 89964 3780 90020 3790
rect 89964 3714 90020 3724
rect 90636 3780 90692 3790
rect 90636 3714 90692 3724
rect 90860 3780 90916 3790
rect 90860 3714 90916 3724
rect 91308 3780 91364 3790
rect 91308 3714 91364 3724
rect 92204 3780 92260 3790
rect 92204 3714 92260 3724
rect 93100 3780 93156 3790
rect 93100 3714 93156 3724
rect 93548 3780 93604 3790
rect 93548 3714 93604 3724
rect 94220 3780 94276 3790
rect 94220 3714 94276 3724
rect 94892 3780 94948 3790
rect 94892 3714 94948 3724
rect 96012 3780 96068 3790
rect 96012 3714 96068 3724
rect 96236 3780 96292 3790
rect 96236 3714 96292 3724
rect 96908 3780 96964 3790
rect 96908 3714 96964 3724
rect 97356 3780 97412 3790
rect 97356 3714 97412 3724
rect 98700 3780 98756 3790
rect 98700 3714 98756 3724
rect 99372 3780 99428 3790
rect 99372 3714 99428 3724
rect 99596 3780 99652 3790
rect 99596 3714 99652 3724
rect 99820 3780 99876 3790
rect 99820 3714 99876 3724
rect 100268 3780 100324 3790
rect 100268 3714 100324 3724
rect 100716 3780 100772 3790
rect 100716 3714 100772 3724
rect 100940 3780 100996 3790
rect 100940 3714 100996 3724
rect 39564 3668 39620 3678
rect 39564 3602 39620 3612
rect 42028 3668 42084 3678
rect 42028 3602 42084 3612
rect 42700 3668 42756 3678
rect 42700 3602 42756 3612
rect 62860 3668 62916 3678
rect 62860 3602 62916 3612
rect 63532 3668 63588 3678
rect 63532 3602 63588 3612
rect 64876 3668 64932 3678
rect 64876 3602 64932 3612
rect 65100 3668 65156 3678
rect 65100 3602 65156 3612
rect 65548 3668 65604 3678
rect 65548 3602 65604 3612
rect 66668 3668 66724 3678
rect 66668 3602 66724 3612
rect 68460 3668 68516 3678
rect 68460 3602 68516 3612
rect 70252 3668 70308 3678
rect 70252 3602 70308 3612
rect 71148 3668 71204 3678
rect 71148 3602 71204 3612
rect 73388 3668 73444 3678
rect 73388 3602 73444 3612
rect 74732 3668 74788 3678
rect 74732 3602 74788 3612
rect 76972 3668 77028 3678
rect 76972 3602 77028 3612
rect 78540 3668 78596 3678
rect 78540 3602 78596 3612
rect 81452 3668 81508 3678
rect 81452 3602 81508 3612
rect 82124 3668 82180 3678
rect 82124 3602 82180 3612
rect 83020 3668 83076 3678
rect 83020 3602 83076 3612
rect 83468 3668 83524 3678
rect 83468 3602 83524 3612
rect 84812 3668 84868 3678
rect 84812 3602 84868 3612
rect 32508 3556 32564 3566
rect 11564 3444 11620 3454
rect 11564 480 11620 3388
rect 15372 3108 15428 3118
rect 13356 1092 13412 1102
rect 13356 480 13412 1036
rect 15372 480 15428 3052
rect 26796 980 26852 990
rect 24892 644 24948 654
rect 23100 532 23156 542
rect 17276 480 17444 532
rect 19180 480 19348 532
rect 21084 480 21252 532
rect 22988 480 23100 532
rect 11368 392 11620 480
rect 11368 -960 11592 392
rect 13272 -960 13496 480
rect 15176 392 15428 480
rect 17080 476 17444 480
rect 17080 392 17332 476
rect 15176 -960 15400 392
rect 17080 -960 17304 392
rect 17388 196 17444 476
rect 17388 130 17444 140
rect 18984 476 19348 480
rect 18984 392 19236 476
rect 18984 -960 19208 392
rect 19292 308 19348 476
rect 19292 242 19348 252
rect 20888 476 21252 480
rect 20888 392 21140 476
rect 21196 420 21252 476
rect 22792 476 23100 480
rect 24892 480 24948 588
rect 26796 480 26852 924
rect 30604 868 30660 878
rect 28700 756 28756 766
rect 28700 480 28756 700
rect 30604 480 30660 812
rect 32508 480 32564 3500
rect 37100 3556 37156 3566
rect 37100 3490 37156 3500
rect 46060 3556 46116 3566
rect 46060 3490 46116 3500
rect 46956 3556 47012 3566
rect 46956 3490 47012 3500
rect 47852 3556 47908 3566
rect 47852 3490 47908 3500
rect 49644 3556 49700 3566
rect 49644 3490 49700 3500
rect 51660 3556 51716 3566
rect 51660 3490 51716 3500
rect 52780 3556 52836 3566
rect 52780 3490 52836 3500
rect 54572 3556 54628 3566
rect 54572 3490 54628 3500
rect 56364 3556 56420 3566
rect 56364 3490 56420 3500
rect 58380 3556 58436 3566
rect 58380 3490 58436 3500
rect 59052 3556 59108 3566
rect 59052 3490 59108 3500
rect 61740 3556 61796 3566
rect 61740 3490 61796 3500
rect 67564 3556 67620 3566
rect 67564 3490 67620 3500
rect 76524 3556 76580 3566
rect 76524 3490 76580 3500
rect 77420 3556 77476 3566
rect 77420 3490 77476 3500
rect 80556 3556 80612 3566
rect 80556 3490 80612 3500
rect 83916 3556 83972 3566
rect 83916 3490 83972 3500
rect 104636 3556 104692 3566
rect 34636 3444 34692 3454
rect 34636 3378 34692 3388
rect 38892 3444 38948 3454
rect 38892 3378 38948 3388
rect 46508 3444 46564 3454
rect 46508 3378 46564 3388
rect 47404 3444 47460 3454
rect 47404 3378 47460 3388
rect 48748 3444 48804 3454
rect 48748 3378 48804 3388
rect 51436 3444 51492 3454
rect 51436 3378 51492 3388
rect 53004 3444 53060 3454
rect 53004 3378 53060 3388
rect 70700 3444 70756 3454
rect 70700 3378 70756 3388
rect 86380 3444 86436 3454
rect 86380 3378 86436 3388
rect 88172 3444 88228 3454
rect 88172 3378 88228 3388
rect 90188 3444 90244 3454
rect 90188 3378 90244 3388
rect 91980 3444 92036 3454
rect 91980 3378 92036 3388
rect 92876 3444 92932 3454
rect 92876 3378 92932 3388
rect 93324 3444 93380 3454
rect 93324 3378 93380 3388
rect 95340 3444 95396 3454
rect 95340 3378 95396 3388
rect 96684 3444 96740 3454
rect 96684 3378 96740 3388
rect 98028 3444 98084 3454
rect 98028 3378 98084 3388
rect 100044 3444 100100 3454
rect 102060 3444 102116 3454
rect 101192 3388 102060 3444
rect 100044 3378 100100 3388
rect 102060 3378 102116 3388
rect 43596 3332 43652 3342
rect 43596 3266 43652 3276
rect 45836 3332 45892 3342
rect 45836 3266 45892 3276
rect 50092 3332 50148 3342
rect 50092 3266 50148 3276
rect 54796 3332 54852 3342
rect 54796 3266 54852 3276
rect 56140 3332 56196 3342
rect 56140 3266 56196 3276
rect 57484 3332 57540 3342
rect 57484 3266 57540 3276
rect 59948 3332 60004 3342
rect 59948 3266 60004 3276
rect 60620 3332 60676 3342
rect 60620 3266 60676 3276
rect 63756 3332 63812 3342
rect 63756 3266 63812 3276
rect 79436 3332 79492 3342
rect 79436 3266 79492 3276
rect 84364 3332 84420 3342
rect 84364 3266 84420 3276
rect 91532 3332 91588 3342
rect 91532 3266 91588 3276
rect 93996 3332 94052 3342
rect 93996 3266 94052 3276
rect 94668 3332 94724 3342
rect 94668 3266 94724 3276
rect 95788 3332 95844 3342
rect 95788 3266 95844 3276
rect 97580 3332 97636 3342
rect 97580 3266 97636 3276
rect 40684 3220 40740 3230
rect 40684 3154 40740 3164
rect 62636 3220 62692 3230
rect 62636 3154 62692 3164
rect 67340 3220 67396 3230
rect 67340 3154 67396 3164
rect 72044 3220 72100 3230
rect 72044 3154 72100 3164
rect 73164 3220 73220 3230
rect 73164 3154 73220 3164
rect 75180 3220 75236 3230
rect 75180 3154 75236 3164
rect 76748 3220 76804 3230
rect 76748 3154 76804 3164
rect 92652 3220 92708 3230
rect 92652 3154 92708 3164
rect 95564 3220 95620 3230
rect 95564 3154 95620 3164
rect 98252 3220 98308 3230
rect 98252 3154 98308 3164
rect 98924 3220 98980 3230
rect 98924 3154 98980 3164
rect 35084 3108 35140 3118
rect 34412 1540 34468 1550
rect 34412 480 34468 1484
rect 34860 1092 34916 3080
rect 42252 3108 42308 3118
rect 35084 3042 35140 3052
rect 34860 1026 34916 1036
rect 21756 420 21812 430
rect 20888 -960 21112 392
rect 21196 364 21756 420
rect 21756 354 21812 364
rect 22792 392 23044 476
rect 23100 466 23156 476
rect 24696 392 24948 480
rect 26600 392 26852 480
rect 28504 392 28756 480
rect 30408 392 30660 480
rect 32312 392 32564 480
rect 34216 392 34468 480
rect 22792 -960 23016 392
rect 24696 -960 24920 392
rect 26600 -960 26824 392
rect 28504 -960 28728 392
rect 30408 -960 30632 392
rect 32312 -960 32536 392
rect 34216 -960 34440 392
rect 35308 196 35364 3080
rect 35420 1204 35476 1214
rect 35420 644 35476 1148
rect 35420 578 35476 588
rect 35420 308 35476 318
rect 35532 308 35588 3080
rect 35756 420 35812 3080
rect 35980 532 36036 3080
rect 36204 1204 36260 3080
rect 36204 1138 36260 1148
rect 36428 980 36484 3080
rect 36652 1428 36708 3080
rect 36652 1362 36708 1372
rect 36428 914 36484 924
rect 36876 868 36932 3080
rect 37324 1876 37380 3080
rect 36988 1820 37380 1876
rect 36988 1540 37044 1820
rect 37548 1652 37604 3080
rect 36988 1474 37044 1484
rect 37100 1596 37604 1652
rect 37772 1652 37828 3080
rect 37996 1764 38052 3080
rect 37996 1708 38164 1764
rect 37772 1596 38052 1652
rect 36876 802 36932 812
rect 36316 480 36484 532
rect 35980 466 36036 476
rect 36120 476 36484 480
rect 35756 354 35812 364
rect 36120 392 36372 476
rect 36428 420 36484 476
rect 37100 420 37156 1596
rect 35476 252 35588 308
rect 35420 242 35476 252
rect 35308 130 35364 140
rect 36120 -960 36344 392
rect 36428 364 37156 420
rect 37996 480 38052 1596
rect 38108 1540 38164 1708
rect 38220 1652 38276 3080
rect 38220 1586 38276 1596
rect 38108 1474 38164 1484
rect 38444 1428 38500 3080
rect 38444 1362 38500 1372
rect 38668 980 38724 3080
rect 39116 1316 39172 3080
rect 39116 1250 39172 1260
rect 38668 914 38724 924
rect 37996 392 38248 480
rect 38024 -960 38248 392
rect 39228 84 39284 94
rect 39340 84 39396 3080
rect 39788 868 39844 3080
rect 39788 802 39844 812
rect 39900 1540 39956 1550
rect 39900 480 39956 1484
rect 40236 1540 40292 3080
rect 40460 2660 40516 3080
rect 41132 2772 41188 3080
rect 41132 2706 41188 2716
rect 40460 2594 40516 2604
rect 41580 2548 41636 3080
rect 41804 2884 41860 3080
rect 43820 3108 43876 3118
rect 42252 3042 42308 3052
rect 41804 2818 41860 2828
rect 41580 2482 41636 2492
rect 40796 1652 40852 1662
rect 40852 1596 41076 1652
rect 40796 1586 40852 1596
rect 40236 1474 40292 1484
rect 39900 392 40152 480
rect 39284 28 39396 84
rect 39228 18 39284 28
rect 39928 -960 40152 392
rect 41020 420 41076 1596
rect 42476 532 42532 3080
rect 42924 2436 42980 3080
rect 42924 2370 42980 2380
rect 43372 1092 43428 3080
rect 56588 3108 56644 3118
rect 43820 3042 43876 3052
rect 44044 1652 44100 3080
rect 44044 1586 44100 1596
rect 44492 1652 44548 3080
rect 44492 1586 44548 1596
rect 43372 1026 43428 1036
rect 43708 1428 43764 1438
rect 41692 480 41860 532
rect 41692 476 42056 480
rect 41692 420 41748 476
rect 41020 364 41748 420
rect 41804 392 42056 476
rect 42476 466 42532 476
rect 43708 480 43764 1372
rect 45164 532 45220 3080
rect 45388 1204 45444 3080
rect 47180 1428 47236 3080
rect 47180 1362 47236 1372
rect 47516 2324 47572 2334
rect 45388 1138 45444 1148
rect 43708 392 43960 480
rect 45164 466 45220 476
rect 45612 980 45668 990
rect 45612 480 45668 924
rect 47516 480 47572 2268
rect 48076 1652 48132 3080
rect 48076 1586 48132 1596
rect 49420 1540 49476 3080
rect 49308 1484 49476 1540
rect 49308 980 49364 1484
rect 50764 1428 50820 3080
rect 50764 1362 50820 1372
rect 49308 914 49364 924
rect 49420 1316 49476 1326
rect 49420 480 49476 1260
rect 52108 756 52164 3080
rect 52556 1316 52612 3080
rect 52556 1250 52612 1260
rect 53228 2324 53284 2334
rect 52108 690 52164 700
rect 51212 480 51380 532
rect 53228 480 53284 2268
rect 53452 1652 53508 3080
rect 53452 1586 53508 1596
rect 55244 1540 55300 3080
rect 55244 1474 55300 1484
rect 55468 980 55524 3080
rect 62188 3108 62244 3118
rect 56588 3042 56644 3052
rect 55468 914 55524 924
rect 55020 868 55076 878
rect 55076 812 55188 868
rect 55020 802 55076 812
rect 55132 480 55188 812
rect 56812 644 56868 3080
rect 57148 2324 57204 2334
rect 56812 578 56868 588
rect 56924 2100 56980 2110
rect 56924 532 56980 2044
rect 45612 392 45864 480
rect 47516 392 47768 480
rect 49420 392 49672 480
rect 41832 -960 42056 392
rect 43736 -960 43960 392
rect 45640 -960 45864 392
rect 47544 -960 47768 392
rect 49448 -960 49672 392
rect 51212 476 51576 480
rect 51212 84 51268 476
rect 51324 392 51576 476
rect 53228 392 53480 480
rect 55132 392 55384 480
rect 57148 480 57204 2268
rect 58156 1652 58212 3080
rect 60956 2660 61012 2670
rect 58156 1586 58212 1596
rect 58940 2324 58996 2334
rect 58940 480 58996 2268
rect 60956 480 61012 2604
rect 61516 1652 61572 3080
rect 68012 3108 68068 3118
rect 62188 3042 62244 3052
rect 61516 1586 61572 1596
rect 62412 1540 62468 3080
rect 62972 2660 63028 2670
rect 63308 2660 63364 3080
rect 63028 2604 63364 2660
rect 64764 2660 64820 2670
rect 62972 2594 63028 2604
rect 62412 1474 62468 1484
rect 62748 2324 62804 2334
rect 62748 480 62804 2268
rect 64764 480 64820 2604
rect 65772 1540 65828 3080
rect 66444 1652 66500 3080
rect 66444 1586 66500 1596
rect 66556 2772 66612 2782
rect 65772 1474 65828 1484
rect 66556 480 66612 2716
rect 66892 532 66948 3080
rect 68012 3042 68068 3052
rect 68236 3108 68292 3118
rect 74284 3108 74340 3118
rect 68236 3042 68292 3052
rect 56924 466 56980 476
rect 51212 18 51268 28
rect 51352 -960 51576 392
rect 53256 -960 53480 392
rect 55160 -960 55384 392
rect 57064 -960 57288 480
rect 58940 392 59192 480
rect 58968 -960 59192 392
rect 60872 -960 61096 480
rect 62748 392 63000 480
rect 62776 -960 63000 392
rect 64680 -960 64904 480
rect 66556 392 66808 480
rect 68572 2772 68628 2782
rect 68572 480 68628 2716
rect 68796 2324 68852 2334
rect 68796 1204 68852 2268
rect 69580 1652 69636 3080
rect 69580 1586 69636 1596
rect 70028 1652 70084 3080
rect 70028 1586 70084 1596
rect 70364 2212 70420 2222
rect 68796 1138 68852 1148
rect 70364 480 70420 2156
rect 70924 1204 70980 3080
rect 71372 2772 71428 3080
rect 72380 2884 72436 2894
rect 71708 2772 71764 2782
rect 71372 2716 71708 2772
rect 71708 2706 71764 2716
rect 72156 2212 72212 2222
rect 72156 1428 72212 2156
rect 72156 1362 72212 1372
rect 70924 1138 70980 1148
rect 72380 480 72436 2828
rect 74060 1316 74116 3080
rect 78092 3108 78148 3118
rect 74284 3042 74340 3052
rect 74060 1250 74116 1260
rect 74172 2884 74228 2894
rect 74172 480 74228 2828
rect 75628 2548 75684 3080
rect 75628 2482 75684 2492
rect 76188 2772 76244 2782
rect 76188 480 76244 2716
rect 76300 1652 76356 3080
rect 78092 3042 78148 3052
rect 76300 1586 76356 1596
rect 77980 2660 78036 2670
rect 77980 480 78036 2604
rect 78316 1428 78372 3080
rect 78316 1362 78372 1372
rect 66892 466 66948 476
rect 66584 -960 66808 392
rect 68488 -960 68712 480
rect 70364 392 70616 480
rect 70392 -960 70616 392
rect 72296 -960 72520 480
rect 74172 392 74424 480
rect 74200 -960 74424 392
rect 76104 -960 76328 480
rect 77980 392 78232 480
rect 78008 -960 78232 392
rect 78764 308 78820 3080
rect 78988 2772 79044 3080
rect 79100 2772 79156 2782
rect 78988 2716 79100 2772
rect 79100 2706 79156 2716
rect 78876 2548 78932 2558
rect 78876 1540 78932 2492
rect 79660 1652 79716 3080
rect 79660 1586 79716 1596
rect 79996 2884 80052 2894
rect 78876 1474 78932 1484
rect 79996 480 80052 2828
rect 80332 1316 80388 3080
rect 81004 1540 81060 3080
rect 81004 1474 81060 1484
rect 80332 1250 80388 1260
rect 81676 1316 81732 3080
rect 81676 1250 81732 1260
rect 81788 2436 81844 2446
rect 81788 480 81844 2380
rect 82348 1316 82404 3080
rect 82348 1250 82404 1260
rect 83804 2884 83860 2894
rect 83804 480 83860 2828
rect 85036 1092 85092 3080
rect 85484 1652 85540 3080
rect 85708 2660 85764 3080
rect 85708 2594 85764 2604
rect 85484 1586 85540 1596
rect 85708 1764 85764 1774
rect 85036 1026 85092 1036
rect 85708 480 85764 1708
rect 87052 1540 87108 3080
rect 87052 1474 87108 1484
rect 87500 2884 87556 2894
rect 87500 480 87556 2828
rect 87724 1204 87780 3080
rect 87724 1138 87780 1148
rect 88396 532 88452 3080
rect 78764 242 78820 252
rect 79912 -960 80136 480
rect 81788 392 82040 480
rect 81816 -960 82040 392
rect 83720 -960 83944 480
rect 85624 -960 85848 480
rect 87500 392 87752 480
rect 88396 466 88452 476
rect 89404 1764 89460 1774
rect 89404 480 89460 1708
rect 89740 1540 89796 3080
rect 90412 2884 90468 3080
rect 90412 2818 90468 2828
rect 91084 2772 91140 3080
rect 91084 2706 91140 2716
rect 89740 1474 89796 1484
rect 91308 2212 91364 2222
rect 91308 480 91364 2156
rect 91756 1652 91812 3080
rect 91756 1586 91812 1596
rect 92428 868 92484 3080
rect 92428 802 92484 812
rect 93212 2660 93268 2670
rect 93212 480 93268 2604
rect 93772 1092 93828 3080
rect 94444 1204 94500 3080
rect 95116 1428 95172 3080
rect 95228 2884 95284 2894
rect 95900 2884 95956 2894
rect 95284 2828 95900 2884
rect 95228 2818 95284 2828
rect 95900 2818 95956 2828
rect 95116 1362 95172 1372
rect 95228 2660 95284 2670
rect 94444 1138 94500 1148
rect 93772 1026 93828 1036
rect 95228 480 95284 2604
rect 95676 2660 95732 2670
rect 95676 1316 95732 2604
rect 96460 1428 96516 3080
rect 96460 1362 96516 1372
rect 97020 2772 97076 2782
rect 95676 1250 95732 1260
rect 97020 480 97076 2716
rect 97132 1540 97188 3080
rect 97804 1540 97860 3080
rect 98476 1652 98532 3080
rect 98476 1586 98532 1596
rect 99036 2772 99092 2782
rect 97132 1484 97412 1540
rect 97356 756 97412 1484
rect 97804 1474 97860 1484
rect 97356 690 97412 700
rect 99036 480 99092 2716
rect 99148 1652 99204 3080
rect 99148 1586 99204 1596
rect 100492 1652 100548 3080
rect 102732 2324 102788 2334
rect 100492 1586 100548 1596
rect 100828 2100 100884 2110
rect 100828 480 100884 2044
rect 102732 480 102788 2268
rect 104636 480 104692 3500
rect 106540 3556 106596 3566
rect 106540 480 106596 3500
rect 108444 3556 108500 3566
rect 108444 480 108500 3500
rect 110348 3556 110404 3566
rect 110348 480 110404 3500
rect 112252 3556 112308 3566
rect 112252 480 112308 3500
rect 116060 3556 116116 3566
rect 114268 3444 114324 3454
rect 114268 480 114324 3388
rect 116060 480 116116 3500
rect 119868 3556 119924 3566
rect 117964 2100 118020 2110
rect 117964 480 118020 2044
rect 119868 480 119924 3500
rect 121772 3556 121828 3566
rect 121772 480 121828 3500
rect 123564 3220 123620 6860
rect 123564 3154 123620 3164
rect 123676 480 123732 80780
rect 124012 8708 124068 8718
rect 124012 2660 124068 8652
rect 124012 2594 124068 2604
rect 125580 480 125636 82348
rect 127036 16884 127092 16894
rect 127036 868 127092 16828
rect 127036 802 127092 812
rect 127484 4228 127540 4238
rect 127484 480 127540 4172
rect 129388 480 129444 82460
rect 315980 80724 316036 80734
rect 272188 79828 272244 79838
rect 218876 76468 218932 76478
rect 213164 73444 213220 73454
rect 205548 4452 205604 4462
rect 131292 4228 131348 4238
rect 131292 480 131348 4172
rect 133196 4228 133252 4238
rect 133196 480 133252 4172
rect 135100 4228 135156 4238
rect 135100 480 135156 4172
rect 138908 4228 138964 4238
rect 137004 4116 137060 4126
rect 137004 480 137060 4060
rect 138908 480 138964 4172
rect 140812 4228 140868 4238
rect 140812 480 140868 4172
rect 142828 4228 142884 4238
rect 142828 480 142884 4172
rect 144620 4228 144676 4238
rect 144620 480 144676 4172
rect 146524 4228 146580 4238
rect 146524 480 146580 4172
rect 148428 4228 148484 4238
rect 148428 480 148484 4172
rect 150332 4228 150388 4238
rect 150332 480 150388 4172
rect 152236 4228 152292 4238
rect 152236 480 152292 4172
rect 154140 4228 154196 4238
rect 154140 480 154196 4172
rect 156044 4228 156100 4238
rect 156044 480 156100 4172
rect 157948 4228 158004 4238
rect 157948 480 158004 4172
rect 161756 4228 161812 4238
rect 159852 4004 159908 4014
rect 159852 480 159908 3948
rect 161756 480 161812 4172
rect 163660 4228 163716 4238
rect 163660 480 163716 4172
rect 165564 4228 165620 4238
rect 165564 480 165620 4172
rect 167468 4228 167524 4238
rect 167468 480 167524 4172
rect 169372 4228 169428 4238
rect 169372 480 169428 4172
rect 173180 4228 173236 4238
rect 171388 3892 171444 3902
rect 171388 480 171444 3836
rect 173180 480 173236 4172
rect 175084 4228 175140 4238
rect 175084 480 175140 4172
rect 178892 4228 178948 4238
rect 176988 3780 177044 3790
rect 176988 480 177044 3724
rect 178892 480 178948 4172
rect 180796 4228 180852 4238
rect 180796 480 180852 4172
rect 184604 4228 184660 4238
rect 182700 3556 182756 3566
rect 182700 480 182756 3500
rect 184604 480 184660 4172
rect 190428 4228 190484 4238
rect 186508 1988 186564 1998
rect 186508 480 186564 1932
rect 188412 980 188468 990
rect 188412 480 188468 924
rect 190428 480 190484 4172
rect 192220 4228 192276 4238
rect 192220 480 192276 4172
rect 196028 4228 196084 4238
rect 194124 3444 194180 3454
rect 194124 480 194180 3388
rect 196028 480 196084 4172
rect 201740 4228 201796 4238
rect 197932 1988 197988 1998
rect 197932 480 197988 1932
rect 199724 480 199892 532
rect 201740 480 201796 4172
rect 203644 4228 203700 4238
rect 203644 480 203700 4172
rect 205548 480 205604 4396
rect 207452 4228 207508 4238
rect 207452 480 207508 4172
rect 209356 3668 209412 3678
rect 209356 480 209412 3612
rect 211260 644 211316 654
rect 211260 480 211316 588
rect 213164 480 213220 73388
rect 215068 4228 215124 4238
rect 215068 480 215124 4172
rect 216972 4228 217028 4238
rect 216972 480 217028 4172
rect 218876 480 218932 76412
rect 230300 76356 230356 76366
rect 226492 73332 226548 73342
rect 220780 4228 220836 4238
rect 220780 480 220836 4172
rect 222684 4228 222740 4238
rect 222684 480 222740 4172
rect 224588 4228 224644 4238
rect 224588 480 224644 4172
rect 226492 480 226548 73276
rect 228508 4228 228564 4238
rect 228508 480 228564 4172
rect 230300 480 230356 76300
rect 247436 76244 247492 76254
rect 241724 74788 241780 74798
rect 232204 4228 232260 4238
rect 232204 480 232260 4172
rect 234108 4228 234164 4238
rect 234108 480 234164 4172
rect 236012 4228 236068 4238
rect 236012 480 236068 4172
rect 237916 4228 237972 4238
rect 237916 480 237972 4172
rect 239820 4228 239876 4238
rect 239820 480 239876 4172
rect 241724 480 241780 74732
rect 243628 4228 243684 4238
rect 243628 480 243684 4172
rect 245532 4228 245588 4238
rect 245532 480 245588 4172
rect 247436 480 247492 76188
rect 270284 74676 270340 74686
rect 249340 4228 249396 4238
rect 249340 480 249396 4172
rect 251244 4228 251300 4238
rect 251244 480 251300 4172
rect 253148 4228 253204 4238
rect 253148 480 253204 4172
rect 255052 4228 255108 4238
rect 255052 480 255108 4172
rect 258860 4228 258916 4238
rect 257068 3556 257124 3566
rect 257068 480 257124 3500
rect 258860 480 258916 4172
rect 260764 4228 260820 4238
rect 260764 480 260820 4172
rect 262668 4228 262724 4238
rect 262668 480 262724 4172
rect 264572 4228 264628 4238
rect 264572 480 264628 4172
rect 266476 4228 266532 4238
rect 266476 480 266532 4172
rect 268380 3444 268436 3454
rect 268380 480 268436 3388
rect 270284 480 270340 74620
rect 272188 480 272244 79772
rect 310268 78260 310324 78270
rect 281708 74564 281764 74574
rect 275996 73108 276052 73118
rect 274092 4228 274148 4238
rect 274092 480 274148 4172
rect 275996 480 276052 73052
rect 277900 72884 277956 72894
rect 277900 480 277956 72828
rect 279804 4228 279860 4238
rect 279804 480 279860 4172
rect 281708 480 281764 74508
rect 293132 74452 293188 74462
rect 287420 72996 287476 73006
rect 283612 4228 283668 4238
rect 283612 480 283668 4172
rect 285740 4228 285796 4238
rect 285740 480 285796 4172
rect 89404 392 89656 480
rect 91308 392 91560 480
rect 93212 392 93464 480
rect 87528 -960 87752 392
rect 89432 -960 89656 392
rect 91336 -960 91560 392
rect 93240 -960 93464 392
rect 95144 -960 95368 480
rect 97020 392 97272 480
rect 97048 -960 97272 392
rect 98952 -960 99176 480
rect 100828 392 101080 480
rect 102732 392 102984 480
rect 104636 392 104888 480
rect 106540 392 106792 480
rect 108444 392 108696 480
rect 110348 392 110600 480
rect 112252 392 112504 480
rect 100856 -960 101080 392
rect 102760 -960 102984 392
rect 104664 -960 104888 392
rect 106568 -960 106792 392
rect 108472 -960 108696 392
rect 110376 -960 110600 392
rect 112280 -960 112504 392
rect 114184 -960 114408 480
rect 116060 392 116312 480
rect 117964 392 118216 480
rect 119868 392 120120 480
rect 121772 392 122024 480
rect 123676 392 123928 480
rect 125580 392 125832 480
rect 127484 392 127736 480
rect 129388 392 129640 480
rect 131292 392 131544 480
rect 133196 392 133448 480
rect 135100 392 135352 480
rect 137004 392 137256 480
rect 138908 392 139160 480
rect 140812 392 141064 480
rect 116088 -960 116312 392
rect 117992 -960 118216 392
rect 119896 -960 120120 392
rect 121800 -960 122024 392
rect 123704 -960 123928 392
rect 125608 -960 125832 392
rect 127512 -960 127736 392
rect 129416 -960 129640 392
rect 131320 -960 131544 392
rect 133224 -960 133448 392
rect 135128 -960 135352 392
rect 137032 -960 137256 392
rect 138936 -960 139160 392
rect 140840 -960 141064 392
rect 142744 -960 142968 480
rect 144620 392 144872 480
rect 146524 392 146776 480
rect 148428 392 148680 480
rect 150332 392 150584 480
rect 152236 392 152488 480
rect 154140 392 154392 480
rect 156044 392 156296 480
rect 157948 392 158200 480
rect 159852 392 160104 480
rect 161756 392 162008 480
rect 163660 392 163912 480
rect 165564 392 165816 480
rect 167468 392 167720 480
rect 169372 392 169624 480
rect 144648 -960 144872 392
rect 146552 -960 146776 392
rect 148456 -960 148680 392
rect 150360 -960 150584 392
rect 152264 -960 152488 392
rect 154168 -960 154392 392
rect 156072 -960 156296 392
rect 157976 -960 158200 392
rect 159880 -960 160104 392
rect 161784 -960 162008 392
rect 163688 -960 163912 392
rect 165592 -960 165816 392
rect 167496 -960 167720 392
rect 169400 -960 169624 392
rect 171304 -960 171528 480
rect 173180 392 173432 480
rect 175084 392 175336 480
rect 176988 392 177240 480
rect 178892 392 179144 480
rect 180796 392 181048 480
rect 182700 392 182952 480
rect 184604 392 184856 480
rect 186508 392 186760 480
rect 188412 392 188664 480
rect 173208 -960 173432 392
rect 175112 -960 175336 392
rect 177016 -960 177240 392
rect 178920 -960 179144 392
rect 180824 -960 181048 392
rect 182728 -960 182952 392
rect 184632 -960 184856 392
rect 186536 -960 186760 392
rect 188440 -960 188664 392
rect 190344 -960 190568 480
rect 192220 392 192472 480
rect 194124 392 194376 480
rect 196028 392 196280 480
rect 197932 392 198184 480
rect 192248 -960 192472 392
rect 194152 -960 194376 392
rect 196056 -960 196280 392
rect 197960 -960 198184 392
rect 199724 476 200088 480
rect 199724 84 199780 476
rect 199836 392 200088 476
rect 201740 392 201992 480
rect 203644 392 203896 480
rect 205548 392 205800 480
rect 207452 392 207704 480
rect 209356 392 209608 480
rect 211260 392 211512 480
rect 213164 392 213416 480
rect 215068 392 215320 480
rect 216972 392 217224 480
rect 218876 392 219128 480
rect 220780 392 221032 480
rect 222684 392 222936 480
rect 224588 392 224840 480
rect 226492 392 226744 480
rect 199724 18 199780 28
rect 199864 -960 200088 392
rect 201768 -960 201992 392
rect 203672 -960 203896 392
rect 205576 -960 205800 392
rect 207480 -960 207704 392
rect 209384 -960 209608 392
rect 211288 -960 211512 392
rect 213192 -960 213416 392
rect 215096 -960 215320 392
rect 217000 -960 217224 392
rect 218904 -960 219128 392
rect 220808 -960 221032 392
rect 222712 -960 222936 392
rect 224616 -960 224840 392
rect 226520 -960 226744 392
rect 228424 -960 228648 480
rect 230300 392 230552 480
rect 232204 392 232456 480
rect 234108 392 234360 480
rect 236012 392 236264 480
rect 237916 392 238168 480
rect 239820 392 240072 480
rect 241724 392 241976 480
rect 243628 392 243880 480
rect 245532 392 245784 480
rect 247436 392 247688 480
rect 249340 392 249592 480
rect 251244 392 251496 480
rect 253148 392 253400 480
rect 255052 392 255304 480
rect 230328 -960 230552 392
rect 232232 -960 232456 392
rect 234136 -960 234360 392
rect 236040 -960 236264 392
rect 237944 -960 238168 392
rect 239848 -960 240072 392
rect 241752 -960 241976 392
rect 243656 -960 243880 392
rect 245560 -960 245784 392
rect 247464 -960 247688 392
rect 249368 -960 249592 392
rect 251272 -960 251496 392
rect 253176 -960 253400 392
rect 255080 -960 255304 392
rect 256984 -960 257208 480
rect 258860 392 259112 480
rect 260764 392 261016 480
rect 262668 392 262920 480
rect 264572 392 264824 480
rect 266476 392 266728 480
rect 268380 392 268632 480
rect 270284 392 270536 480
rect 272188 392 272440 480
rect 274092 392 274344 480
rect 275996 392 276248 480
rect 277900 392 278152 480
rect 279804 392 280056 480
rect 281708 392 281960 480
rect 283612 392 283864 480
rect 258888 -960 259112 392
rect 260792 -960 261016 392
rect 262696 -960 262920 392
rect 264600 -960 264824 392
rect 266504 -960 266728 392
rect 268408 -960 268632 392
rect 270312 -960 270536 392
rect 272216 -960 272440 392
rect 274120 -960 274344 392
rect 276024 -960 276248 392
rect 277928 -960 278152 392
rect 279832 -960 280056 392
rect 281736 -960 281960 392
rect 283640 -960 283864 392
rect 285544 392 285796 480
rect 287420 480 287476 72940
rect 289324 4228 289380 4238
rect 289324 480 289380 4172
rect 291228 4228 291284 4238
rect 291228 480 291284 4172
rect 293132 480 293188 74396
rect 304556 74340 304612 74350
rect 298844 72772 298900 72782
rect 295036 4228 295092 4238
rect 295036 480 295092 4172
rect 296940 4228 296996 4238
rect 296940 480 296996 4172
rect 298844 480 298900 72716
rect 299068 7028 299124 7038
rect 299068 1092 299124 6972
rect 299068 1026 299124 1036
rect 300748 4228 300804 4238
rect 300748 480 300804 4172
rect 302652 4228 302708 4238
rect 302652 480 302708 4172
rect 304556 480 304612 74284
rect 306460 4228 306516 4238
rect 306460 480 306516 4172
rect 308364 3444 308420 3454
rect 308364 480 308420 3388
rect 310268 480 310324 78204
rect 312172 4228 312228 4238
rect 312172 480 312228 4172
rect 314188 4228 314244 4238
rect 314188 480 314244 4172
rect 315980 480 316036 80668
rect 430220 79940 430276 79950
rect 355964 79716 356020 79726
rect 321692 78148 321748 78158
rect 317884 4228 317940 4238
rect 317884 480 317940 4172
rect 319788 4228 319844 4238
rect 319788 480 319844 4172
rect 321692 480 321748 78092
rect 327404 78036 327460 78046
rect 323596 4228 323652 4238
rect 323596 480 323652 4172
rect 325500 4228 325556 4238
rect 325500 480 325556 4172
rect 327404 480 327460 77980
rect 329308 77924 329364 77934
rect 329308 480 329364 77868
rect 350252 77812 350308 77822
rect 333116 76132 333172 76142
rect 331212 4228 331268 4238
rect 331212 480 331268 4172
rect 333116 480 333172 76076
rect 344540 76020 344596 76030
rect 335020 74228 335076 74238
rect 335020 480 335076 74172
rect 338828 73556 338884 73566
rect 336924 4228 336980 4238
rect 336924 480 336980 4172
rect 338828 480 338884 73500
rect 340732 4228 340788 4238
rect 340732 480 340788 4172
rect 342748 4228 342804 4238
rect 342748 480 342804 4172
rect 344540 480 344596 75964
rect 346444 4228 346500 4238
rect 346444 480 346500 4172
rect 348348 4228 348404 4238
rect 348348 480 348404 4172
rect 350252 480 350308 77756
rect 352156 4228 352212 4238
rect 352156 480 352212 4172
rect 354060 4228 354116 4238
rect 354060 480 354116 4172
rect 355964 480 356020 79660
rect 361676 79604 361732 79614
rect 357868 75908 357924 75918
rect 357868 480 357924 75852
rect 359772 4228 359828 4238
rect 359772 480 359828 4172
rect 361676 480 361732 79548
rect 369292 79492 369348 79502
rect 367388 74116 367444 74126
rect 363580 4228 363636 4238
rect 363580 480 363636 4172
rect 365484 4228 365540 4238
rect 365484 480 365540 4172
rect 367388 480 367444 74060
rect 369292 480 369348 79436
rect 373100 79380 373156 79390
rect 371308 4228 371364 4238
rect 371308 480 371364 4172
rect 373100 480 373156 79324
rect 378812 79268 378868 79278
rect 375004 4228 375060 4238
rect 375004 480 375060 4172
rect 376908 4228 376964 4238
rect 376908 480 376964 4172
rect 378812 480 378868 79212
rect 413084 79156 413140 79166
rect 390236 77700 390292 77710
rect 380716 4228 380772 4238
rect 380716 480 380772 4172
rect 384524 4228 384580 4238
rect 382620 1876 382676 1886
rect 382620 480 382676 1820
rect 384524 480 384580 4172
rect 386428 4228 386484 4238
rect 386428 480 386484 4172
rect 388332 4228 388388 4238
rect 388332 480 388388 4172
rect 390236 480 390292 77644
rect 401660 75796 401716 75806
rect 399868 8708 399924 8718
rect 392140 4228 392196 4238
rect 392140 480 392196 4172
rect 394044 4228 394100 4238
rect 394044 480 394100 4172
rect 395948 4228 396004 4238
rect 395948 480 396004 4172
rect 397852 4228 397908 4238
rect 397852 480 397908 4172
rect 399868 480 399924 8652
rect 401660 480 401716 75740
rect 403564 4228 403620 4238
rect 403564 480 403620 4172
rect 407372 4228 407428 4238
rect 405468 1764 405524 1774
rect 405468 480 405524 1708
rect 407372 480 407428 4172
rect 411180 4228 411236 4238
rect 409276 3444 409332 3454
rect 409276 480 409332 3388
rect 411180 480 411236 4172
rect 413084 480 413140 79100
rect 424508 77588 424564 77598
rect 418796 74900 418852 74910
rect 416892 4228 416948 4238
rect 414988 3444 415044 3454
rect 414988 480 415044 3388
rect 416892 480 416948 4172
rect 418796 480 418852 74844
rect 420700 4228 420756 4238
rect 420700 480 420756 4172
rect 422604 4228 422660 4238
rect 422604 480 422660 4172
rect 424508 480 424564 77532
rect 426412 4228 426468 4238
rect 426412 480 426468 4172
rect 428428 4228 428484 4238
rect 426748 1764 426804 1774
rect 426748 1204 426804 1708
rect 426748 1138 426804 1148
rect 428428 480 428484 4172
rect 430220 480 430276 79884
rect 441644 77476 441700 77486
rect 434028 11060 434084 11070
rect 432124 4228 432180 4238
rect 432124 480 432180 4172
rect 434028 480 434084 11004
rect 435932 4228 435988 4238
rect 435932 480 435988 4172
rect 437836 4228 437892 4238
rect 437836 480 437892 4172
rect 439740 4228 439796 4238
rect 439740 480 439796 4172
rect 441644 480 441700 77420
rect 569212 77364 569268 77374
rect 464492 76580 464548 76590
rect 443548 4228 443604 4238
rect 443548 480 443604 4172
rect 447356 4228 447412 4238
rect 445452 2548 445508 2558
rect 445452 480 445508 2492
rect 447356 480 447412 4172
rect 449260 4228 449316 4238
rect 449260 480 449316 4172
rect 451164 4228 451220 4238
rect 451164 480 451220 4172
rect 453068 4228 453124 4238
rect 453068 480 453124 4172
rect 454972 4228 455028 4238
rect 454972 480 455028 4172
rect 456988 4228 457044 4238
rect 456876 1876 456932 1886
rect 456876 1316 456932 1820
rect 456876 1250 456932 1260
rect 456988 480 457044 4172
rect 458780 4228 458836 4238
rect 458780 480 458836 4172
rect 460684 4228 460740 4238
rect 460684 480 460740 4172
rect 462588 3444 462644 3454
rect 462588 480 462644 3388
rect 464492 480 464548 76524
rect 553980 23604 554036 23614
rect 502572 16884 502628 16894
rect 491148 6916 491204 6926
rect 466396 4228 466452 4238
rect 466396 480 466452 4172
rect 470204 4228 470260 4238
rect 468300 3556 468356 3566
rect 468300 480 468356 3500
rect 470204 480 470260 4172
rect 472108 4228 472164 4238
rect 472108 480 472164 4172
rect 474012 4228 474068 4238
rect 474012 480 474068 4172
rect 475916 4228 475972 4238
rect 475916 480 475972 4172
rect 477820 4228 477876 4238
rect 477820 480 477876 4172
rect 479724 4228 479780 4238
rect 479724 480 479780 4172
rect 481628 4228 481684 4238
rect 481628 480 481684 4172
rect 483532 4228 483588 4238
rect 483532 480 483588 4172
rect 487340 4228 487396 4238
rect 485548 3108 485604 3118
rect 485548 480 485604 3052
rect 487340 480 487396 4172
rect 489244 4228 489300 4238
rect 489244 480 489300 4172
rect 491148 480 491204 6860
rect 493052 4228 493108 4238
rect 493052 480 493108 4172
rect 494956 4228 495012 4238
rect 494956 480 495012 4172
rect 496860 4228 496916 4238
rect 496860 480 496916 4172
rect 498764 4228 498820 4238
rect 498764 480 498820 4172
rect 500892 4228 500948 4238
rect 498988 1988 499044 1998
rect 498988 1428 499044 1932
rect 498988 1362 499044 1372
rect 500892 480 500948 4172
rect 287420 392 287672 480
rect 289324 392 289576 480
rect 291228 392 291480 480
rect 293132 392 293384 480
rect 295036 392 295288 480
rect 296940 392 297192 480
rect 298844 392 299096 480
rect 300748 392 301000 480
rect 302652 392 302904 480
rect 304556 392 304808 480
rect 306460 392 306712 480
rect 308364 392 308616 480
rect 310268 392 310520 480
rect 312172 392 312424 480
rect 285544 -960 285768 392
rect 287448 -960 287672 392
rect 289352 -960 289576 392
rect 291256 -960 291480 392
rect 293160 -960 293384 392
rect 295064 -960 295288 392
rect 296968 -960 297192 392
rect 298872 -960 299096 392
rect 300776 -960 301000 392
rect 302680 -960 302904 392
rect 304584 -960 304808 392
rect 306488 -960 306712 392
rect 308392 -960 308616 392
rect 310296 -960 310520 392
rect 312200 -960 312424 392
rect 314104 -960 314328 480
rect 315980 392 316232 480
rect 317884 392 318136 480
rect 319788 392 320040 480
rect 321692 392 321944 480
rect 323596 392 323848 480
rect 325500 392 325752 480
rect 327404 392 327656 480
rect 329308 392 329560 480
rect 331212 392 331464 480
rect 333116 392 333368 480
rect 335020 392 335272 480
rect 336924 392 337176 480
rect 338828 392 339080 480
rect 340732 392 340984 480
rect 316008 -960 316232 392
rect 317912 -960 318136 392
rect 319816 -960 320040 392
rect 321720 -960 321944 392
rect 323624 -960 323848 392
rect 325528 -960 325752 392
rect 327432 -960 327656 392
rect 329336 -960 329560 392
rect 331240 -960 331464 392
rect 333144 -960 333368 392
rect 335048 -960 335272 392
rect 336952 -960 337176 392
rect 338856 -960 339080 392
rect 340760 -960 340984 392
rect 342664 -960 342888 480
rect 344540 392 344792 480
rect 346444 392 346696 480
rect 348348 392 348600 480
rect 350252 392 350504 480
rect 352156 392 352408 480
rect 354060 392 354312 480
rect 355964 392 356216 480
rect 357868 392 358120 480
rect 359772 392 360024 480
rect 361676 392 361928 480
rect 363580 392 363832 480
rect 365484 392 365736 480
rect 367388 392 367640 480
rect 369292 392 369544 480
rect 344568 -960 344792 392
rect 346472 -960 346696 392
rect 348376 -960 348600 392
rect 350280 -960 350504 392
rect 352184 -960 352408 392
rect 354088 -960 354312 392
rect 355992 -960 356216 392
rect 357896 -960 358120 392
rect 359800 -960 360024 392
rect 361704 -960 361928 392
rect 363608 -960 363832 392
rect 365512 -960 365736 392
rect 367416 -960 367640 392
rect 369320 -960 369544 392
rect 371224 -960 371448 480
rect 373100 392 373352 480
rect 375004 392 375256 480
rect 376908 392 377160 480
rect 378812 392 379064 480
rect 380716 392 380968 480
rect 382620 392 382872 480
rect 384524 392 384776 480
rect 386428 392 386680 480
rect 388332 392 388584 480
rect 390236 392 390488 480
rect 392140 392 392392 480
rect 394044 392 394296 480
rect 395948 392 396200 480
rect 397852 392 398104 480
rect 373128 -960 373352 392
rect 375032 -960 375256 392
rect 376936 -960 377160 392
rect 378840 -960 379064 392
rect 380744 -960 380968 392
rect 382648 -960 382872 392
rect 384552 -960 384776 392
rect 386456 -960 386680 392
rect 388360 -960 388584 392
rect 390264 -960 390488 392
rect 392168 -960 392392 392
rect 394072 -960 394296 392
rect 395976 -960 396200 392
rect 397880 -960 398104 392
rect 399784 -960 400008 480
rect 401660 392 401912 480
rect 403564 392 403816 480
rect 405468 392 405720 480
rect 407372 392 407624 480
rect 409276 392 409528 480
rect 411180 392 411432 480
rect 413084 392 413336 480
rect 414988 392 415240 480
rect 416892 392 417144 480
rect 418796 392 419048 480
rect 420700 392 420952 480
rect 422604 392 422856 480
rect 424508 392 424760 480
rect 426412 392 426664 480
rect 401688 -960 401912 392
rect 403592 -960 403816 392
rect 405496 -960 405720 392
rect 407400 -960 407624 392
rect 409304 -960 409528 392
rect 411208 -960 411432 392
rect 413112 -960 413336 392
rect 415016 -960 415240 392
rect 416920 -960 417144 392
rect 418824 -960 419048 392
rect 420728 -960 420952 392
rect 422632 -960 422856 392
rect 424536 -960 424760 392
rect 426440 -960 426664 392
rect 428344 -960 428568 480
rect 430220 392 430472 480
rect 432124 392 432376 480
rect 434028 392 434280 480
rect 435932 392 436184 480
rect 437836 392 438088 480
rect 439740 392 439992 480
rect 441644 392 441896 480
rect 443548 392 443800 480
rect 445452 392 445704 480
rect 447356 392 447608 480
rect 449260 392 449512 480
rect 451164 392 451416 480
rect 453068 392 453320 480
rect 454972 392 455224 480
rect 430248 -960 430472 392
rect 432152 -960 432376 392
rect 434056 -960 434280 392
rect 435960 -960 436184 392
rect 437864 -960 438088 392
rect 439768 -960 439992 392
rect 441672 -960 441896 392
rect 443576 -960 443800 392
rect 445480 -960 445704 392
rect 447384 -960 447608 392
rect 449288 -960 449512 392
rect 451192 -960 451416 392
rect 453096 -960 453320 392
rect 455000 -960 455224 392
rect 456904 -960 457128 480
rect 458780 392 459032 480
rect 460684 392 460936 480
rect 462588 392 462840 480
rect 464492 392 464744 480
rect 466396 392 466648 480
rect 468300 392 468552 480
rect 470204 392 470456 480
rect 472108 392 472360 480
rect 474012 392 474264 480
rect 475916 392 476168 480
rect 477820 392 478072 480
rect 479724 392 479976 480
rect 481628 392 481880 480
rect 483532 392 483784 480
rect 458808 -960 459032 392
rect 460712 -960 460936 392
rect 462616 -960 462840 392
rect 464520 -960 464744 392
rect 466424 -960 466648 392
rect 468328 -960 468552 392
rect 470232 -960 470456 392
rect 472136 -960 472360 392
rect 474040 -960 474264 392
rect 475944 -960 476168 392
rect 477848 -960 478072 392
rect 479752 -960 479976 392
rect 481656 -960 481880 392
rect 483560 -960 483784 392
rect 485464 -960 485688 480
rect 487340 392 487592 480
rect 489244 392 489496 480
rect 491148 392 491400 480
rect 493052 392 493304 480
rect 494956 392 495208 480
rect 496860 392 497112 480
rect 498764 392 499016 480
rect 487368 -960 487592 392
rect 489272 -960 489496 392
rect 491176 -960 491400 392
rect 493080 -960 493304 392
rect 494984 -960 495208 392
rect 496888 -960 497112 392
rect 498792 -960 499016 392
rect 500696 392 500948 480
rect 502572 480 502628 16828
rect 546364 10948 546420 10958
rect 514108 7028 514164 7038
rect 504476 4228 504532 4238
rect 504476 480 504532 4172
rect 506380 4228 506436 4238
rect 506380 480 506436 4172
rect 508284 4228 508340 4238
rect 508284 480 508340 4172
rect 510188 4228 510244 4238
rect 510188 480 510244 4172
rect 512092 4228 512148 4238
rect 512092 480 512148 4172
rect 514108 480 514164 6972
rect 529228 5908 529284 5918
rect 515900 4228 515956 4238
rect 515900 480 515956 4172
rect 517804 4228 517860 4238
rect 517804 480 517860 4172
rect 521612 4228 521668 4238
rect 519708 1764 519764 1774
rect 519708 480 519764 1708
rect 521612 480 521668 4172
rect 523516 4228 523572 4238
rect 523516 480 523572 4172
rect 527324 4228 527380 4238
rect 524188 2100 524244 2110
rect 524188 756 524244 2044
rect 524188 690 524244 700
rect 525420 1876 525476 1886
rect 525420 480 525476 1820
rect 527324 480 527380 4172
rect 529228 480 529284 5852
rect 531132 4228 531188 4238
rect 531132 480 531188 4172
rect 533036 4228 533092 4238
rect 533036 480 533092 4172
rect 534940 4228 534996 4238
rect 534940 480 534996 4172
rect 538748 4228 538804 4238
rect 536844 1988 536900 1998
rect 536844 480 536900 1932
rect 538748 480 538804 4172
rect 540652 4228 540708 4238
rect 540652 480 540708 4172
rect 544460 4228 544516 4238
rect 542668 2100 542724 2110
rect 542668 480 542724 2044
rect 544460 480 544516 4172
rect 546364 480 546420 10892
rect 552076 6804 552132 6814
rect 550172 4228 550228 4238
rect 548268 1764 548324 1774
rect 548268 480 548324 1708
rect 550172 480 550228 4172
rect 552076 480 552132 6748
rect 553980 480 554036 23548
rect 555884 4228 555940 4238
rect 555884 480 555940 4172
rect 561596 4228 561652 4238
rect 559692 1876 559748 1886
rect 557788 1764 557844 1774
rect 557788 480 557844 1708
rect 559692 480 559748 1820
rect 561596 480 561652 4172
rect 565404 4228 565460 4238
rect 563500 3444 563556 3454
rect 563500 480 563556 3388
rect 565404 480 565460 4172
rect 567308 4228 567364 4238
rect 567308 480 567364 4172
rect 569212 480 569268 77308
rect 573020 4228 573076 4238
rect 571228 1764 571284 1774
rect 571228 480 571284 1708
rect 573020 480 573076 4172
rect 574924 4228 574980 4238
rect 574924 480 574980 4172
rect 576828 4228 576884 4238
rect 576828 480 576884 4172
rect 502572 392 502824 480
rect 504476 392 504728 480
rect 506380 392 506632 480
rect 508284 392 508536 480
rect 510188 392 510440 480
rect 512092 392 512344 480
rect 500696 -960 500920 392
rect 502600 -960 502824 392
rect 504504 -960 504728 392
rect 506408 -960 506632 392
rect 508312 -960 508536 392
rect 510216 -960 510440 392
rect 512120 -960 512344 392
rect 514024 -960 514248 480
rect 515900 392 516152 480
rect 517804 392 518056 480
rect 519708 392 519960 480
rect 521612 392 521864 480
rect 523516 392 523768 480
rect 525420 392 525672 480
rect 527324 392 527576 480
rect 529228 392 529480 480
rect 531132 392 531384 480
rect 533036 392 533288 480
rect 534940 392 535192 480
rect 536844 392 537096 480
rect 538748 392 539000 480
rect 540652 392 540904 480
rect 515928 -960 516152 392
rect 517832 -960 518056 392
rect 519736 -960 519960 392
rect 521640 -960 521864 392
rect 523544 -960 523768 392
rect 525448 -960 525672 392
rect 527352 -960 527576 392
rect 529256 -960 529480 392
rect 531160 -960 531384 392
rect 533064 -960 533288 392
rect 534968 -960 535192 392
rect 536872 -960 537096 392
rect 538776 -960 539000 392
rect 540680 -960 540904 392
rect 542584 -960 542808 480
rect 544460 392 544712 480
rect 546364 392 546616 480
rect 548268 392 548520 480
rect 550172 392 550424 480
rect 552076 392 552328 480
rect 553980 392 554232 480
rect 555884 392 556136 480
rect 557788 392 558040 480
rect 559692 392 559944 480
rect 561596 392 561848 480
rect 563500 392 563752 480
rect 565404 392 565656 480
rect 567308 392 567560 480
rect 569212 392 569464 480
rect 544488 -960 544712 392
rect 546392 -960 546616 392
rect 548296 -960 548520 392
rect 550200 -960 550424 392
rect 552104 -960 552328 392
rect 554008 -960 554232 392
rect 555912 -960 556136 392
rect 557816 -960 558040 392
rect 559720 -960 559944 392
rect 561624 -960 561848 392
rect 563528 -960 563752 392
rect 565432 -960 565656 392
rect 567336 -960 567560 392
rect 569240 -960 569464 392
rect 571144 -960 571368 480
rect 573020 392 573272 480
rect 574924 392 575176 480
rect 576828 392 577080 480
rect 573048 -960 573272 392
rect 574952 -960 575176 392
rect 576856 -960 577080 392
rect 578760 -960 578984 480
rect 580664 -960 580888 480
rect 582568 -960 582792 480
rect 584472 -960 584696 480
<< via2 >>
rect 9996 590492 10052 590548
rect 1596 583772 1652 583828
rect 1484 86492 1540 86548
rect 8316 91532 8372 91588
rect 8204 89852 8260 89908
rect 1596 38444 1652 38500
rect 3276 86604 3332 86660
rect 1484 36652 1540 36708
rect 4956 84924 5012 84980
rect 4844 83132 4900 83188
rect 4844 42924 4900 42980
rect 7980 84812 8036 84868
rect 4956 37548 5012 37604
rect 6636 73164 6692 73220
rect 3276 33964 3332 34020
rect 7980 49196 8036 49252
rect 8092 74844 8148 74900
rect 8204 43820 8260 43876
rect 9772 76412 9828 76468
rect 9660 73388 9716 73444
rect 9772 69580 9828 69636
rect 9884 73276 9940 73332
rect 9660 65548 9716 65604
rect 9884 57148 9940 57204
rect 9996 51884 10052 51940
rect 8316 41132 8372 41188
rect 8092 31276 8148 31332
rect 6636 29484 6692 29540
rect 22652 469644 22708 469700
rect 12124 103292 12180 103348
rect 12012 101612 12068 101668
rect 11676 96572 11732 96628
rect 11564 88172 11620 88228
rect 11452 73052 11508 73108
rect 11676 50092 11732 50148
rect 11564 46508 11620 46564
rect 12236 98252 12292 98308
rect 22652 73388 22708 73444
rect 34412 535724 34468 535780
rect 46172 377132 46228 377188
rect 46172 76412 46228 76468
rect 34412 73276 34468 73332
rect 33068 73164 33124 73220
rect 99260 590156 99316 590212
rect 121324 590156 121380 590212
rect 165452 590156 165508 590212
rect 187516 590156 187572 590212
rect 143388 86604 143444 86660
rect 209580 86492 209636 86548
rect 253708 583772 253764 583828
rect 297836 590156 297892 590212
rect 275772 101612 275828 101668
rect 341964 590156 342020 590212
rect 319900 91532 319956 91588
rect 231644 84924 231700 84980
rect 408268 590604 408324 590660
rect 430220 103292 430276 103348
rect 386092 89852 386148 89908
rect 496412 578732 496468 578788
rect 474348 98252 474404 98308
rect 452284 88172 452340 88228
rect 584668 590492 584724 590548
rect 562604 582092 562660 582148
rect 540540 96572 540596 96628
rect 518476 84812 518532 84868
rect 364028 83132 364084 83188
rect 129388 82460 129444 82516
rect 125580 82348 125636 82404
rect 123676 80780 123732 80836
rect 123564 78988 123620 79044
rect 77308 74844 77364 74900
rect 123452 75628 123508 75684
rect 55132 73052 55188 73108
rect 12236 48076 12292 48132
rect 12124 46284 12180 46340
rect 12012 39900 12068 39956
rect 11452 30380 11508 30436
rect 11004 28588 11060 28644
rect 123564 11004 123620 11060
rect 123452 6188 123508 6244
rect 123564 6860 123620 6916
rect 40012 3724 40068 3780
rect 40908 3724 40964 3780
rect 41356 3724 41412 3780
rect 43148 3724 43204 3780
rect 44268 3724 44324 3780
rect 44716 3724 44772 3780
rect 44940 3724 44996 3780
rect 45612 3724 45668 3780
rect 46284 3724 46340 3780
rect 46732 3724 46788 3780
rect 47628 3724 47684 3780
rect 48300 3724 48356 3780
rect 48524 3724 48580 3780
rect 48972 3724 49028 3780
rect 49196 3724 49252 3780
rect 49868 3724 49924 3780
rect 50316 3724 50372 3780
rect 50540 3724 50596 3780
rect 50988 3724 51044 3780
rect 51212 3724 51268 3780
rect 51884 3724 51940 3780
rect 52332 3724 52388 3780
rect 53228 3724 53284 3780
rect 53676 3724 53732 3780
rect 53900 3724 53956 3780
rect 54124 3724 54180 3780
rect 54348 3724 54404 3780
rect 55020 3724 55076 3780
rect 55692 3724 55748 3780
rect 55916 3724 55972 3780
rect 57036 3724 57092 3780
rect 57260 3724 57316 3780
rect 57708 3724 57764 3780
rect 57932 3724 57988 3780
rect 58604 3724 58660 3780
rect 58828 3724 58884 3780
rect 59276 3724 59332 3780
rect 59500 3724 59556 3780
rect 59724 3724 59780 3780
rect 60172 3724 60228 3780
rect 60396 3724 60452 3780
rect 60844 3724 60900 3780
rect 61068 3724 61124 3780
rect 61292 3724 61348 3780
rect 61964 3724 62020 3780
rect 63084 3724 63140 3780
rect 63980 3724 64036 3780
rect 64204 3724 64260 3780
rect 64428 3724 64484 3780
rect 64652 3724 64708 3780
rect 65324 3724 65380 3780
rect 65996 3724 66052 3780
rect 66220 3724 66276 3780
rect 67116 3724 67172 3780
rect 67788 3724 67844 3780
rect 68684 3724 68740 3780
rect 68908 3724 68964 3780
rect 69132 3724 69188 3780
rect 69356 3724 69412 3780
rect 69804 3724 69860 3780
rect 70476 3724 70532 3780
rect 71596 3724 71652 3780
rect 71820 3724 71876 3780
rect 72268 3724 72324 3780
rect 72492 3724 72548 3780
rect 72716 3724 72772 3780
rect 72940 3724 72996 3780
rect 73612 3724 73668 3780
rect 73836 3724 73892 3780
rect 74508 3724 74564 3780
rect 74956 3724 75012 3780
rect 75404 3724 75460 3780
rect 75852 3724 75908 3780
rect 76076 3724 76132 3780
rect 77196 3724 77252 3780
rect 77644 3724 77700 3780
rect 77868 3724 77924 3780
rect 79212 3724 79268 3780
rect 79884 3724 79940 3780
rect 80108 3724 80164 3780
rect 80780 3724 80836 3780
rect 81228 3724 81284 3780
rect 81900 3724 81956 3780
rect 82572 3724 82628 3780
rect 82796 3724 82852 3780
rect 83244 3724 83300 3780
rect 83692 3724 83748 3780
rect 84140 3724 84196 3780
rect 84588 3724 84644 3780
rect 85260 3724 85316 3780
rect 85932 3724 85988 3780
rect 86156 3724 86212 3780
rect 86604 3724 86660 3780
rect 86828 3724 86884 3780
rect 87276 3724 87332 3780
rect 87500 3724 87556 3780
rect 87948 3724 88004 3780
rect 88620 3724 88676 3780
rect 88844 3724 88900 3780
rect 89068 3724 89124 3780
rect 89292 3724 89348 3780
rect 89516 3724 89572 3780
rect 89964 3724 90020 3780
rect 90636 3724 90692 3780
rect 90860 3724 90916 3780
rect 91308 3724 91364 3780
rect 92204 3724 92260 3780
rect 93100 3724 93156 3780
rect 93548 3724 93604 3780
rect 94220 3724 94276 3780
rect 94892 3724 94948 3780
rect 96012 3724 96068 3780
rect 96236 3724 96292 3780
rect 96908 3724 96964 3780
rect 97356 3724 97412 3780
rect 98700 3724 98756 3780
rect 99372 3724 99428 3780
rect 99596 3724 99652 3780
rect 99820 3724 99876 3780
rect 100268 3724 100324 3780
rect 100716 3724 100772 3780
rect 100940 3724 100996 3780
rect 39564 3612 39620 3668
rect 42028 3612 42084 3668
rect 42700 3612 42756 3668
rect 62860 3612 62916 3668
rect 63532 3612 63588 3668
rect 64876 3612 64932 3668
rect 65100 3612 65156 3668
rect 65548 3612 65604 3668
rect 66668 3612 66724 3668
rect 68460 3612 68516 3668
rect 70252 3612 70308 3668
rect 71148 3612 71204 3668
rect 73388 3612 73444 3668
rect 74732 3612 74788 3668
rect 76972 3612 77028 3668
rect 78540 3612 78596 3668
rect 81452 3612 81508 3668
rect 82124 3612 82180 3668
rect 83020 3612 83076 3668
rect 83468 3612 83524 3668
rect 84812 3612 84868 3668
rect 32508 3500 32564 3556
rect 11564 3388 11620 3444
rect 15372 3052 15428 3108
rect 13356 1036 13412 1092
rect 26796 924 26852 980
rect 24892 588 24948 644
rect 17388 140 17444 196
rect 19292 252 19348 308
rect 23100 476 23156 532
rect 30604 812 30660 868
rect 28700 700 28756 756
rect 37100 3500 37156 3556
rect 46060 3500 46116 3556
rect 46956 3500 47012 3556
rect 47852 3500 47908 3556
rect 49644 3500 49700 3556
rect 51660 3500 51716 3556
rect 52780 3500 52836 3556
rect 54572 3500 54628 3556
rect 56364 3500 56420 3556
rect 58380 3500 58436 3556
rect 59052 3500 59108 3556
rect 61740 3500 61796 3556
rect 67564 3500 67620 3556
rect 76524 3500 76580 3556
rect 77420 3500 77476 3556
rect 80556 3500 80612 3556
rect 83916 3500 83972 3556
rect 104636 3500 104692 3556
rect 34636 3388 34692 3444
rect 38892 3388 38948 3444
rect 46508 3388 46564 3444
rect 47404 3388 47460 3444
rect 48748 3388 48804 3444
rect 51436 3388 51492 3444
rect 53004 3388 53060 3444
rect 70700 3388 70756 3444
rect 86380 3388 86436 3444
rect 88172 3388 88228 3444
rect 90188 3388 90244 3444
rect 91980 3388 92036 3444
rect 92876 3388 92932 3444
rect 93324 3388 93380 3444
rect 95340 3388 95396 3444
rect 96684 3388 96740 3444
rect 98028 3388 98084 3444
rect 100044 3388 100100 3444
rect 102060 3388 102116 3444
rect 43596 3276 43652 3332
rect 45836 3276 45892 3332
rect 50092 3276 50148 3332
rect 54796 3276 54852 3332
rect 56140 3276 56196 3332
rect 57484 3276 57540 3332
rect 59948 3276 60004 3332
rect 60620 3276 60676 3332
rect 63756 3276 63812 3332
rect 79436 3276 79492 3332
rect 84364 3276 84420 3332
rect 91532 3276 91588 3332
rect 93996 3276 94052 3332
rect 94668 3276 94724 3332
rect 95788 3276 95844 3332
rect 97580 3276 97636 3332
rect 40684 3164 40740 3220
rect 62636 3164 62692 3220
rect 67340 3164 67396 3220
rect 72044 3164 72100 3220
rect 73164 3164 73220 3220
rect 75180 3164 75236 3220
rect 76748 3164 76804 3220
rect 92652 3164 92708 3220
rect 95564 3164 95620 3220
rect 98252 3164 98308 3220
rect 98924 3164 98980 3220
rect 34412 1484 34468 1540
rect 35084 3052 35140 3108
rect 34860 1036 34916 1092
rect 21756 364 21812 420
rect 35420 1148 35476 1204
rect 35420 588 35476 644
rect 36204 1148 36260 1204
rect 36652 1372 36708 1428
rect 36428 924 36484 980
rect 36988 1484 37044 1540
rect 36876 812 36932 868
rect 35980 476 36036 532
rect 35756 364 35812 420
rect 35420 252 35476 308
rect 35308 140 35364 196
rect 38220 1596 38276 1652
rect 38108 1484 38164 1540
rect 38444 1372 38500 1428
rect 39116 1260 39172 1316
rect 38668 924 38724 980
rect 39788 812 39844 868
rect 39900 1484 39956 1540
rect 41132 2716 41188 2772
rect 40460 2604 40516 2660
rect 42252 3052 42308 3108
rect 41804 2828 41860 2884
rect 41580 2492 41636 2548
rect 40796 1596 40852 1652
rect 40236 1484 40292 1540
rect 39228 28 39284 84
rect 42924 2380 42980 2436
rect 43820 3052 43876 3108
rect 44044 1596 44100 1652
rect 44492 1596 44548 1652
rect 43372 1036 43428 1092
rect 43708 1372 43764 1428
rect 42476 476 42532 532
rect 47180 1372 47236 1428
rect 47516 2268 47572 2324
rect 45388 1148 45444 1204
rect 45164 476 45220 532
rect 45612 924 45668 980
rect 48076 1596 48132 1652
rect 50764 1372 50820 1428
rect 49308 924 49364 980
rect 49420 1260 49476 1316
rect 52556 1260 52612 1316
rect 53228 2268 53284 2324
rect 52108 700 52164 756
rect 53452 1596 53508 1652
rect 55244 1484 55300 1540
rect 56588 3052 56644 3108
rect 55468 924 55524 980
rect 55020 812 55076 868
rect 57148 2268 57204 2324
rect 56812 588 56868 644
rect 56924 2044 56980 2100
rect 56924 476 56980 532
rect 60956 2604 61012 2660
rect 58156 1596 58212 1652
rect 58940 2268 58996 2324
rect 62188 3052 62244 3108
rect 61516 1596 61572 1652
rect 62972 2604 63028 2660
rect 64764 2604 64820 2660
rect 62412 1484 62468 1540
rect 62748 2268 62804 2324
rect 66444 1596 66500 1652
rect 66556 2716 66612 2772
rect 65772 1484 65828 1540
rect 68012 3052 68068 3108
rect 68236 3052 68292 3108
rect 51212 28 51268 84
rect 66892 476 66948 532
rect 68572 2716 68628 2772
rect 68796 2268 68852 2324
rect 69580 1596 69636 1652
rect 70028 1596 70084 1652
rect 70364 2156 70420 2212
rect 68796 1148 68852 1204
rect 72380 2828 72436 2884
rect 71708 2716 71764 2772
rect 72156 2156 72212 2212
rect 72156 1372 72212 1428
rect 70924 1148 70980 1204
rect 74284 3052 74340 3108
rect 74060 1260 74116 1316
rect 74172 2828 74228 2884
rect 75628 2492 75684 2548
rect 76188 2716 76244 2772
rect 78092 3052 78148 3108
rect 76300 1596 76356 1652
rect 77980 2604 78036 2660
rect 78316 1372 78372 1428
rect 79100 2716 79156 2772
rect 78876 2492 78932 2548
rect 79660 1596 79716 1652
rect 79996 2828 80052 2884
rect 78876 1484 78932 1540
rect 81004 1484 81060 1540
rect 80332 1260 80388 1316
rect 81676 1260 81732 1316
rect 81788 2380 81844 2436
rect 82348 1260 82404 1316
rect 83804 2828 83860 2884
rect 85708 2604 85764 2660
rect 85484 1596 85540 1652
rect 85708 1708 85764 1764
rect 85036 1036 85092 1092
rect 87052 1484 87108 1540
rect 87500 2828 87556 2884
rect 87724 1148 87780 1204
rect 78764 252 78820 308
rect 88396 476 88452 532
rect 89404 1708 89460 1764
rect 90412 2828 90468 2884
rect 91084 2716 91140 2772
rect 89740 1484 89796 1540
rect 91308 2156 91364 2212
rect 91756 1596 91812 1652
rect 92428 812 92484 868
rect 93212 2604 93268 2660
rect 95228 2828 95284 2884
rect 95900 2828 95956 2884
rect 95116 1372 95172 1428
rect 95228 2604 95284 2660
rect 94444 1148 94500 1204
rect 93772 1036 93828 1092
rect 95676 2604 95732 2660
rect 96460 1372 96516 1428
rect 97020 2716 97076 2772
rect 95676 1260 95732 1316
rect 98476 1596 98532 1652
rect 99036 2716 99092 2772
rect 97804 1484 97860 1540
rect 97356 700 97412 756
rect 99148 1596 99204 1652
rect 102732 2268 102788 2324
rect 100492 1596 100548 1652
rect 100828 2044 100884 2100
rect 106540 3500 106596 3556
rect 108444 3500 108500 3556
rect 110348 3500 110404 3556
rect 112252 3500 112308 3556
rect 116060 3500 116116 3556
rect 114268 3388 114324 3444
rect 119868 3500 119924 3556
rect 117964 2044 118020 2100
rect 121772 3500 121828 3556
rect 123564 3164 123620 3220
rect 124012 8652 124068 8708
rect 124012 2604 124068 2660
rect 127036 16828 127092 16884
rect 127036 812 127092 868
rect 127484 4172 127540 4228
rect 315980 80668 316036 80724
rect 272188 79772 272244 79828
rect 218876 76412 218932 76468
rect 213164 73388 213220 73444
rect 205548 4396 205604 4452
rect 131292 4172 131348 4228
rect 133196 4172 133252 4228
rect 135100 4172 135156 4228
rect 138908 4172 138964 4228
rect 137004 4060 137060 4116
rect 140812 4172 140868 4228
rect 142828 4172 142884 4228
rect 144620 4172 144676 4228
rect 146524 4172 146580 4228
rect 148428 4172 148484 4228
rect 150332 4172 150388 4228
rect 152236 4172 152292 4228
rect 154140 4172 154196 4228
rect 156044 4172 156100 4228
rect 157948 4172 158004 4228
rect 161756 4172 161812 4228
rect 159852 3948 159908 4004
rect 163660 4172 163716 4228
rect 165564 4172 165620 4228
rect 167468 4172 167524 4228
rect 169372 4172 169428 4228
rect 173180 4172 173236 4228
rect 171388 3836 171444 3892
rect 175084 4172 175140 4228
rect 178892 4172 178948 4228
rect 176988 3724 177044 3780
rect 180796 4172 180852 4228
rect 184604 4172 184660 4228
rect 182700 3500 182756 3556
rect 190428 4172 190484 4228
rect 186508 1932 186564 1988
rect 188412 924 188468 980
rect 192220 4172 192276 4228
rect 196028 4172 196084 4228
rect 194124 3388 194180 3444
rect 201740 4172 201796 4228
rect 197932 1932 197988 1988
rect 203644 4172 203700 4228
rect 207452 4172 207508 4228
rect 209356 3612 209412 3668
rect 211260 588 211316 644
rect 215068 4172 215124 4228
rect 216972 4172 217028 4228
rect 230300 76300 230356 76356
rect 226492 73276 226548 73332
rect 220780 4172 220836 4228
rect 222684 4172 222740 4228
rect 224588 4172 224644 4228
rect 228508 4172 228564 4228
rect 247436 76188 247492 76244
rect 241724 74732 241780 74788
rect 232204 4172 232260 4228
rect 234108 4172 234164 4228
rect 236012 4172 236068 4228
rect 237916 4172 237972 4228
rect 239820 4172 239876 4228
rect 243628 4172 243684 4228
rect 245532 4172 245588 4228
rect 270284 74620 270340 74676
rect 249340 4172 249396 4228
rect 251244 4172 251300 4228
rect 253148 4172 253204 4228
rect 255052 4172 255108 4228
rect 258860 4172 258916 4228
rect 257068 3500 257124 3556
rect 260764 4172 260820 4228
rect 262668 4172 262724 4228
rect 264572 4172 264628 4228
rect 266476 4172 266532 4228
rect 268380 3388 268436 3444
rect 310268 78204 310324 78260
rect 281708 74508 281764 74564
rect 275996 73052 276052 73108
rect 274092 4172 274148 4228
rect 277900 72828 277956 72884
rect 279804 4172 279860 4228
rect 293132 74396 293188 74452
rect 287420 72940 287476 72996
rect 283612 4172 283668 4228
rect 285740 4172 285796 4228
rect 199724 28 199780 84
rect 289324 4172 289380 4228
rect 291228 4172 291284 4228
rect 304556 74284 304612 74340
rect 298844 72716 298900 72772
rect 295036 4172 295092 4228
rect 296940 4172 296996 4228
rect 299068 6972 299124 7028
rect 299068 1036 299124 1092
rect 300748 4172 300804 4228
rect 302652 4172 302708 4228
rect 306460 4172 306516 4228
rect 308364 3388 308420 3444
rect 312172 4172 312228 4228
rect 314188 4172 314244 4228
rect 430220 79884 430276 79940
rect 355964 79660 356020 79716
rect 321692 78092 321748 78148
rect 317884 4172 317940 4228
rect 319788 4172 319844 4228
rect 327404 77980 327460 78036
rect 323596 4172 323652 4228
rect 325500 4172 325556 4228
rect 329308 77868 329364 77924
rect 350252 77756 350308 77812
rect 333116 76076 333172 76132
rect 331212 4172 331268 4228
rect 344540 75964 344596 76020
rect 335020 74172 335076 74228
rect 338828 73500 338884 73556
rect 336924 4172 336980 4228
rect 340732 4172 340788 4228
rect 342748 4172 342804 4228
rect 346444 4172 346500 4228
rect 348348 4172 348404 4228
rect 352156 4172 352212 4228
rect 354060 4172 354116 4228
rect 361676 79548 361732 79604
rect 357868 75852 357924 75908
rect 359772 4172 359828 4228
rect 369292 79436 369348 79492
rect 367388 74060 367444 74116
rect 363580 4172 363636 4228
rect 365484 4172 365540 4228
rect 373100 79324 373156 79380
rect 371308 4172 371364 4228
rect 378812 79212 378868 79268
rect 375004 4172 375060 4228
rect 376908 4172 376964 4228
rect 413084 79100 413140 79156
rect 390236 77644 390292 77700
rect 380716 4172 380772 4228
rect 384524 4172 384580 4228
rect 382620 1820 382676 1876
rect 386428 4172 386484 4228
rect 388332 4172 388388 4228
rect 401660 75740 401716 75796
rect 399868 8652 399924 8708
rect 392140 4172 392196 4228
rect 394044 4172 394100 4228
rect 395948 4172 396004 4228
rect 397852 4172 397908 4228
rect 403564 4172 403620 4228
rect 407372 4172 407428 4228
rect 405468 1708 405524 1764
rect 411180 4172 411236 4228
rect 409276 3388 409332 3444
rect 424508 77532 424564 77588
rect 418796 74844 418852 74900
rect 416892 4172 416948 4228
rect 414988 3388 415044 3444
rect 420700 4172 420756 4228
rect 422604 4172 422660 4228
rect 426412 4172 426468 4228
rect 428428 4172 428484 4228
rect 426748 1708 426804 1764
rect 426748 1148 426804 1204
rect 441644 77420 441700 77476
rect 434028 11004 434084 11060
rect 432124 4172 432180 4228
rect 435932 4172 435988 4228
rect 437836 4172 437892 4228
rect 439740 4172 439796 4228
rect 569212 77308 569268 77364
rect 464492 76524 464548 76580
rect 443548 4172 443604 4228
rect 447356 4172 447412 4228
rect 445452 2492 445508 2548
rect 449260 4172 449316 4228
rect 451164 4172 451220 4228
rect 453068 4172 453124 4228
rect 454972 4172 455028 4228
rect 456988 4172 457044 4228
rect 456876 1820 456932 1876
rect 456876 1260 456932 1316
rect 458780 4172 458836 4228
rect 460684 4172 460740 4228
rect 462588 3388 462644 3444
rect 553980 23548 554036 23604
rect 502572 16828 502628 16884
rect 491148 6860 491204 6916
rect 466396 4172 466452 4228
rect 470204 4172 470260 4228
rect 468300 3500 468356 3556
rect 472108 4172 472164 4228
rect 474012 4172 474068 4228
rect 475916 4172 475972 4228
rect 477820 4172 477876 4228
rect 479724 4172 479780 4228
rect 481628 4172 481684 4228
rect 483532 4172 483588 4228
rect 487340 4172 487396 4228
rect 485548 3052 485604 3108
rect 489244 4172 489300 4228
rect 493052 4172 493108 4228
rect 494956 4172 495012 4228
rect 496860 4172 496916 4228
rect 498764 4172 498820 4228
rect 500892 4172 500948 4228
rect 498988 1932 499044 1988
rect 498988 1372 499044 1428
rect 546364 10892 546420 10948
rect 514108 6972 514164 7028
rect 504476 4172 504532 4228
rect 506380 4172 506436 4228
rect 508284 4172 508340 4228
rect 510188 4172 510244 4228
rect 512092 4172 512148 4228
rect 529228 5852 529284 5908
rect 515900 4172 515956 4228
rect 517804 4172 517860 4228
rect 521612 4172 521668 4228
rect 519708 1708 519764 1764
rect 523516 4172 523572 4228
rect 527324 4172 527380 4228
rect 524188 2044 524244 2100
rect 524188 700 524244 756
rect 525420 1820 525476 1876
rect 531132 4172 531188 4228
rect 533036 4172 533092 4228
rect 534940 4172 534996 4228
rect 538748 4172 538804 4228
rect 536844 1932 536900 1988
rect 540652 4172 540708 4228
rect 544460 4172 544516 4228
rect 542668 2044 542724 2100
rect 552076 6748 552132 6804
rect 550172 4172 550228 4228
rect 548268 1708 548324 1764
rect 555884 4172 555940 4228
rect 561596 4172 561652 4228
rect 559692 1820 559748 1876
rect 557788 1708 557844 1764
rect 565404 4172 565460 4228
rect 563500 3388 563556 3444
rect 567308 4172 567364 4228
rect 573020 4172 573076 4228
rect 571228 1708 571284 1764
rect 574924 4172 574980 4228
rect 576828 4172 576884 4228
<< metal3 >>
rect 27682 590604 27692 590660
rect 27748 590604 408268 590660
rect 408324 590604 408334 590660
rect 9986 590492 9996 590548
rect 10052 590492 584668 590548
rect 584724 590492 584734 590548
rect 99222 590156 99260 590212
rect 99316 590156 99326 590212
rect 120978 590156 120988 590212
rect 121044 590156 121324 590212
rect 121380 590156 121390 590212
rect 164658 590156 164668 590212
rect 164724 590156 165452 590212
rect 165508 590156 165518 590212
rect 186498 590156 186508 590212
rect 186564 590156 187516 590212
rect 187572 590156 187582 590212
rect 297378 590156 297388 590212
rect 297444 590156 297836 590212
rect 297892 590156 297902 590212
rect 341058 590156 341068 590212
rect 341124 590156 341964 590212
rect 342020 590156 342030 590212
rect 595560 588644 597000 588840
rect 26002 588588 26012 588644
rect 26068 588616 597000 588644
rect 26068 588588 595672 588616
rect -960 587188 480 587384
rect -960 587160 3388 587188
rect 392 587132 3388 587160
rect 3444 587132 3454 587188
rect 1586 583772 1596 583828
rect 1652 583772 253708 583828
rect 253764 583772 253774 583828
rect 22642 582092 22652 582148
rect 22708 582092 562604 582148
rect 562660 582092 562670 582148
rect 19282 578732 19292 578788
rect 19348 578732 496412 578788
rect 496468 578732 496478 578788
rect 595560 575428 597000 575624
rect 17602 575372 17612 575428
rect 17668 575400 597000 575428
rect 17668 575372 595672 575400
rect -960 573076 480 573272
rect -960 573048 12012 573076
rect 392 573020 12012 573048
rect 12068 573020 12078 573076
rect 595560 562212 597000 562408
rect 590706 562156 590716 562212
rect 590772 562184 597000 562212
rect 590772 562156 595672 562184
rect -960 558964 480 559160
rect -960 558936 10892 558964
rect 392 558908 10892 558936
rect 10948 558908 10958 558964
rect 595560 548996 597000 549192
rect 24322 548940 24332 548996
rect 24388 548968 597000 548996
rect 24388 548940 595672 548968
rect -960 544852 480 545048
rect -960 544824 532 544852
rect 392 544796 532 544824
rect 476 544740 532 544796
rect 18 544684 28 544740
rect 84 544684 532 544740
rect 595560 535780 597000 535976
rect 34402 535724 34412 535780
rect 34468 535752 597000 535780
rect 34468 535724 595672 535752
rect -960 530740 480 530936
rect -960 530712 15148 530740
rect 392 530684 15148 530712
rect 15204 530684 15214 530740
rect 3154 523292 3164 523348
rect 3220 523292 590716 523348
rect 590772 523292 590782 523348
rect 595560 522564 597000 522760
rect 590482 522508 590492 522564
rect 590548 522536 597000 522564
rect 590548 522508 595672 522536
rect -960 516628 480 516824
rect -960 516600 11900 516628
rect 392 516572 11900 516600
rect 11956 516572 11966 516628
rect 595560 509348 597000 509544
rect 14242 509292 14252 509348
rect 14308 509320 597000 509348
rect 14308 509292 595672 509320
rect -960 502516 480 502712
rect -960 502488 2492 502516
rect 392 502460 2492 502488
rect 2548 502460 2558 502516
rect 595560 496132 597000 496328
rect 590146 496076 590156 496132
rect 590212 496104 597000 496132
rect 590212 496076 595672 496104
rect 31042 494732 31052 494788
rect 31108 494732 590156 494788
rect 590212 494732 590222 494788
rect -960 488404 480 488600
rect -960 488376 13468 488404
rect 392 488348 13468 488376
rect 13524 488348 13534 488404
rect 595560 482916 597000 483112
rect 8306 482860 8316 482916
rect 8372 482888 597000 482916
rect 8372 482860 595672 482888
rect -960 474292 480 474488
rect -960 474264 532 474292
rect 392 474236 532 474264
rect 476 474180 532 474236
rect 130 474124 140 474180
rect 196 474124 532 474180
rect 595560 469700 597000 469896
rect 22642 469644 22652 469700
rect 22708 469672 597000 469700
rect 22708 469644 595672 469672
rect -960 460180 480 460376
rect -960 460152 7532 460180
rect 392 460124 7532 460152
rect 7588 460124 7598 460180
rect 595560 456484 597000 456680
rect 20962 456428 20972 456484
rect 21028 456456 597000 456484
rect 21028 456428 595672 456456
rect -960 446068 480 446264
rect -960 446040 4620 446068
rect 392 446012 4620 446040
rect 4676 446012 4686 446068
rect 595560 443268 597000 443464
rect 86482 443212 86492 443268
rect 86548 443240 597000 443268
rect 86548 443212 595672 443240
rect -960 431956 480 432152
rect -960 431928 4172 431956
rect 392 431900 4172 431928
rect 4228 431900 4238 431956
rect 595560 430164 597000 430248
rect 11666 430108 11676 430164
rect 11732 430108 597000 430164
rect 595560 430024 597000 430108
rect -960 417844 480 418040
rect -960 417816 532 417844
rect 392 417788 532 417816
rect 476 417732 532 417788
rect 242 417676 252 417732
rect 308 417676 532 417732
rect 595560 416836 597000 417032
rect 76402 416780 76412 416836
rect 76468 416808 597000 416836
rect 76468 416780 595672 416808
rect -960 403732 480 403928
rect -960 403704 13580 403732
rect 392 403676 13580 403704
rect 13636 403676 13646 403732
rect 595560 403620 597000 403816
rect 8194 403564 8204 403620
rect 8260 403592 597000 403620
rect 8260 403564 595672 403592
rect 595560 390404 597000 390600
rect 29362 390348 29372 390404
rect 29428 390376 597000 390404
rect 29428 390348 595672 390376
rect -960 389620 480 389816
rect -960 389592 4284 389620
rect 392 389564 4284 389592
rect 4340 389564 4350 389620
rect 595560 377188 597000 377384
rect 46162 377132 46172 377188
rect 46228 377160 597000 377188
rect 46228 377132 595672 377160
rect -960 375508 480 375704
rect -960 375480 2604 375508
rect 392 375452 2604 375480
rect 2660 375452 2670 375508
rect 595560 363972 597000 364168
rect 587122 363916 587132 363972
rect 587188 363944 597000 363972
rect 587188 363916 595672 363944
rect -960 361396 480 361592
rect -960 361368 4732 361396
rect 392 361340 4732 361368
rect 4788 361340 4798 361396
rect 595560 350756 597000 350952
rect 15922 350700 15932 350756
rect 15988 350728 597000 350756
rect 15988 350700 595672 350728
rect -960 347284 480 347480
rect -960 347256 2716 347284
rect 392 347228 2716 347256
rect 2772 347228 2782 347284
rect 595560 337540 597000 337736
rect 21074 337484 21084 337540
rect 21140 337512 597000 337540
rect 21140 337484 595672 337512
rect -960 333172 480 333368
rect -960 333144 588 333172
rect 392 333116 588 333144
rect 644 333116 654 333172
rect 595560 324324 597000 324520
rect 47842 324268 47852 324324
rect 47908 324296 597000 324324
rect 47908 324268 595672 324296
rect -960 319060 480 319256
rect -960 319032 11788 319060
rect 392 319004 11788 319032
rect 11844 319004 11854 319060
rect 595560 311108 597000 311304
rect 126802 311052 126812 311108
rect 126868 311080 597000 311108
rect 126868 311052 595672 311080
rect -960 304948 480 305144
rect -960 304920 4396 304948
rect 392 304892 4396 304920
rect 4452 304892 4462 304948
rect 4610 304108 4620 304164
rect 4676 304108 11004 304164
rect 11060 304108 11070 304164
rect 595560 297892 597000 298088
rect 590146 297836 590156 297892
rect 590212 297864 597000 297892
rect 590212 297836 595672 297864
rect 150322 296492 150332 296548
rect 150388 296492 590156 296548
rect 590212 296492 590222 296548
rect -960 290836 480 291032
rect -960 290808 7644 290836
rect 392 290780 7644 290808
rect 7700 290780 7710 290836
rect 595560 284676 597000 284872
rect 173842 284620 173852 284676
rect 173908 284648 597000 284676
rect 173908 284620 595672 284648
rect -960 276724 480 276920
rect -960 276696 4508 276724
rect 392 276668 4508 276696
rect 4564 276668 4574 276724
rect 4722 275548 4732 275604
rect 4788 275548 6188 275604
rect 6244 275548 6254 275604
rect 595560 271460 597000 271656
rect 145282 271404 145292 271460
rect 145348 271432 597000 271460
rect 145348 271404 595672 271432
rect -960 262612 480 262808
rect -960 262584 4620 262612
rect 392 262556 4620 262584
rect 4676 262556 4686 262612
rect 595560 258244 597000 258440
rect 126914 258188 126924 258244
rect 126980 258216 597000 258244
rect 126980 258188 595672 258216
rect -960 248472 480 248696
rect 595560 245028 597000 245224
rect 591266 244972 591276 245028
rect 591332 245000 597000 245028
rect 591332 244972 595672 245000
rect 136882 242732 136892 242788
rect 136948 242732 591276 242788
rect 591332 242732 591342 242788
rect -960 234360 480 234584
rect 595560 231924 597000 232008
rect 148642 231868 148652 231924
rect 148708 231868 597000 231924
rect 595560 231784 597000 231868
rect -960 220248 480 220472
rect 595560 218596 597000 218792
rect 127026 218540 127036 218596
rect 127092 218568 597000 218596
rect 127092 218540 595672 218568
rect -960 206136 480 206360
rect 595560 205380 597000 205576
rect 135202 205324 135212 205380
rect 135268 205352 597000 205380
rect 135268 205324 595672 205352
rect -960 192024 480 192248
rect 595560 192164 597000 192360
rect 141922 192108 141932 192164
rect 141988 192136 597000 192164
rect 141988 192108 595672 192136
rect 595560 178948 597000 179144
rect 127138 178892 127148 178948
rect 127204 178920 597000 178948
rect 127204 178892 595672 178920
rect -960 177912 480 178136
rect 595560 165732 597000 165928
rect 590146 165676 590156 165732
rect 590212 165704 597000 165732
rect 590212 165676 595672 165704
rect -960 163800 480 164024
rect 133522 163772 133532 163828
rect 133588 163772 590156 163828
rect 590212 163772 590222 163828
rect 595560 152516 597000 152712
rect 140242 152460 140252 152516
rect 140308 152488 597000 152516
rect 140308 152460 595672 152488
rect -960 149688 480 149912
rect 595560 139300 597000 139496
rect 127250 139244 127260 139300
rect 127316 139272 597000 139300
rect 127316 139244 595672 139272
rect -960 135576 480 135800
rect 595560 126084 597000 126280
rect 129042 126028 129052 126084
rect 129108 126056 597000 126084
rect 129108 126028 595672 126056
rect -960 121464 480 121688
rect 595560 112868 597000 113064
rect 138562 112812 138572 112868
rect 138628 112840 597000 112868
rect 138628 112812 595672 112840
rect -960 107352 480 107576
rect 8642 104972 8652 105028
rect 8708 104972 587132 105028
rect 587188 104972 587198 105028
rect 12114 103292 12124 103348
rect 12180 103292 430220 103348
rect 430276 103292 430286 103348
rect 12002 101612 12012 101668
rect 12068 101612 275772 101668
rect 275828 101612 275838 101668
rect 595560 99652 597000 99848
rect 590146 99596 590156 99652
rect 590212 99624 597000 99652
rect 590212 99596 595672 99624
rect 12226 98252 12236 98308
rect 12292 98252 474348 98308
rect 474404 98252 474414 98308
rect 474562 98252 474572 98308
rect 474628 98252 590156 98308
rect 590212 98252 590222 98308
rect 11666 96572 11676 96628
rect 11732 96572 540540 96628
rect 540596 96572 540606 96628
rect -960 93240 480 93464
rect 8306 91532 8316 91588
rect 8372 91532 319900 91588
rect 319956 91532 319966 91588
rect 8194 89852 8204 89908
rect 8260 89852 386092 89908
rect 386148 89852 386158 89908
rect 11554 88172 11564 88228
rect 11620 88172 452284 88228
rect 452340 88172 452350 88228
rect 3266 86604 3276 86660
rect 3332 86604 143388 86660
rect 143444 86604 143454 86660
rect 1474 86492 1484 86548
rect 1540 86492 209580 86548
rect 209636 86492 209646 86548
rect 595560 86436 597000 86632
rect 504802 86380 504812 86436
rect 504868 86408 597000 86436
rect 504868 86380 595672 86408
rect 4946 84924 4956 84980
rect 5012 84924 231644 84980
rect 231700 84924 231710 84980
rect 7970 84812 7980 84868
rect 8036 84812 518476 84868
rect 518532 84812 518542 84868
rect 4834 83132 4844 83188
rect 4900 83132 364028 83188
rect 364084 83132 364094 83188
rect 46946 82684 46956 82740
rect 47012 82684 114268 82740
rect 114324 82684 114334 82740
rect 47618 82572 47628 82628
rect 47684 82572 121100 82628
rect 121156 82572 121166 82628
rect 48514 82460 48524 82516
rect 48580 82460 129388 82516
rect 129444 82460 129454 82516
rect 43586 82348 43596 82404
rect 43652 82348 125580 82404
rect 125636 82348 125646 82404
rect 9874 81452 9884 81508
rect 9940 81452 47852 81508
rect 47908 81452 47918 81508
rect 46834 81004 46844 81060
rect 46900 81004 110908 81060
rect 110964 81004 110974 81060
rect 48290 80892 48300 80948
rect 48356 80892 119308 80948
rect 119364 80892 119374 80948
rect 48402 80780 48412 80836
rect 48468 80780 123676 80836
rect 123732 80780 123742 80836
rect 70354 80668 70364 80724
rect 70420 80668 315980 80724
rect 316036 80668 316046 80724
rect 84802 79884 84812 79940
rect 84868 79884 430220 79940
rect 430276 79884 430286 79940
rect 65426 79772 65436 79828
rect 65492 79772 272188 79828
rect 272244 79772 272254 79828
rect 76514 79660 76524 79716
rect 76580 79660 355964 79716
rect 356020 79660 356030 79716
rect 75842 79548 75852 79604
rect 75908 79548 361676 79604
rect 361732 79548 361742 79604
rect 81554 79436 81564 79492
rect 81620 79436 369292 79492
rect 369348 79436 369358 79492
rect -960 79128 480 79352
rect 78306 79324 78316 79380
rect 78372 79324 373100 79380
rect 373156 79324 373166 79380
rect 78866 79212 78876 79268
rect 78932 79212 378812 79268
rect 378868 79212 378878 79268
rect 81778 79100 81788 79156
rect 81844 79100 413084 79156
rect 413140 79100 413150 79156
rect 99036 78988 123564 79044
rect 123620 78988 123630 79044
rect 99036 78372 99092 78988
rect 86594 78316 86604 78372
rect 86660 78316 99092 78372
rect 70242 78204 70252 78260
rect 70308 78204 310268 78260
rect 310324 78204 310334 78260
rect 71698 78092 71708 78148
rect 71764 78092 321692 78148
rect 321748 78092 321758 78148
rect 76626 77980 76636 78036
rect 76692 77980 327404 78036
rect 327460 77980 327470 78036
rect 73042 77868 73052 77924
rect 73108 77868 329308 77924
rect 329364 77868 329374 77924
rect 74498 77756 74508 77812
rect 74564 77756 350252 77812
rect 350308 77756 350318 77812
rect 79426 77644 79436 77700
rect 79492 77644 390236 77700
rect 390292 77644 390302 77700
rect 83010 77532 83020 77588
rect 83076 77532 424508 77588
rect 424564 77532 424574 77588
rect 85586 77420 85596 77476
rect 85652 77420 441644 77476
rect 441700 77420 441710 77476
rect 100146 77308 100156 77364
rect 100212 77308 569212 77364
rect 569268 77308 569278 77364
rect 87938 76524 87948 76580
rect 88004 76524 464492 76580
rect 464548 76524 464558 76580
rect 9762 76412 9772 76468
rect 9828 76412 46172 76468
rect 46228 76412 46238 76468
rect 60274 76412 60284 76468
rect 60340 76412 218876 76468
rect 218932 76412 218942 76468
rect 60386 76300 60396 76356
rect 60452 76300 230300 76356
rect 230356 76300 230366 76356
rect 52770 76188 52780 76244
rect 52836 76188 247436 76244
rect 247492 76188 247502 76244
rect 72482 76076 72492 76132
rect 72548 76076 333116 76132
rect 333172 76076 333182 76132
rect 73826 75964 73836 76020
rect 73892 75964 344540 76020
rect 344596 75964 344606 76020
rect 75394 75852 75404 75908
rect 75460 75852 357868 75908
rect 357924 75852 357934 75908
rect 81442 75740 81452 75796
rect 81508 75740 401660 75796
rect 401716 75740 401726 75796
rect 94434 75628 94444 75684
rect 94500 75628 123452 75684
rect 123508 75628 123518 75684
rect 8082 74844 8092 74900
rect 8148 74844 77308 74900
rect 77364 74844 77374 74900
rect 82562 74844 82572 74900
rect 82628 74844 418796 74900
rect 418852 74844 418862 74900
rect 9986 74732 9996 74788
rect 10052 74732 21084 74788
rect 21140 74732 21150 74788
rect 62066 74732 62076 74788
rect 62132 74732 241724 74788
rect 241780 74732 241790 74788
rect 65314 74620 65324 74676
rect 65380 74620 270284 74676
rect 270340 74620 270350 74676
rect 61954 74508 61964 74564
rect 62020 74508 281708 74564
rect 281764 74508 281774 74564
rect 67778 74396 67788 74452
rect 67844 74396 293132 74452
rect 293188 74396 293198 74452
rect 69122 74284 69132 74340
rect 69188 74284 304556 74340
rect 304612 74284 304622 74340
rect 72706 74172 72716 74228
rect 72772 74172 335020 74228
rect 335076 74172 335086 74228
rect 77074 74060 77084 74116
rect 77140 74060 367388 74116
rect 367444 74060 367454 74116
rect 8754 73948 8764 74004
rect 8820 73948 11788 74004
rect 11844 73948 11854 74004
rect 91522 73948 91532 74004
rect 91588 73948 121772 74004
rect 121828 73948 121838 74004
rect 74722 73500 74732 73556
rect 74788 73500 338828 73556
rect 338884 73500 338894 73556
rect 9650 73388 9660 73444
rect 9716 73388 22652 73444
rect 22708 73388 22718 73444
rect 57474 73388 57484 73444
rect 57540 73388 213164 73444
rect 213220 73388 213230 73444
rect 9874 73276 9884 73332
rect 9940 73276 34412 73332
rect 34468 73276 34478 73332
rect 58482 73276 58492 73332
rect 58548 73276 226492 73332
rect 226548 73276 226558 73332
rect 595560 73220 597000 73416
rect 6626 73164 6636 73220
rect 6692 73164 33068 73220
rect 33124 73164 33134 73220
rect 130162 73164 130172 73220
rect 130228 73192 597000 73220
rect 130228 73164 595672 73192
rect 11442 73052 11452 73108
rect 11508 73052 55132 73108
rect 55188 73052 55198 73108
rect 58034 73052 58044 73108
rect 58100 73052 275996 73108
rect 276052 73052 276062 73108
rect 8530 72940 8540 72996
rect 8596 72940 13580 72996
rect 13636 72940 13646 72996
rect 66658 72940 66668 72996
rect 66724 72940 287420 72996
rect 287476 72940 287486 72996
rect 56354 72828 56364 72884
rect 56420 72828 277900 72884
rect 277956 72828 277966 72884
rect 68786 72716 68796 72772
rect 68852 72716 298844 72772
rect 298900 72716 298910 72772
rect 123928 72492 126812 72548
rect 126868 72492 126878 72548
rect 9874 70700 9884 70756
rect 9940 70700 12040 70756
rect 9986 69804 9996 69860
rect 10052 69804 12040 69860
rect 9762 69580 9772 69636
rect 9828 69580 9996 69636
rect 10052 69580 10062 69636
rect 123928 69580 150332 69636
rect 150388 69580 150398 69636
rect 12674 68908 12684 68964
rect 12740 68908 12750 68964
rect 8642 68012 8652 68068
rect 8708 68012 12040 68068
rect 9986 67116 9996 67172
rect 10052 67116 12040 67172
rect 12562 66892 12572 66948
rect 12628 66892 12638 66948
rect 12572 66248 12628 66892
rect 123928 66668 173852 66724
rect 173908 66668 173918 66724
rect 9650 65548 9660 65604
rect 9716 65548 9996 65604
rect 10052 65548 10062 65604
rect 8194 65324 8204 65380
rect 8260 65324 12040 65380
rect -960 65016 480 65240
rect 12450 64988 12460 65044
rect 12516 64988 12526 65044
rect 12460 64456 12516 64988
rect 123928 63756 145292 63812
rect 145348 63756 145358 63812
rect 11330 63532 11340 63588
rect 11396 63532 12040 63588
rect 12450 63308 12460 63364
rect 12516 63308 12526 63364
rect 12460 62664 12516 63308
rect 12674 61740 12684 61796
rect 12740 61740 12750 61796
rect 9986 60844 9996 60900
rect 10052 60844 12040 60900
rect 123928 60844 126924 60900
rect 126980 60844 126990 60900
rect 595560 60004 597000 60200
rect 8306 59948 8316 60004
rect 8372 59948 12040 60004
rect 126802 59948 126812 60004
rect 126868 59976 597000 60004
rect 126868 59948 595672 59976
rect 12450 59612 12460 59668
rect 12516 59612 12526 59668
rect 12460 59080 12516 59612
rect 12562 58716 12572 58772
rect 12628 58716 12638 58772
rect 12572 58184 12628 58716
rect 123928 57932 136892 57988
rect 136948 57932 136958 57988
rect 11442 57260 11452 57316
rect 11508 57260 12040 57316
rect 9874 57148 9884 57204
rect 9940 57148 9950 57204
rect 9884 57092 9940 57148
rect 9884 57036 12068 57092
rect 12012 56392 12068 57036
rect 12338 56140 12348 56196
rect 12404 56140 12414 56196
rect 12348 55496 12404 56140
rect 123928 55020 148652 55076
rect 148708 55020 148718 55076
rect 3154 54572 3164 54628
rect 3220 54572 12040 54628
rect 12674 53676 12684 53732
rect 12740 53676 12750 53732
rect 12338 53452 12348 53508
rect 12404 53452 12414 53508
rect 12348 52808 12404 53452
rect 123928 52108 127036 52164
rect 127092 52108 127102 52164
rect 9986 51884 9996 51940
rect 10052 51884 12040 51940
rect 12338 51660 12348 51716
rect 12404 51660 12414 51716
rect -960 50904 480 51128
rect 12348 51016 12404 51660
rect 11666 50092 11676 50148
rect 11732 50092 12040 50148
rect 7970 49196 7980 49252
rect 8036 49196 12040 49252
rect 123928 49196 135212 49252
rect 135268 49196 135278 49252
rect 12674 48300 12684 48356
rect 12740 48300 12750 48356
rect 12226 48076 12236 48132
rect 12292 48076 12302 48132
rect 12236 47432 12292 48076
rect 127586 47852 127596 47908
rect 127652 47852 141932 47908
rect 141988 47852 141998 47908
rect 595560 46788 597000 46984
rect 590482 46732 590492 46788
rect 590548 46760 597000 46788
rect 590548 46732 595672 46760
rect 11554 46508 11564 46564
rect 11620 46508 12040 46564
rect 12114 46284 12124 46340
rect 12180 46284 12190 46340
rect 123928 46284 127596 46340
rect 127652 46284 127662 46340
rect 12124 45640 12180 46284
rect 9986 44716 9996 44772
rect 10052 44716 12040 44772
rect 8194 43820 8204 43876
rect 8260 43820 12040 43876
rect 123928 43372 127148 43428
rect 127204 43372 127214 43428
rect 4834 42924 4844 42980
rect 4900 42924 12040 42980
rect 6514 42028 6524 42084
rect 6580 42028 12040 42084
rect 8306 41132 8316 41188
rect 8372 41132 12040 41188
rect 123928 40460 133532 40516
rect 133588 40460 133598 40516
rect 6626 40236 6636 40292
rect 6692 40236 12040 40292
rect 12002 39900 12012 39956
rect 12068 39900 12078 39956
rect 12012 39368 12068 39900
rect 1586 38444 1596 38500
rect 1652 38444 12040 38500
rect 4946 37548 4956 37604
rect 5012 37548 12040 37604
rect 123928 37548 140252 37604
rect 140308 37548 140318 37604
rect -960 36792 480 37016
rect 1474 36652 1484 36708
rect 1540 36652 12040 36708
rect 11554 35756 11564 35812
rect 11620 35756 12040 35812
rect 7970 34860 7980 34916
rect 8036 34860 12040 34916
rect 123928 34636 127260 34692
rect 127316 34636 127326 34692
rect 3266 33964 3276 34020
rect 3332 33964 12040 34020
rect 595560 33684 597000 33768
rect 127026 33628 127036 33684
rect 127092 33628 597000 33684
rect 4610 33516 4620 33572
rect 4676 33516 7756 33572
rect 7812 33516 7822 33572
rect 595560 33544 597000 33628
rect 8082 33068 8092 33124
rect 8148 33068 12040 33124
rect 127362 32732 127372 32788
rect 127428 32732 504812 32788
rect 504868 32732 504878 32788
rect 3042 32172 3052 32228
rect 3108 32172 12040 32228
rect 127138 31948 127148 32004
rect 127204 31948 587132 32004
rect 587188 31948 587198 32004
rect 123928 31724 129052 31780
rect 129108 31724 129118 31780
rect 8082 31276 8092 31332
rect 8148 31276 12040 31332
rect 127250 31052 127260 31108
rect 127316 31052 590492 31108
rect 590548 31052 590558 31108
rect 11442 30380 11452 30436
rect 11508 30380 12040 30436
rect 126914 30380 126924 30436
rect 126980 30380 137788 30436
rect 137732 30324 137788 30380
rect 127474 30268 127484 30324
rect 127540 30268 130172 30324
rect 130228 30268 130238 30324
rect 137732 30268 575372 30324
rect 575428 30268 575438 30324
rect 6626 29484 6636 29540
rect 6692 29484 12040 29540
rect 123928 28812 138572 28868
rect 138628 28812 138638 28868
rect 10994 28588 11004 28644
rect 11060 28588 12040 28644
rect 3266 27692 3276 27748
rect 3332 27692 12040 27748
rect 12002 26796 12012 26852
rect 12068 26796 12078 26852
rect 10882 25900 10892 25956
rect 10948 25900 12040 25956
rect 123928 25900 474572 25956
rect 474628 25900 474638 25956
rect 18 25004 28 25060
rect 84 25004 12040 25060
rect 8978 24108 8988 24164
rect 9044 24108 12040 24164
rect 130162 23548 130172 23604
rect 130228 23548 553980 23604
rect 554036 23548 554046 23604
rect 12002 23212 12012 23268
rect 12068 23212 12078 23268
rect 123928 22988 127372 23044
rect 127428 22988 127438 23044
rect -960 22680 480 22904
rect 2482 22316 2492 22372
rect 2548 22316 12040 22372
rect 8866 21420 8876 21476
rect 8932 21420 12040 21476
rect 130 20524 140 20580
rect 196 20524 12040 20580
rect 587122 20524 587132 20580
rect 587188 20552 595672 20580
rect 587188 20524 597000 20552
rect 595560 20328 597000 20524
rect 123928 20076 127484 20132
rect 127540 20076 127550 20132
rect 7522 19628 7532 19684
rect 7588 19628 12040 19684
rect 10994 18732 11004 18788
rect 11060 18732 12040 18788
rect 4162 17836 4172 17892
rect 4228 17836 12040 17892
rect 123928 17164 126812 17220
rect 126868 17164 126878 17220
rect 242 16940 252 16996
rect 308 16940 12040 16996
rect 127026 16828 127036 16884
rect 127092 16828 502572 16884
rect 502628 16828 502638 16884
rect 8530 16044 8540 16100
rect 8596 16044 12040 16100
rect 4274 15148 4284 15204
rect 4340 15148 12040 15204
rect 2594 14252 2604 14308
rect 2660 14252 12040 14308
rect 123928 14252 127260 14308
rect 127316 14252 127326 14308
rect 6178 13356 6188 13412
rect 6244 13356 12040 13412
rect 2706 12460 2716 12516
rect 2772 12460 12040 12516
rect 354 11564 364 11620
rect 420 11564 12040 11620
rect 123928 11340 127036 11396
rect 127092 11340 127102 11396
rect 123554 11004 123564 11060
rect 123620 11004 434028 11060
rect 434084 11004 434094 11060
rect 124002 10892 124012 10948
rect 124068 10892 546364 10948
rect 546420 10892 546430 10948
rect 8754 10668 8764 10724
rect 8820 10668 12040 10724
rect 4386 9772 4396 9828
rect 4452 9772 12040 9828
rect 7634 8876 7644 8932
rect 7700 8876 12040 8932
rect -960 8568 480 8792
rect 124002 8652 124012 8708
rect 124068 8652 399868 8708
rect 399924 8652 399934 8708
rect 123928 8428 127148 8484
rect 127204 8428 127214 8484
rect 4498 7980 4508 8036
rect 4564 7980 12040 8036
rect 595560 7140 597000 7336
rect 7746 7084 7756 7140
rect 7812 7084 12040 7140
rect 575362 7084 575372 7140
rect 575428 7112 597000 7140
rect 575428 7084 595672 7112
rect 299058 6972 299068 7028
rect 299124 6972 514108 7028
rect 514164 6972 514174 7028
rect 123554 6860 123564 6916
rect 123620 6860 491148 6916
rect 491204 6860 491214 6916
rect 123442 6748 123452 6804
rect 123508 6748 552076 6804
rect 552132 6748 552142 6804
rect 123442 6188 123452 6244
rect 123508 6188 123518 6244
rect 123452 5908 123508 6188
rect 123452 5852 529228 5908
rect 529284 5852 529294 5908
rect 123928 5516 126924 5572
rect 126980 5516 126990 5572
rect 75058 4508 75068 4564
rect 75124 4508 76524 4564
rect 76580 4508 76590 4564
rect 79538 4508 79548 4564
rect 79604 4508 80668 4564
rect 80724 4508 80734 4564
rect 85698 4508 85708 4564
rect 85764 4508 93324 4564
rect 93380 4508 93390 4564
rect 57586 4396 57596 4452
rect 57652 4396 205548 4452
rect 205604 4396 205614 4452
rect 62850 4284 62860 4340
rect 62916 4284 79828 4340
rect 84690 4284 84700 4340
rect 84756 4284 91420 4340
rect 91476 4284 91486 4340
rect 92754 4284 92764 4340
rect 92820 4284 93436 4340
rect 93492 4284 93502 4340
rect 79772 4228 79828 4284
rect 40684 4172 57148 4228
rect 57204 4172 57214 4228
rect 61180 4172 61628 4228
rect 61684 4172 61694 4228
rect 62178 4172 62188 4228
rect 62244 4172 73948 4228
rect 79762 4172 79772 4228
rect 79828 4172 79838 4228
rect 82114 4172 82124 4228
rect 82180 4172 120988 4228
rect 121044 4172 121054 4228
rect 126018 4172 126028 4228
rect 126084 4172 127484 4228
rect 127540 4172 127550 4228
rect 131254 4172 131292 4228
rect 131348 4172 131358 4228
rect 132738 4172 132748 4228
rect 132804 4172 133196 4228
rect 133252 4172 133262 4228
rect 134418 4172 134428 4228
rect 134484 4172 135100 4228
rect 135156 4172 135166 4228
rect 137778 4172 137788 4228
rect 137844 4172 138908 4228
rect 138964 4172 138974 4228
rect 139458 4172 139468 4228
rect 139524 4172 140812 4228
rect 140868 4172 140878 4228
rect 142790 4172 142828 4228
rect 142884 4172 142894 4228
rect 144582 4172 144620 4228
rect 144676 4172 144686 4228
rect 146178 4172 146188 4228
rect 146244 4172 146524 4228
rect 146580 4172 146590 4228
rect 147858 4172 147868 4228
rect 147924 4172 148428 4228
rect 148484 4172 148494 4228
rect 149538 4172 149548 4228
rect 149604 4172 150332 4228
rect 150388 4172 150398 4228
rect 151218 4172 151228 4228
rect 151284 4172 152236 4228
rect 152292 4172 152302 4228
rect 152898 4172 152908 4228
rect 152964 4172 154140 4228
rect 154196 4172 154206 4228
rect 154578 4172 154588 4228
rect 154644 4172 156044 4228
rect 156100 4172 156110 4228
rect 157910 4172 157948 4228
rect 158004 4172 158014 4228
rect 161298 4172 161308 4228
rect 161364 4172 161756 4228
rect 161812 4172 161822 4228
rect 163622 4172 163660 4228
rect 163716 4172 163726 4228
rect 164658 4172 164668 4228
rect 164724 4172 165564 4228
rect 165620 4172 165630 4228
rect 166338 4172 166348 4228
rect 166404 4172 167468 4228
rect 167524 4172 167534 4228
rect 169334 4172 169372 4228
rect 169428 4172 169438 4228
rect 173142 4172 173180 4228
rect 173236 4172 173246 4228
rect 174738 4172 174748 4228
rect 174804 4172 175084 4228
rect 175140 4172 175150 4228
rect 178098 4172 178108 4228
rect 178164 4172 178892 4228
rect 178948 4172 178958 4228
rect 179778 4172 179788 4228
rect 179844 4172 180796 4228
rect 180852 4172 180862 4228
rect 183138 4172 183148 4228
rect 183204 4172 184604 4228
rect 184660 4172 184670 4228
rect 190390 4172 190428 4228
rect 190484 4172 190494 4228
rect 191538 4172 191548 4228
rect 191604 4172 192220 4228
rect 192276 4172 192286 4228
rect 194898 4172 194908 4228
rect 194964 4172 196028 4228
rect 196084 4172 196094 4228
rect 201702 4172 201740 4228
rect 201796 4172 201806 4228
rect 203606 4172 203644 4228
rect 203700 4172 203710 4228
rect 206658 4172 206668 4228
rect 206724 4172 207452 4228
rect 207508 4172 207518 4228
rect 215030 4172 215068 4228
rect 215124 4172 215134 4228
rect 216934 4172 216972 4228
rect 217028 4172 217038 4228
rect 220098 4172 220108 4228
rect 220164 4172 220780 4228
rect 220836 4172 220846 4228
rect 221778 4172 221788 4228
rect 221844 4172 222684 4228
rect 222740 4172 222750 4228
rect 223458 4172 223468 4228
rect 223524 4172 224588 4228
rect 224644 4172 224654 4228
rect 228470 4172 228508 4228
rect 228564 4172 228574 4228
rect 231858 4172 231868 4228
rect 231924 4172 232204 4228
rect 232260 4172 232270 4228
rect 233538 4172 233548 4228
rect 233604 4172 234108 4228
rect 234164 4172 234174 4228
rect 235218 4172 235228 4228
rect 235284 4172 236012 4228
rect 236068 4172 236078 4228
rect 236898 4172 236908 4228
rect 236964 4172 237916 4228
rect 237972 4172 237982 4228
rect 238578 4172 238588 4228
rect 238644 4172 239820 4228
rect 239876 4172 239886 4228
rect 243618 4172 243628 4228
rect 243684 4172 243722 4228
rect 245494 4172 245532 4228
rect 245588 4172 245598 4228
rect 248658 4172 248668 4228
rect 248724 4172 249340 4228
rect 249396 4172 249406 4228
rect 250338 4172 250348 4228
rect 250404 4172 251244 4228
rect 251300 4172 251310 4228
rect 252018 4172 252028 4228
rect 252084 4172 253148 4228
rect 253204 4172 253214 4228
rect 253698 4172 253708 4228
rect 253764 4172 255052 4228
rect 255108 4172 255118 4228
rect 258822 4172 258860 4228
rect 258916 4172 258926 4228
rect 260418 4172 260428 4228
rect 260484 4172 260764 4228
rect 260820 4172 260830 4228
rect 262098 4172 262108 4228
rect 262164 4172 262668 4228
rect 262724 4172 262734 4228
rect 263778 4172 263788 4228
rect 263844 4172 264572 4228
rect 264628 4172 264638 4228
rect 265458 4172 265468 4228
rect 265524 4172 266476 4228
rect 266532 4172 266542 4228
rect 274054 4172 274092 4228
rect 274148 4172 274158 4228
rect 278898 4172 278908 4228
rect 278964 4172 279804 4228
rect 279860 4172 279870 4228
rect 282594 4172 282604 4228
rect 282660 4172 283612 4228
rect 283668 4172 283678 4228
rect 285730 4172 285740 4228
rect 285796 4172 286300 4228
rect 286356 4172 286366 4228
rect 288978 4172 288988 4228
rect 289044 4172 289324 4228
rect 289380 4172 289390 4228
rect 290658 4172 290668 4228
rect 290724 4172 291228 4228
rect 291284 4172 291294 4228
rect 294018 4172 294028 4228
rect 294084 4172 295036 4228
rect 295092 4172 295102 4228
rect 295698 4172 295708 4228
rect 295764 4172 296940 4228
rect 296996 4172 297006 4228
rect 300710 4172 300748 4228
rect 300804 4172 300814 4228
rect 302614 4172 302652 4228
rect 302708 4172 302718 4228
rect 305778 4172 305788 4228
rect 305844 4172 306460 4228
rect 306516 4172 306526 4228
rect 310818 4172 310828 4228
rect 310884 4172 312172 4228
rect 312228 4172 312238 4228
rect 314178 4172 314188 4228
rect 314244 4172 314282 4228
rect 317538 4172 317548 4228
rect 317604 4172 317884 4228
rect 317940 4172 317950 4228
rect 319218 4172 319228 4228
rect 319284 4172 319788 4228
rect 319844 4172 319854 4228
rect 322578 4172 322588 4228
rect 322644 4172 323596 4228
rect 323652 4172 323662 4228
rect 324258 4172 324268 4228
rect 324324 4172 325500 4228
rect 325556 4172 325566 4228
rect 331174 4172 331212 4228
rect 331268 4172 331278 4228
rect 336018 4172 336028 4228
rect 336084 4172 336924 4228
rect 336980 4172 336990 4228
rect 339378 4172 339388 4228
rect 339444 4172 340732 4228
rect 340788 4172 340798 4228
rect 342710 4172 342748 4228
rect 342804 4172 342814 4228
rect 346098 4172 346108 4228
rect 346164 4172 346444 4228
rect 346500 4172 346510 4228
rect 347778 4172 347788 4228
rect 347844 4172 348348 4228
rect 348404 4172 348414 4228
rect 351138 4172 351148 4228
rect 351204 4172 352156 4228
rect 352212 4172 352222 4228
rect 352818 4172 352828 4228
rect 352884 4172 354060 4228
rect 354116 4172 354126 4228
rect 359734 4172 359772 4228
rect 359828 4172 359838 4228
rect 362898 4172 362908 4228
rect 362964 4172 363580 4228
rect 363636 4172 363646 4228
rect 364578 4172 364588 4228
rect 364644 4172 365484 4228
rect 365540 4172 365550 4228
rect 371270 4172 371308 4228
rect 371364 4172 371374 4228
rect 374966 4172 375004 4228
rect 375060 4172 375070 4228
rect 376338 4172 376348 4228
rect 376404 4172 376908 4228
rect 376964 4172 376974 4228
rect 379698 4172 379708 4228
rect 379764 4172 380716 4228
rect 380772 4172 380782 4228
rect 383058 4172 383068 4228
rect 383124 4172 384524 4228
rect 384580 4172 384590 4228
rect 386390 4172 386428 4228
rect 386484 4172 386494 4228
rect 388294 4172 388332 4228
rect 388388 4172 388398 4228
rect 391458 4172 391468 4228
rect 391524 4172 392140 4228
rect 392196 4172 392206 4228
rect 393138 4172 393148 4228
rect 393204 4172 394044 4228
rect 394100 4172 394110 4228
rect 394818 4172 394828 4228
rect 394884 4172 395948 4228
rect 396004 4172 396014 4228
rect 396498 4172 396508 4228
rect 396564 4172 397852 4228
rect 397908 4172 397918 4228
rect 403218 4172 403228 4228
rect 403284 4172 403564 4228
rect 403620 4172 403630 4228
rect 406578 4172 406588 4228
rect 406644 4172 407372 4228
rect 407428 4172 407438 4228
rect 409938 4172 409948 4228
rect 410004 4172 411180 4228
rect 411236 4172 411246 4228
rect 416854 4172 416892 4228
rect 416948 4172 416958 4228
rect 420018 4172 420028 4228
rect 420084 4172 420700 4228
rect 420756 4172 420766 4228
rect 422566 4172 422604 4228
rect 422660 4172 422670 4228
rect 425058 4172 425068 4228
rect 425124 4172 426412 4228
rect 426468 4172 426478 4228
rect 428390 4172 428428 4228
rect 428484 4172 428494 4228
rect 431778 4172 431788 4228
rect 431844 4172 432124 4228
rect 432180 4172 432190 4228
rect 435138 4172 435148 4228
rect 435204 4172 435932 4228
rect 435988 4172 435998 4228
rect 436818 4172 436828 4228
rect 436884 4172 437836 4228
rect 437892 4172 437902 4228
rect 438498 4172 438508 4228
rect 438564 4172 439740 4228
rect 439796 4172 439806 4228
rect 443538 4172 443548 4228
rect 443604 4172 443642 4228
rect 446898 4172 446908 4228
rect 446964 4172 447356 4228
rect 447412 4172 447422 4228
rect 448578 4172 448588 4228
rect 448644 4172 449260 4228
rect 449316 4172 449326 4228
rect 450258 4172 450268 4228
rect 450324 4172 451164 4228
rect 451220 4172 451230 4228
rect 451938 4172 451948 4228
rect 452004 4172 453068 4228
rect 453124 4172 453134 4228
rect 453618 4172 453628 4228
rect 453684 4172 454972 4228
rect 455028 4172 455038 4228
rect 456950 4172 456988 4228
rect 457044 4172 457054 4228
rect 458742 4172 458780 4228
rect 458836 4172 458846 4228
rect 460338 4172 460348 4228
rect 460404 4172 460684 4228
rect 460740 4172 460750 4228
rect 465378 4172 465388 4228
rect 465444 4172 466396 4228
rect 466452 4172 466462 4228
rect 468738 4172 468748 4228
rect 468804 4172 470204 4228
rect 470260 4172 470270 4228
rect 472070 4172 472108 4228
rect 472164 4172 472174 4228
rect 473974 4172 474012 4228
rect 474068 4172 474078 4228
rect 475458 4172 475468 4228
rect 475524 4172 475916 4228
rect 475972 4172 475982 4228
rect 477138 4172 477148 4228
rect 477204 4172 477820 4228
rect 477876 4172 477886 4228
rect 478818 4172 478828 4228
rect 478884 4172 479724 4228
rect 479780 4172 479790 4228
rect 480498 4172 480508 4228
rect 480564 4172 481628 4228
rect 481684 4172 481694 4228
rect 482178 4172 482188 4228
rect 482244 4172 483532 4228
rect 483588 4172 483598 4228
rect 487302 4172 487340 4228
rect 487396 4172 487406 4228
rect 488898 4172 488908 4228
rect 488964 4172 489244 4228
rect 489300 4172 489310 4228
rect 492258 4172 492268 4228
rect 492324 4172 493052 4228
rect 493108 4172 493118 4228
rect 493938 4172 493948 4228
rect 494004 4172 494956 4228
rect 495012 4172 495022 4228
rect 495618 4172 495628 4228
rect 495684 4172 496860 4228
rect 496916 4172 496926 4228
rect 497634 4172 497644 4228
rect 497700 4172 498764 4228
rect 498820 4172 498830 4228
rect 500882 4172 500892 4228
rect 500948 4172 501340 4228
rect 501396 4172 501406 4228
rect 504018 4172 504028 4228
rect 504084 4172 504476 4228
rect 504532 4172 504542 4228
rect 505698 4172 505708 4228
rect 505764 4172 506380 4228
rect 506436 4172 506446 4228
rect 508246 4172 508284 4228
rect 508340 4172 508350 4228
rect 509058 4172 509068 4228
rect 509124 4172 510188 4228
rect 510244 4172 510254 4228
rect 510738 4172 510748 4228
rect 510804 4172 512092 4228
rect 512148 4172 512158 4228
rect 515862 4172 515900 4228
rect 515956 4172 515966 4228
rect 517458 4172 517468 4228
rect 517524 4172 517804 4228
rect 517860 4172 517870 4228
rect 520818 4172 520828 4228
rect 520884 4172 521612 4228
rect 521668 4172 521678 4228
rect 522498 4172 522508 4228
rect 522564 4172 523516 4228
rect 523572 4172 523582 4228
rect 525858 4172 525868 4228
rect 525924 4172 527324 4228
rect 527380 4172 527390 4228
rect 531094 4172 531132 4228
rect 531188 4172 531198 4228
rect 532578 4172 532588 4228
rect 532644 4172 533036 4228
rect 533092 4172 533102 4228
rect 534258 4172 534268 4228
rect 534324 4172 534940 4228
rect 534996 4172 535006 4228
rect 537618 4172 537628 4228
rect 537684 4172 538748 4228
rect 538804 4172 538814 4228
rect 539298 4172 539308 4228
rect 539364 4172 540652 4228
rect 540708 4172 540718 4228
rect 544422 4172 544460 4228
rect 544516 4172 544526 4228
rect 549378 4172 549388 4228
rect 549444 4172 550172 4228
rect 550228 4172 550238 4228
rect 554418 4172 554428 4228
rect 554484 4172 555884 4228
rect 555940 4172 555950 4228
rect 561138 4172 561148 4228
rect 561204 4172 561596 4228
rect 561652 4172 561662 4228
rect 564498 4172 564508 4228
rect 564564 4172 565404 4228
rect 565460 4172 565470 4228
rect 566178 4172 566188 4228
rect 566244 4172 567308 4228
rect 567364 4172 567374 4228
rect 572982 4172 573020 4228
rect 573076 4172 573086 4228
rect 574578 4172 574588 4228
rect 574644 4172 574924 4228
rect 574980 4172 574990 4228
rect 576258 4172 576268 4228
rect 576324 4172 576828 4228
rect 576884 4172 576894 4228
rect 40684 3780 40740 4172
rect 61180 4116 61236 4172
rect 73892 4116 73948 4172
rect 41132 4060 53116 4116
rect 53172 4060 53182 4116
rect 54114 4060 54124 4116
rect 54180 4060 61236 4116
rect 61292 4060 68124 4116
rect 68180 4060 68190 4116
rect 68898 4060 68908 4116
rect 68964 4060 70140 4116
rect 70196 4060 70206 4116
rect 72258 4060 72268 4116
rect 72324 4060 73724 4116
rect 73780 4060 73790 4116
rect 73892 4060 137004 4116
rect 137060 4060 137070 4116
rect 40002 3724 40012 3780
rect 40068 3724 40740 3780
rect 40870 3724 40908 3780
rect 40964 3724 40974 3780
rect 41132 3668 41188 4060
rect 61292 4004 61348 4060
rect 42140 3948 61348 4004
rect 61404 3948 74172 4004
rect 74228 3948 74238 4004
rect 79538 3948 79548 4004
rect 79604 3948 79614 4004
rect 91410 3948 91420 4004
rect 91476 3948 159852 4004
rect 159908 3948 159918 4004
rect 42140 3780 42196 3948
rect 61404 3892 61460 3948
rect 79548 3892 79604 3948
rect 41346 3724 41356 3780
rect 41412 3724 42196 3780
rect 42252 3836 61460 3892
rect 61618 3836 61628 3892
rect 61684 3836 79604 3892
rect 79884 3836 79996 3892
rect 80052 3836 80062 3892
rect 80658 3836 80668 3892
rect 80724 3836 85708 3892
rect 42252 3668 42308 3836
rect 79884 3780 79940 3836
rect 43110 3724 43148 3780
rect 43204 3724 43214 3780
rect 44230 3724 44268 3780
rect 44324 3724 44334 3780
rect 44678 3724 44716 3780
rect 44772 3724 44782 3780
rect 44930 3724 44940 3780
rect 44996 3724 45034 3780
rect 45574 3724 45612 3780
rect 45668 3724 45678 3780
rect 46274 3724 46284 3780
rect 46340 3724 46508 3780
rect 46564 3724 46574 3780
rect 46722 3724 46732 3780
rect 46788 3724 46844 3780
rect 46900 3724 46910 3780
rect 47590 3724 47628 3780
rect 47684 3724 47694 3780
rect 48178 3724 48188 3780
rect 48244 3724 48300 3780
rect 48356 3724 48366 3780
rect 48486 3724 48524 3780
rect 48580 3724 48590 3780
rect 48934 3724 48972 3780
rect 49028 3724 49038 3780
rect 49186 3724 49196 3780
rect 49252 3724 49290 3780
rect 49830 3724 49868 3780
rect 49924 3724 49934 3780
rect 50278 3724 50316 3780
rect 50372 3724 50382 3780
rect 50530 3724 50540 3780
rect 50596 3724 50634 3780
rect 50950 3724 50988 3780
rect 51044 3724 51054 3780
rect 51202 3724 51212 3780
rect 51268 3724 51306 3780
rect 51762 3724 51772 3780
rect 51828 3724 51884 3780
rect 51940 3724 51950 3780
rect 52294 3724 52332 3780
rect 52388 3724 52398 3780
rect 53190 3724 53228 3780
rect 53284 3724 53294 3780
rect 53442 3724 53452 3780
rect 53508 3724 53676 3780
rect 53732 3724 53742 3780
rect 53862 3724 53900 3780
rect 53956 3724 53966 3780
rect 54114 3724 54124 3780
rect 54180 3724 54218 3780
rect 54310 3724 54348 3780
rect 54404 3724 54414 3780
rect 55010 3724 55020 3780
rect 55076 3724 55244 3780
rect 55300 3724 55310 3780
rect 55654 3724 55692 3780
rect 55748 3724 55758 3780
rect 55906 3724 55916 3780
rect 55972 3724 56700 3780
rect 56756 3724 56766 3780
rect 56914 3724 56924 3780
rect 56980 3724 57036 3780
rect 57092 3724 57102 3780
rect 57222 3724 57260 3780
rect 57316 3724 57326 3780
rect 57670 3724 57708 3780
rect 57764 3724 57774 3780
rect 57922 3724 57932 3780
rect 57988 3724 58026 3780
rect 58370 3724 58380 3780
rect 58436 3724 58604 3780
rect 58660 3724 58670 3780
rect 58818 3724 58828 3780
rect 58884 3724 59052 3780
rect 59108 3724 59118 3780
rect 59238 3724 59276 3780
rect 59332 3724 59342 3780
rect 59490 3724 59500 3780
rect 59556 3724 59594 3780
rect 59714 3724 59724 3780
rect 59780 3724 59818 3780
rect 60134 3724 60172 3780
rect 60228 3724 60238 3780
rect 60358 3724 60396 3780
rect 60452 3724 60462 3780
rect 60806 3724 60844 3780
rect 60900 3724 60910 3780
rect 61030 3724 61068 3780
rect 61124 3724 61134 3780
rect 61282 3724 61292 3780
rect 61348 3724 61386 3780
rect 61730 3724 61740 3780
rect 61796 3724 61964 3780
rect 62020 3724 62030 3780
rect 62132 3724 62860 3780
rect 62916 3724 62926 3780
rect 63074 3724 63084 3780
rect 63140 3724 63644 3780
rect 63700 3724 63710 3780
rect 63942 3724 63980 3780
rect 64036 3724 64046 3780
rect 64194 3724 64204 3780
rect 64260 3724 64298 3780
rect 64390 3724 64428 3780
rect 64484 3724 64494 3780
rect 64642 3724 64652 3780
rect 64708 3724 65100 3780
rect 65156 3724 65166 3780
rect 65314 3724 65324 3780
rect 65380 3724 65436 3780
rect 65492 3724 65502 3780
rect 65958 3724 65996 3780
rect 66052 3724 66062 3780
rect 66210 3724 66220 3780
rect 66276 3724 66332 3780
rect 66388 3724 66398 3780
rect 66658 3724 66668 3780
rect 66724 3724 67116 3780
rect 67172 3724 67182 3780
rect 67750 3724 67788 3780
rect 67844 3724 67854 3780
rect 68450 3724 68460 3780
rect 68516 3724 68684 3780
rect 68740 3724 68750 3780
rect 68898 3724 68908 3780
rect 68964 3724 69002 3780
rect 69094 3724 69132 3780
rect 69188 3724 69198 3780
rect 69346 3724 69356 3780
rect 69412 3724 69468 3780
rect 69524 3724 69534 3780
rect 69794 3724 69804 3780
rect 69860 3724 70140 3780
rect 70196 3724 70206 3780
rect 70354 3724 70364 3780
rect 70420 3724 70476 3780
rect 70532 3724 70542 3780
rect 71558 3724 71596 3780
rect 71652 3724 71662 3780
rect 71810 3724 71820 3780
rect 71876 3724 71932 3780
rect 71988 3724 71998 3780
rect 72230 3724 72268 3780
rect 72324 3724 72334 3780
rect 72454 3724 72492 3780
rect 72548 3724 72558 3780
rect 72706 3724 72716 3780
rect 72772 3724 72810 3780
rect 72930 3724 72940 3780
rect 72996 3724 73164 3780
rect 73220 3724 73230 3780
rect 73490 3724 73500 3780
rect 73556 3724 73612 3780
rect 73668 3724 73678 3780
rect 73798 3724 73836 3780
rect 73892 3724 73902 3780
rect 74470 3724 74508 3780
rect 74564 3724 74574 3780
rect 74946 3724 74956 3780
rect 75012 3724 75180 3780
rect 75236 3724 75246 3780
rect 75366 3724 75404 3780
rect 75460 3724 75470 3780
rect 75814 3724 75852 3780
rect 75908 3724 75918 3780
rect 76066 3724 76076 3780
rect 76132 3724 76170 3780
rect 76962 3724 76972 3780
rect 77028 3724 77196 3780
rect 77252 3724 77262 3780
rect 77606 3724 77644 3780
rect 77700 3724 77710 3780
rect 77858 3724 77868 3780
rect 77924 3724 78876 3780
rect 78932 3724 78942 3780
rect 79202 3724 79212 3780
rect 79268 3724 79436 3780
rect 79492 3724 79502 3780
rect 79874 3724 79884 3780
rect 79940 3724 79950 3780
rect 80098 3724 80108 3780
rect 80164 3724 80556 3780
rect 80612 3724 80622 3780
rect 80742 3724 80780 3780
rect 80836 3724 80846 3780
rect 81190 3724 81228 3780
rect 81284 3724 81294 3780
rect 81890 3724 81900 3780
rect 81956 3724 82012 3780
rect 82068 3724 82078 3780
rect 82534 3724 82572 3780
rect 82628 3724 82638 3780
rect 82786 3724 82796 3780
rect 82852 3724 82890 3780
rect 83010 3724 83020 3780
rect 83076 3724 83244 3780
rect 83300 3724 83310 3780
rect 83654 3724 83692 3780
rect 83748 3724 83758 3780
rect 84102 3724 84140 3780
rect 84196 3724 84206 3780
rect 84550 3724 84588 3780
rect 84644 3724 84654 3780
rect 85250 3724 85260 3780
rect 85316 3724 85484 3780
rect 85540 3724 85550 3780
rect 62132 3668 62188 3724
rect 85652 3668 85708 3836
rect 86604 3836 87276 3892
rect 87332 3836 87342 3892
rect 88620 3836 88956 3892
rect 89012 3836 89022 3892
rect 92978 3836 92988 3892
rect 93044 3836 93156 3892
rect 93314 3836 93324 3892
rect 93380 3836 171388 3892
rect 171444 3836 171454 3892
rect 86604 3780 86660 3836
rect 88620 3780 88676 3836
rect 93100 3780 93156 3836
rect 85894 3724 85932 3780
rect 85988 3724 85998 3780
rect 86146 3724 86156 3780
rect 86212 3724 86250 3780
rect 86594 3724 86604 3780
rect 86660 3724 86670 3780
rect 86790 3724 86828 3780
rect 86884 3724 86894 3780
rect 87154 3724 87164 3780
rect 87220 3724 87276 3780
rect 87332 3724 87342 3780
rect 87490 3724 87500 3780
rect 87556 3724 87724 3780
rect 87780 3724 87790 3780
rect 87910 3724 87948 3780
rect 88004 3724 88014 3780
rect 88610 3724 88620 3780
rect 88676 3724 88686 3780
rect 88806 3724 88844 3780
rect 88900 3724 88910 3780
rect 89058 3724 89068 3780
rect 89124 3724 89162 3780
rect 89254 3724 89292 3780
rect 89348 3724 89358 3780
rect 89506 3724 89516 3780
rect 89572 3724 89610 3780
rect 89730 3724 89740 3780
rect 89796 3724 89964 3780
rect 90020 3724 90030 3780
rect 90402 3724 90412 3780
rect 90468 3724 90636 3780
rect 90692 3724 90702 3780
rect 90822 3724 90860 3780
rect 90916 3724 90926 3780
rect 91270 3724 91308 3780
rect 91364 3724 91374 3780
rect 92082 3724 92092 3780
rect 92148 3724 92204 3780
rect 92260 3724 92270 3780
rect 93090 3724 93100 3780
rect 93156 3724 93166 3780
rect 93538 3724 93548 3780
rect 93604 3724 93660 3780
rect 93716 3724 93726 3780
rect 94182 3724 94220 3780
rect 94276 3724 94286 3780
rect 94882 3724 94892 3780
rect 94948 3724 95452 3780
rect 95508 3724 95518 3780
rect 95974 3724 96012 3780
rect 96068 3724 96078 3780
rect 96226 3724 96236 3780
rect 96292 3724 96330 3780
rect 96450 3724 96460 3780
rect 96516 3724 96908 3780
rect 96964 3724 96974 3780
rect 97234 3724 97244 3780
rect 97300 3724 97356 3780
rect 97412 3724 97422 3780
rect 98578 3724 98588 3780
rect 98644 3724 98700 3780
rect 98756 3724 98766 3780
rect 99334 3724 99372 3780
rect 99428 3724 99438 3780
rect 99586 3724 99596 3780
rect 99652 3724 99690 3780
rect 99782 3724 99820 3780
rect 99876 3724 99886 3780
rect 100146 3724 100156 3780
rect 100212 3724 100268 3780
rect 100324 3724 100334 3780
rect 100594 3724 100604 3780
rect 100660 3724 100716 3780
rect 100772 3724 100782 3780
rect 100930 3724 100940 3780
rect 100996 3724 102396 3780
rect 102452 3724 102462 3780
rect 108332 3724 176988 3780
rect 177044 3724 177054 3780
rect 108332 3668 108388 3724
rect 39554 3612 39564 3668
rect 39620 3612 41188 3668
rect 42018 3612 42028 3668
rect 42084 3612 42308 3668
rect 42690 3612 42700 3668
rect 42756 3612 62188 3668
rect 62850 3612 62860 3668
rect 62916 3612 63308 3668
rect 63364 3612 63374 3668
rect 63522 3612 63532 3668
rect 63588 3612 63756 3668
rect 63812 3612 63822 3668
rect 64838 3612 64876 3668
rect 64932 3612 64942 3668
rect 65090 3612 65100 3668
rect 65156 3612 65324 3668
rect 65380 3612 65390 3668
rect 65538 3612 65548 3668
rect 65604 3612 66220 3668
rect 66276 3612 66286 3668
rect 66434 3612 66444 3668
rect 66500 3612 66668 3668
rect 66724 3612 66734 3668
rect 68450 3612 68460 3668
rect 68516 3612 68796 3668
rect 68852 3612 68862 3668
rect 69906 3612 69916 3668
rect 69972 3612 70252 3668
rect 70308 3612 70318 3668
rect 71138 3612 71148 3668
rect 71204 3612 71708 3668
rect 71764 3612 71774 3668
rect 71932 3612 72324 3668
rect 73378 3612 73388 3668
rect 73444 3612 73612 3668
rect 73668 3612 73678 3668
rect 74722 3612 74732 3668
rect 74788 3612 75292 3668
rect 75348 3612 75358 3668
rect 76738 3612 76748 3668
rect 76804 3612 76972 3668
rect 77028 3612 77038 3668
rect 78530 3612 78540 3668
rect 78596 3612 80108 3668
rect 80164 3612 80174 3668
rect 81442 3612 81452 3668
rect 81508 3612 81900 3668
rect 81956 3612 81966 3668
rect 82086 3612 82124 3668
rect 82180 3612 82190 3668
rect 82898 3612 82908 3668
rect 82964 3612 83020 3668
rect 83076 3612 83086 3668
rect 83458 3612 83468 3668
rect 83524 3612 83804 3668
rect 83860 3612 83870 3668
rect 84802 3612 84812 3668
rect 84868 3612 85372 3668
rect 85428 3612 85438 3668
rect 85652 3612 108388 3668
rect 108668 3612 126028 3668
rect 209318 3612 209356 3668
rect 209412 3612 209422 3668
rect 71932 3556 71988 3612
rect 32498 3500 32508 3556
rect 32564 3500 37100 3556
rect 37156 3500 37166 3556
rect 46050 3500 46060 3556
rect 46116 3500 46396 3556
rect 46452 3500 46462 3556
rect 46722 3500 46732 3556
rect 46788 3500 46956 3556
rect 47012 3500 47022 3556
rect 47842 3500 47852 3556
rect 47908 3500 48412 3556
rect 48468 3500 48478 3556
rect 49634 3500 49644 3556
rect 49700 3500 50204 3556
rect 50260 3500 50270 3556
rect 51650 3500 51660 3556
rect 51716 3500 51996 3556
rect 52052 3500 52062 3556
rect 52770 3500 52780 3556
rect 52836 3500 53564 3556
rect 53620 3500 53630 3556
rect 54562 3500 54572 3556
rect 54628 3500 55356 3556
rect 55412 3500 55422 3556
rect 55570 3500 55580 3556
rect 55636 3500 56364 3556
rect 56420 3500 56430 3556
rect 57474 3500 57484 3556
rect 57540 3500 58380 3556
rect 58436 3500 58446 3556
rect 59042 3500 59052 3556
rect 59108 3500 60284 3556
rect 60340 3500 60350 3556
rect 61730 3500 61740 3556
rect 61796 3500 62076 3556
rect 62132 3500 62142 3556
rect 67554 3500 67564 3556
rect 67620 3500 68572 3556
rect 68628 3500 68638 3556
rect 68796 3500 71988 3556
rect 68796 3444 68852 3500
rect 72268 3444 72324 3612
rect 76514 3500 76524 3556
rect 76580 3500 77084 3556
rect 77140 3500 77150 3556
rect 77410 3500 77420 3556
rect 77476 3500 79884 3556
rect 79940 3500 79950 3556
rect 80546 3500 80556 3556
rect 80612 3500 81452 3556
rect 81508 3500 81518 3556
rect 83906 3500 83916 3556
rect 83972 3500 84812 3556
rect 84868 3500 84878 3556
rect 85652 3500 102508 3556
rect 104178 3500 104188 3556
rect 104244 3500 104636 3556
rect 104692 3500 104702 3556
rect 106502 3500 106540 3556
rect 106596 3500 106606 3556
rect 107538 3500 107548 3556
rect 107604 3500 108444 3556
rect 108500 3500 108510 3556
rect 85652 3444 85708 3500
rect 102452 3444 102508 3500
rect 108668 3444 108724 3612
rect 125972 3556 126028 3612
rect 109218 3500 109228 3556
rect 109284 3500 110348 3556
rect 110404 3500 110414 3556
rect 110898 3500 110908 3556
rect 110964 3500 112252 3556
rect 112308 3500 112318 3556
rect 116022 3500 116060 3556
rect 116116 3500 116126 3556
rect 119298 3500 119308 3556
rect 119364 3500 119868 3556
rect 119924 3500 119934 3556
rect 121090 3500 121100 3556
rect 121156 3500 121772 3556
rect 121828 3500 121838 3556
rect 125972 3500 182700 3556
rect 182756 3500 182766 3556
rect 257030 3500 257068 3556
rect 257124 3500 257134 3556
rect 468262 3500 468300 3556
rect 468356 3500 468366 3556
rect 11554 3388 11564 3444
rect 11620 3388 34636 3444
rect 34692 3388 34702 3444
rect 38882 3388 38892 3444
rect 38948 3388 46284 3444
rect 46340 3388 46350 3444
rect 46498 3388 46508 3444
rect 46564 3388 46956 3444
rect 47012 3388 47022 3444
rect 47394 3388 47404 3444
rect 47460 3388 48300 3444
rect 48356 3388 48366 3444
rect 48738 3388 48748 3444
rect 48804 3388 50092 3444
rect 50148 3388 50158 3444
rect 51426 3388 51436 3444
rect 51492 3388 51884 3444
rect 51940 3388 51950 3444
rect 52994 3388 53004 3444
rect 53060 3388 54572 3444
rect 54628 3388 54638 3444
rect 55412 3388 68852 3444
rect 70690 3388 70700 3444
rect 70756 3388 72044 3444
rect 72100 3388 72110 3444
rect 72268 3388 85708 3444
rect 86370 3388 86380 3444
rect 86436 3388 86716 3444
rect 86772 3388 86782 3444
rect 88162 3388 88172 3444
rect 88228 3388 88732 3444
rect 88788 3388 88798 3444
rect 90178 3388 90188 3444
rect 90244 3388 90636 3444
rect 90692 3388 90702 3444
rect 91970 3388 91980 3444
rect 92036 3388 92316 3444
rect 92372 3388 92382 3444
rect 92866 3388 92876 3444
rect 92932 3388 93100 3444
rect 93156 3388 93166 3444
rect 93314 3388 93324 3444
rect 93380 3388 93436 3444
rect 93492 3388 93502 3444
rect 95330 3388 95340 3444
rect 95396 3388 95676 3444
rect 95732 3388 95742 3444
rect 96674 3388 96684 3444
rect 96740 3388 97356 3444
rect 97412 3388 97422 3444
rect 98018 3388 98028 3444
rect 98084 3388 98700 3444
rect 98756 3388 98766 3444
rect 100034 3388 100044 3444
rect 100100 3388 100492 3444
rect 100548 3388 100558 3444
rect 102022 3388 102060 3444
rect 102116 3388 102126 3444
rect 102452 3388 108724 3444
rect 114258 3388 114268 3444
rect 114324 3388 114362 3444
rect 193218 3388 193228 3444
rect 193284 3388 194124 3444
rect 194180 3388 194190 3444
rect 268342 3388 268380 3444
rect 268436 3388 268446 3444
rect 308326 3388 308364 3444
rect 308420 3388 308430 3444
rect 409238 3388 409276 3444
rect 409332 3388 409342 3444
rect 414950 3388 414988 3444
rect 415044 3388 415054 3444
rect 462550 3388 462588 3444
rect 462644 3388 462654 3444
rect 563462 3388 563500 3444
rect 563556 3388 563566 3444
rect 55412 3332 55468 3388
rect 42466 3276 42476 3332
rect 42532 3276 43596 3332
rect 43652 3276 43662 3332
rect 45798 3276 45836 3332
rect 45892 3276 45902 3332
rect 50082 3276 50092 3332
rect 50148 3276 52556 3332
rect 52612 3276 52622 3332
rect 54786 3276 54796 3332
rect 54852 3276 55468 3332
rect 56102 3276 56140 3332
rect 56196 3276 56206 3332
rect 57474 3276 57484 3332
rect 57540 3276 57596 3332
rect 57652 3276 57662 3332
rect 58482 3276 58492 3332
rect 58548 3276 59948 3332
rect 60004 3276 60014 3332
rect 60610 3276 60620 3332
rect 60676 3276 61852 3332
rect 61908 3276 61918 3332
rect 63186 3276 63196 3332
rect 63252 3276 63756 3332
rect 63812 3276 63822 3332
rect 63970 3276 63980 3332
rect 64036 3276 79268 3332
rect 79426 3276 79436 3332
rect 79492 3276 81676 3332
rect 81732 3276 81742 3332
rect 84354 3276 84364 3332
rect 84420 3276 86604 3332
rect 86660 3276 86670 3332
rect 91522 3276 91532 3332
rect 91588 3276 92204 3332
rect 92260 3276 92270 3332
rect 92866 3276 92876 3332
rect 92932 3276 93996 3332
rect 94052 3276 94062 3332
rect 94658 3276 94668 3332
rect 94724 3276 95564 3332
rect 95620 3276 95630 3332
rect 95778 3276 95788 3332
rect 95844 3276 97132 3332
rect 97188 3276 97198 3332
rect 97570 3276 97580 3332
rect 97636 3276 98812 3332
rect 98868 3276 98878 3332
rect 101388 3276 123452 3332
rect 123508 3276 123518 3332
rect 40674 3164 40684 3220
rect 40740 3164 60508 3220
rect 60564 3164 60574 3220
rect 62626 3164 62636 3220
rect 62692 3164 63532 3220
rect 63588 3164 63598 3220
rect 67330 3164 67340 3220
rect 67396 3164 68684 3220
rect 68740 3164 68750 3220
rect 69794 3164 69804 3220
rect 69860 3164 72044 3220
rect 72100 3164 72110 3220
rect 73154 3164 73164 3220
rect 73220 3164 74732 3220
rect 74788 3164 74798 3220
rect 75058 3164 75068 3220
rect 75124 3164 75180 3220
rect 75236 3164 75246 3220
rect 76738 3164 76748 3220
rect 76804 3164 78428 3220
rect 78484 3164 78494 3220
rect 79212 3108 79268 3276
rect 92642 3164 92652 3220
rect 92708 3164 93772 3220
rect 93828 3164 93838 3220
rect 94434 3164 94444 3220
rect 94500 3164 95564 3220
rect 95620 3164 95630 3220
rect 98242 3164 98252 3220
rect 98308 3164 98318 3220
rect 98886 3164 98924 3220
rect 98980 3164 98990 3220
rect 98252 3108 98308 3164
rect 101388 3108 101444 3276
rect 15362 3052 15372 3108
rect 15428 3052 35084 3108
rect 35140 3052 35150 3108
rect 42242 3052 42252 3108
rect 42308 3052 43708 3108
rect 43782 3052 43820 3108
rect 43876 3052 43886 3108
rect 56550 3052 56588 3108
rect 56644 3052 56654 3108
rect 62178 3052 62188 3108
rect 62244 3052 63420 3108
rect 63476 3052 63486 3108
rect 66658 3052 66668 3108
rect 66724 3052 68012 3108
rect 68068 3052 68078 3108
rect 68226 3052 68236 3108
rect 68292 3052 68348 3108
rect 68404 3052 68414 3108
rect 74274 3052 74284 3108
rect 74340 3052 76860 3108
rect 76916 3052 76926 3108
rect 78082 3052 78092 3108
rect 78148 3052 78988 3108
rect 79212 3052 95284 3108
rect 98252 3052 101444 3108
rect 102452 3164 123564 3220
rect 123620 3164 123630 3220
rect 43652 2996 43708 3052
rect 78932 2996 78988 3052
rect 95228 2996 95284 3052
rect 102452 2996 102508 3164
rect 43652 2940 76244 2996
rect 78932 2940 85036 2996
rect 85092 2940 85102 2996
rect 95218 2940 95228 2996
rect 95284 2940 95294 2996
rect 95564 2940 102508 2996
rect 114212 3052 485548 3108
rect 485604 3052 485614 3108
rect 41794 2828 41804 2884
rect 41860 2828 72380 2884
rect 72436 2828 72446 2884
rect 74134 2828 74172 2884
rect 74228 2828 74238 2884
rect 76188 2772 76244 2940
rect 79762 2828 79772 2884
rect 79828 2828 79996 2884
rect 80052 2828 80062 2884
rect 83570 2828 83580 2884
rect 83636 2828 83804 2884
rect 83860 2828 83870 2884
rect 87462 2828 87500 2884
rect 87556 2828 87566 2884
rect 90402 2828 90412 2884
rect 90468 2828 95228 2884
rect 95284 2828 95294 2884
rect 95564 2772 95620 2940
rect 114212 2884 114268 3052
rect 95890 2828 95900 2884
rect 95956 2828 114268 2884
rect 41122 2716 41132 2772
rect 41188 2716 66556 2772
rect 66612 2716 66622 2772
rect 68114 2716 68124 2772
rect 68180 2716 68572 2772
rect 68628 2716 68638 2772
rect 71698 2716 71708 2772
rect 71764 2716 74844 2772
rect 74900 2716 74910 2772
rect 76178 2716 76188 2772
rect 76244 2716 76254 2772
rect 79090 2716 79100 2772
rect 79156 2716 80444 2772
rect 80500 2716 80510 2772
rect 91074 2716 91084 2772
rect 91140 2716 95620 2772
rect 95890 2716 95900 2772
rect 95956 2716 97020 2772
rect 97076 2716 97086 2772
rect 98998 2716 99036 2772
rect 99092 2716 99102 2772
rect 40450 2604 40460 2660
rect 40516 2604 60956 2660
rect 61012 2604 61022 2660
rect 62934 2604 62972 2660
rect 63028 2604 63038 2660
rect 63186 2604 63196 2660
rect 63252 2604 64372 2660
rect 64726 2604 64764 2660
rect 64820 2604 64830 2660
rect 77942 2604 77980 2660
rect 78036 2604 78046 2660
rect 85698 2604 85708 2660
rect 85764 2604 91532 2660
rect 91588 2604 91598 2660
rect 93174 2604 93212 2660
rect 93268 2604 93278 2660
rect 95190 2604 95228 2660
rect 95284 2604 95294 2660
rect 95666 2604 95676 2660
rect 95732 2604 124012 2660
rect 124068 2604 124078 2660
rect 64316 2548 64372 2604
rect 41570 2492 41580 2548
rect 41636 2492 64260 2548
rect 64316 2492 67228 2548
rect 75618 2492 75628 2548
rect 75684 2492 78652 2548
rect 78708 2492 78718 2548
rect 78866 2492 78876 2548
rect 78932 2492 96348 2548
rect 96404 2492 96414 2548
rect 121762 2492 121772 2548
rect 121828 2492 445452 2548
rect 445508 2492 445518 2548
rect 42914 2380 42924 2436
rect 42980 2380 63196 2436
rect 63252 2380 63262 2436
rect 64204 2324 64260 2492
rect 67172 2436 67228 2492
rect 67172 2380 81788 2436
rect 81844 2380 81854 2436
rect 46274 2268 46284 2324
rect 46340 2268 47516 2324
rect 47572 2268 47582 2324
rect 53106 2268 53116 2324
rect 53172 2268 53228 2324
rect 53284 2268 53294 2324
rect 57110 2268 57148 2324
rect 57204 2268 57214 2324
rect 58902 2268 58940 2324
rect 58996 2268 59006 2324
rect 60498 2268 60508 2324
rect 60564 2268 62748 2324
rect 62804 2268 62814 2324
rect 63970 2268 63980 2324
rect 64036 2268 64046 2324
rect 64204 2268 67228 2324
rect 68786 2268 68796 2324
rect 68852 2268 102732 2324
rect 102788 2268 102798 2324
rect 63980 2212 64036 2268
rect 49858 2156 49868 2212
rect 49924 2156 64036 2212
rect 67172 2212 67228 2268
rect 67172 2156 70364 2212
rect 70420 2156 70430 2212
rect 72146 2156 72156 2212
rect 72212 2156 91308 2212
rect 91364 2156 91374 2212
rect 56914 2044 56924 2100
rect 56980 2044 100828 2100
rect 100884 2044 100894 2100
rect 117926 2044 117964 2100
rect 118020 2044 118030 2100
rect 524178 2044 524188 2100
rect 524244 2044 542668 2100
rect 542724 2044 542734 2100
rect 67172 1932 186508 1988
rect 186564 1932 186574 1988
rect 197894 1932 197932 1988
rect 197988 1932 197998 1988
rect 498978 1932 498988 1988
rect 499044 1932 536844 1988
rect 536900 1932 536910 1988
rect 67172 1764 67228 1932
rect 85932 1820 90748 1876
rect 93986 1820 93996 1876
rect 94052 1820 382620 1876
rect 382676 1820 382686 1876
rect 456866 1820 456876 1876
rect 456932 1820 525420 1876
rect 525476 1820 525486 1876
rect 542546 1820 542556 1876
rect 542612 1820 559692 1876
rect 559748 1820 559758 1876
rect 85932 1764 85988 1820
rect 90692 1764 90748 1820
rect 44268 1708 44772 1764
rect 44268 1652 44324 1708
rect 44716 1652 44772 1708
rect 47852 1708 48356 1764
rect 47852 1652 47908 1708
rect 48300 1652 48356 1708
rect 61292 1708 67228 1764
rect 80546 1708 80556 1764
rect 80612 1708 85708 1764
rect 85764 1708 85774 1764
rect 85922 1708 85932 1764
rect 85988 1708 85998 1764
rect 89366 1708 89404 1764
rect 89460 1708 89470 1764
rect 90692 1708 405468 1764
rect 405524 1708 405534 1764
rect 426738 1708 426748 1764
rect 426804 1708 519708 1764
rect 519764 1708 519774 1764
rect 519932 1708 548268 1764
rect 548324 1708 548334 1764
rect 557750 1708 557788 1764
rect 557844 1708 557854 1764
rect 569538 1708 569548 1764
rect 569604 1708 571228 1764
rect 571284 1708 571294 1764
rect 38210 1596 38220 1652
rect 38276 1596 40796 1652
rect 40852 1596 40862 1652
rect 44034 1596 44044 1652
rect 44100 1596 44324 1652
rect 44482 1596 44492 1652
rect 44548 1596 44558 1652
rect 44716 1596 47908 1652
rect 48038 1596 48076 1652
rect 48132 1596 48142 1652
rect 48300 1596 53284 1652
rect 53414 1596 53452 1652
rect 53508 1596 53518 1652
rect 58118 1596 58156 1652
rect 58212 1596 58222 1652
rect 44492 1540 44548 1596
rect 53228 1540 53284 1596
rect 61292 1540 61348 1708
rect 61478 1596 61516 1652
rect 61572 1596 61582 1652
rect 61954 1596 61964 1652
rect 62020 1596 66444 1652
rect 66500 1596 66510 1652
rect 69570 1596 69580 1652
rect 69636 1596 69646 1652
rect 70018 1596 70028 1652
rect 70084 1596 74956 1652
rect 75012 1596 75022 1652
rect 76262 1596 76300 1652
rect 76356 1596 76366 1652
rect 79650 1596 79660 1652
rect 79716 1596 83244 1652
rect 83300 1596 83310 1652
rect 85474 1596 85484 1652
rect 85540 1596 88172 1652
rect 88228 1596 88238 1652
rect 88844 1596 90748 1652
rect 90804 1596 90814 1652
rect 91746 1596 91756 1652
rect 91812 1596 95340 1652
rect 95396 1596 95406 1652
rect 98438 1596 98476 1652
rect 98532 1596 98542 1652
rect 99110 1596 99148 1652
rect 99204 1596 99214 1652
rect 100454 1596 100492 1652
rect 100548 1596 100558 1652
rect 69580 1540 69636 1596
rect 88844 1540 88900 1596
rect 519932 1540 519988 1708
rect 34402 1484 34412 1540
rect 34468 1484 36988 1540
rect 37044 1484 37054 1540
rect 38098 1484 38108 1540
rect 38164 1484 39900 1540
rect 39956 1484 39966 1540
rect 40226 1484 40236 1540
rect 40292 1484 44436 1540
rect 44492 1484 49868 1540
rect 49924 1484 49934 1540
rect 53228 1484 54292 1540
rect 55234 1484 55244 1540
rect 55300 1484 61348 1540
rect 62374 1484 62412 1540
rect 62468 1484 62478 1540
rect 65734 1484 65772 1540
rect 65828 1484 65838 1540
rect 69580 1484 78876 1540
rect 78932 1484 78942 1540
rect 80994 1484 81004 1540
rect 81060 1484 85932 1540
rect 85988 1484 85998 1540
rect 87042 1484 87052 1540
rect 87108 1484 88900 1540
rect 89730 1484 89740 1540
rect 89796 1484 95004 1540
rect 95060 1484 95070 1540
rect 97794 1484 97804 1540
rect 97860 1484 519988 1540
rect 44380 1428 44436 1484
rect 54236 1428 54292 1484
rect 31938 1372 31948 1428
rect 32004 1372 36652 1428
rect 36708 1372 36718 1428
rect 38434 1372 38444 1428
rect 38500 1372 43708 1428
rect 43764 1372 43774 1428
rect 44380 1372 46620 1428
rect 46676 1372 46686 1428
rect 47170 1372 47180 1428
rect 47236 1372 48636 1428
rect 48692 1372 48702 1428
rect 50754 1372 50764 1428
rect 50820 1372 54012 1428
rect 54068 1372 54078 1428
rect 54236 1372 72156 1428
rect 72212 1372 72222 1428
rect 72380 1372 77308 1428
rect 77364 1372 77374 1428
rect 78306 1372 78316 1428
rect 78372 1372 93996 1428
rect 94052 1372 94062 1428
rect 95106 1372 95116 1428
rect 95172 1372 96292 1428
rect 96450 1372 96460 1428
rect 96516 1372 498988 1428
rect 499044 1372 499054 1428
rect 72380 1316 72436 1372
rect 96236 1316 96292 1372
rect 39106 1260 39116 1316
rect 39172 1260 49420 1316
rect 49476 1260 49486 1316
rect 52546 1260 52556 1316
rect 52612 1260 72436 1316
rect 74050 1260 74060 1316
rect 74116 1260 79660 1316
rect 79716 1260 79726 1316
rect 80322 1260 80332 1316
rect 80388 1260 80398 1316
rect 81666 1260 81676 1316
rect 81732 1260 81788 1316
rect 81844 1260 81854 1316
rect 82338 1260 82348 1316
rect 82404 1260 87276 1316
rect 87332 1260 87342 1316
rect 87500 1260 95676 1316
rect 95732 1260 95742 1316
rect 96236 1260 456876 1316
rect 456932 1260 456942 1316
rect 80332 1204 80388 1260
rect 87500 1204 87556 1260
rect 35410 1148 35420 1204
rect 35476 1148 36204 1204
rect 36260 1148 36270 1204
rect 45378 1148 45388 1204
rect 45444 1148 68796 1204
rect 68852 1148 68862 1204
rect 70914 1148 70924 1204
rect 70980 1148 80108 1204
rect 80164 1148 80174 1204
rect 80332 1148 87556 1204
rect 87714 1148 87724 1204
rect 87780 1148 93884 1204
rect 93940 1148 93950 1204
rect 94434 1148 94444 1204
rect 94500 1148 426748 1204
rect 426804 1148 426814 1204
rect 13346 1036 13356 1092
rect 13412 1036 34860 1092
rect 34916 1036 34926 1092
rect 43362 1036 43372 1092
rect 43428 1036 80556 1092
rect 80612 1036 80622 1092
rect 85026 1036 85036 1092
rect 85092 1036 90972 1092
rect 91028 1036 91038 1092
rect 93762 1036 93772 1092
rect 93828 1036 299068 1092
rect 299124 1036 299134 1092
rect 26786 924 26796 980
rect 26852 924 36428 980
rect 36484 924 36494 980
rect 38658 924 38668 980
rect 38724 924 45612 980
rect 45668 924 45678 980
rect 49298 924 49308 980
rect 49364 924 55300 980
rect 55458 924 55468 980
rect 55524 924 188412 980
rect 188468 924 188478 980
rect 55244 868 55300 924
rect 30594 812 30604 868
rect 30660 812 32228 868
rect 36866 812 36876 868
rect 36932 812 36942 868
rect 39778 812 39788 868
rect 39844 812 55020 868
rect 55076 812 55086 868
rect 55244 812 62188 868
rect 62244 812 62254 868
rect 80098 812 80108 868
rect 80164 812 83020 868
rect 83076 812 83086 868
rect 92418 812 92428 868
rect 92484 812 127036 868
rect 127092 812 127102 868
rect 32172 756 32228 812
rect 36876 756 36932 812
rect 28690 700 28700 756
rect 28756 700 31892 756
rect 31948 700 31958 756
rect 32172 700 36932 756
rect 52098 700 52108 756
rect 52164 700 84700 756
rect 84756 700 84766 756
rect 97346 700 97356 756
rect 97412 700 524188 756
rect 524244 700 524254 756
rect 24882 588 24892 644
rect 24948 588 35420 644
rect 35476 588 35486 644
rect 56802 588 56812 644
rect 56868 588 61908 644
rect 211222 588 211260 644
rect 211316 588 211326 644
rect 23090 476 23100 532
rect 23156 476 35980 532
rect 36036 476 36046 532
rect 42466 476 42476 532
rect 42532 476 43708 532
rect 45154 476 45164 532
rect 45220 476 56924 532
rect 56980 476 56990 532
rect 43652 420 43708 476
rect 21746 364 21756 420
rect 21812 364 35756 420
rect 35812 364 35822 420
rect 43652 364 53788 420
rect 53844 364 53854 420
rect 19282 252 19292 308
rect 19348 252 35420 308
rect 35476 252 35486 308
rect 17378 140 17388 196
rect 17444 140 35308 196
rect 35364 140 35374 196
rect 61852 84 61908 588
rect 66882 476 66892 532
rect 66948 476 78540 532
rect 78596 476 78606 532
rect 88386 476 88396 532
rect 88452 476 94892 532
rect 94948 476 94958 532
rect 78754 252 78764 308
rect 78820 252 84924 308
rect 84980 252 84990 308
rect 39218 28 39228 84
rect 39284 28 51212 84
rect 51268 28 51278 84
rect 61852 28 199724 84
rect 199780 28 199790 84
<< via3 >>
rect 27692 590604 27748 590660
rect 99260 590156 99316 590212
rect 120988 590156 121044 590212
rect 164668 590156 164724 590212
rect 186508 590156 186564 590212
rect 297388 590156 297444 590212
rect 341068 590156 341124 590212
rect 26012 588588 26068 588644
rect 3388 587132 3444 587188
rect 22652 582092 22708 582148
rect 19292 578732 19348 578788
rect 17612 575372 17668 575428
rect 12012 573020 12068 573076
rect 590716 562156 590772 562212
rect 10892 558908 10948 558964
rect 24332 548940 24388 548996
rect 28 544684 84 544740
rect 15148 530684 15204 530740
rect 3164 523292 3220 523348
rect 590716 523292 590772 523348
rect 590492 522508 590548 522564
rect 11900 516572 11956 516628
rect 14252 509292 14308 509348
rect 2492 502460 2548 502516
rect 590156 496076 590212 496132
rect 31052 494732 31108 494788
rect 590156 494732 590212 494788
rect 13468 488348 13524 488404
rect 8316 482860 8372 482916
rect 140 474124 196 474180
rect 7532 460124 7588 460180
rect 20972 456428 21028 456484
rect 4620 446012 4676 446068
rect 86492 443212 86548 443268
rect 4172 431900 4228 431956
rect 11676 430108 11732 430164
rect 252 417676 308 417732
rect 76412 416780 76468 416836
rect 13580 403676 13636 403732
rect 8204 403564 8260 403620
rect 29372 390348 29428 390404
rect 4284 389564 4340 389620
rect 2604 375452 2660 375508
rect 587132 363916 587188 363972
rect 4732 361340 4788 361396
rect 15932 350700 15988 350756
rect 2716 347228 2772 347284
rect 21084 337484 21140 337540
rect 588 333116 644 333172
rect 47852 324268 47908 324324
rect 11788 319004 11844 319060
rect 126812 311052 126868 311108
rect 4396 304892 4452 304948
rect 4620 304108 4676 304164
rect 11004 304108 11060 304164
rect 590156 297836 590212 297892
rect 150332 296492 150388 296548
rect 590156 296492 590212 296548
rect 7644 290780 7700 290836
rect 173852 284620 173908 284676
rect 4508 276668 4564 276724
rect 4732 275548 4788 275604
rect 6188 275548 6244 275604
rect 145292 271404 145348 271460
rect 4620 262556 4676 262612
rect 126924 258188 126980 258244
rect 591276 244972 591332 245028
rect 136892 242732 136948 242788
rect 591276 242732 591332 242788
rect 148652 231868 148708 231924
rect 127036 218540 127092 218596
rect 135212 205324 135268 205380
rect 141932 192108 141988 192164
rect 127148 178892 127204 178948
rect 590156 165676 590212 165732
rect 133532 163772 133588 163828
rect 590156 163772 590212 163828
rect 140252 152460 140308 152516
rect 127260 139244 127316 139300
rect 129052 126028 129108 126084
rect 138572 112812 138628 112868
rect 8652 104972 8708 105028
rect 587132 104972 587188 105028
rect 590156 99596 590212 99652
rect 474572 98252 474628 98308
rect 590156 98252 590212 98308
rect 504812 86380 504868 86436
rect 46956 82684 47012 82740
rect 114268 82684 114324 82740
rect 47628 82572 47684 82628
rect 121100 82572 121156 82628
rect 48524 82460 48580 82516
rect 43596 82348 43652 82404
rect 9884 81452 9940 81508
rect 47852 81452 47908 81508
rect 46844 81004 46900 81060
rect 110908 81004 110964 81060
rect 48300 80892 48356 80948
rect 119308 80892 119364 80948
rect 48412 80780 48468 80836
rect 70364 80668 70420 80724
rect 84812 79884 84868 79940
rect 65436 79772 65492 79828
rect 76524 79660 76580 79716
rect 75852 79548 75908 79604
rect 81564 79436 81620 79492
rect 78316 79324 78372 79380
rect 78876 79212 78932 79268
rect 81788 79100 81844 79156
rect 86604 78316 86660 78372
rect 70252 78204 70308 78260
rect 71708 78092 71764 78148
rect 76636 77980 76692 78036
rect 73052 77868 73108 77924
rect 74508 77756 74564 77812
rect 79436 77644 79492 77700
rect 83020 77532 83076 77588
rect 85596 77420 85652 77476
rect 100156 77308 100212 77364
rect 87948 76524 88004 76580
rect 60284 76412 60340 76468
rect 60396 76300 60452 76356
rect 52780 76188 52836 76244
rect 72492 76076 72548 76132
rect 73836 75964 73892 76020
rect 75404 75852 75460 75908
rect 81452 75740 81508 75796
rect 94444 75628 94500 75684
rect 82572 74844 82628 74900
rect 9996 74732 10052 74788
rect 21084 74732 21140 74788
rect 62076 74732 62132 74788
rect 65324 74620 65380 74676
rect 61964 74508 62020 74564
rect 67788 74396 67844 74452
rect 69132 74284 69188 74340
rect 72716 74172 72772 74228
rect 77084 74060 77140 74116
rect 8764 73948 8820 74004
rect 11788 73948 11844 74004
rect 91532 73948 91588 74004
rect 121772 73948 121828 74004
rect 74732 73500 74788 73556
rect 57484 73388 57540 73444
rect 58492 73276 58548 73332
rect 130172 73164 130228 73220
rect 58044 73052 58100 73108
rect 8540 72940 8596 72996
rect 13580 72940 13636 72996
rect 66668 72940 66724 72996
rect 56364 72828 56420 72884
rect 68796 72716 68852 72772
rect 126812 72492 126868 72548
rect 9884 70700 9940 70756
rect 9996 69804 10052 69860
rect 9996 69580 10052 69636
rect 150332 69580 150388 69636
rect 12684 68908 12740 68964
rect 8652 68012 8708 68068
rect 9996 67116 10052 67172
rect 12572 66892 12628 66948
rect 173852 66668 173908 66724
rect 9996 65548 10052 65604
rect 8204 65324 8260 65380
rect 12460 64988 12516 65044
rect 145292 63756 145348 63812
rect 11340 63532 11396 63588
rect 12460 63308 12516 63364
rect 12684 61740 12740 61796
rect 9996 60844 10052 60900
rect 126924 60844 126980 60900
rect 8316 59948 8372 60004
rect 126812 59948 126868 60004
rect 12460 59612 12516 59668
rect 12572 58716 12628 58772
rect 136892 57932 136948 57988
rect 11452 57260 11508 57316
rect 12348 56140 12404 56196
rect 148652 55020 148708 55076
rect 3164 54572 3220 54628
rect 12684 53676 12740 53732
rect 12348 53452 12404 53508
rect 127036 52108 127092 52164
rect 12348 51660 12404 51716
rect 135212 49196 135268 49252
rect 12684 48300 12740 48356
rect 127596 47852 127652 47908
rect 141932 47852 141988 47908
rect 590492 46732 590548 46788
rect 127596 46284 127652 46340
rect 9996 44716 10052 44772
rect 127148 43372 127204 43428
rect 6524 42028 6580 42084
rect 133532 40460 133588 40516
rect 6636 40236 6692 40292
rect 140252 37548 140308 37604
rect 11564 35756 11620 35812
rect 7980 34860 8036 34916
rect 127260 34636 127316 34692
rect 127036 33628 127092 33684
rect 4620 33516 4676 33572
rect 7756 33516 7812 33572
rect 8092 33068 8148 33124
rect 127372 32732 127428 32788
rect 504812 32732 504868 32788
rect 3052 32172 3108 32228
rect 127148 31948 127204 32004
rect 587132 31948 587188 32004
rect 129052 31724 129108 31780
rect 127260 31052 127316 31108
rect 590492 31052 590548 31108
rect 126924 30380 126980 30436
rect 127484 30268 127540 30324
rect 130172 30268 130228 30324
rect 575372 30268 575428 30324
rect 138572 28812 138628 28868
rect 3276 27692 3332 27748
rect 12012 26796 12068 26852
rect 10892 25900 10948 25956
rect 474572 25900 474628 25956
rect 28 25004 84 25060
rect 8988 24108 9044 24164
rect 130172 23548 130228 23604
rect 12012 23212 12068 23268
rect 127372 22988 127428 23044
rect 2492 22316 2548 22372
rect 8876 21420 8932 21476
rect 140 20524 196 20580
rect 587132 20524 587188 20580
rect 127484 20076 127540 20132
rect 7532 19628 7588 19684
rect 11004 18732 11060 18788
rect 4172 17836 4228 17892
rect 126812 17164 126868 17220
rect 252 16940 308 16996
rect 8540 16044 8596 16100
rect 4284 15148 4340 15204
rect 2604 14252 2660 14308
rect 127260 14252 127316 14308
rect 6188 13356 6244 13412
rect 2716 12460 2772 12516
rect 364 11564 420 11620
rect 127036 11340 127092 11396
rect 124012 10892 124068 10948
rect 8764 10668 8820 10724
rect 4396 9772 4452 9828
rect 7644 8876 7700 8932
rect 127148 8428 127204 8484
rect 4508 7980 4564 8036
rect 7756 7084 7812 7140
rect 575372 7084 575428 7140
rect 123452 6748 123508 6804
rect 126924 5516 126980 5572
rect 75068 4508 75124 4564
rect 76524 4508 76580 4564
rect 79548 4508 79604 4564
rect 80668 4508 80724 4564
rect 85708 4508 85764 4564
rect 93324 4508 93380 4564
rect 57596 4396 57652 4452
rect 62860 4284 62916 4340
rect 84700 4284 84756 4340
rect 91420 4284 91476 4340
rect 92764 4284 92820 4340
rect 93436 4284 93492 4340
rect 57148 4172 57204 4228
rect 61628 4172 61684 4228
rect 62188 4172 62244 4228
rect 79772 4172 79828 4228
rect 82124 4172 82180 4228
rect 120988 4172 121044 4228
rect 126028 4172 126084 4228
rect 131292 4172 131348 4228
rect 132748 4172 132804 4228
rect 134428 4172 134484 4228
rect 137788 4172 137844 4228
rect 139468 4172 139524 4228
rect 142828 4172 142884 4228
rect 144620 4172 144676 4228
rect 146188 4172 146244 4228
rect 147868 4172 147924 4228
rect 149548 4172 149604 4228
rect 151228 4172 151284 4228
rect 152908 4172 152964 4228
rect 154588 4172 154644 4228
rect 157948 4172 158004 4228
rect 161308 4172 161364 4228
rect 163660 4172 163716 4228
rect 164668 4172 164724 4228
rect 166348 4172 166404 4228
rect 169372 4172 169428 4228
rect 173180 4172 173236 4228
rect 174748 4172 174804 4228
rect 178108 4172 178164 4228
rect 179788 4172 179844 4228
rect 183148 4172 183204 4228
rect 190428 4172 190484 4228
rect 191548 4172 191604 4228
rect 194908 4172 194964 4228
rect 201740 4172 201796 4228
rect 203644 4172 203700 4228
rect 206668 4172 206724 4228
rect 215068 4172 215124 4228
rect 216972 4172 217028 4228
rect 220108 4172 220164 4228
rect 221788 4172 221844 4228
rect 223468 4172 223524 4228
rect 228508 4172 228564 4228
rect 231868 4172 231924 4228
rect 233548 4172 233604 4228
rect 235228 4172 235284 4228
rect 236908 4172 236964 4228
rect 238588 4172 238644 4228
rect 243628 4172 243684 4228
rect 245532 4172 245588 4228
rect 248668 4172 248724 4228
rect 250348 4172 250404 4228
rect 252028 4172 252084 4228
rect 253708 4172 253764 4228
rect 258860 4172 258916 4228
rect 260428 4172 260484 4228
rect 262108 4172 262164 4228
rect 263788 4172 263844 4228
rect 265468 4172 265524 4228
rect 274092 4172 274148 4228
rect 278908 4172 278964 4228
rect 282604 4172 282660 4228
rect 286300 4172 286356 4228
rect 288988 4172 289044 4228
rect 290668 4172 290724 4228
rect 294028 4172 294084 4228
rect 295708 4172 295764 4228
rect 300748 4172 300804 4228
rect 302652 4172 302708 4228
rect 305788 4172 305844 4228
rect 310828 4172 310884 4228
rect 314188 4172 314244 4228
rect 317548 4172 317604 4228
rect 319228 4172 319284 4228
rect 322588 4172 322644 4228
rect 324268 4172 324324 4228
rect 331212 4172 331268 4228
rect 336028 4172 336084 4228
rect 339388 4172 339444 4228
rect 342748 4172 342804 4228
rect 346108 4172 346164 4228
rect 347788 4172 347844 4228
rect 351148 4172 351204 4228
rect 352828 4172 352884 4228
rect 359772 4172 359828 4228
rect 362908 4172 362964 4228
rect 364588 4172 364644 4228
rect 371308 4172 371364 4228
rect 375004 4172 375060 4228
rect 376348 4172 376404 4228
rect 379708 4172 379764 4228
rect 383068 4172 383124 4228
rect 386428 4172 386484 4228
rect 388332 4172 388388 4228
rect 391468 4172 391524 4228
rect 393148 4172 393204 4228
rect 394828 4172 394884 4228
rect 396508 4172 396564 4228
rect 403228 4172 403284 4228
rect 406588 4172 406644 4228
rect 409948 4172 410004 4228
rect 416892 4172 416948 4228
rect 420028 4172 420084 4228
rect 422604 4172 422660 4228
rect 425068 4172 425124 4228
rect 428428 4172 428484 4228
rect 431788 4172 431844 4228
rect 435148 4172 435204 4228
rect 436828 4172 436884 4228
rect 438508 4172 438564 4228
rect 443548 4172 443604 4228
rect 446908 4172 446964 4228
rect 448588 4172 448644 4228
rect 450268 4172 450324 4228
rect 451948 4172 452004 4228
rect 453628 4172 453684 4228
rect 456988 4172 457044 4228
rect 458780 4172 458836 4228
rect 460348 4172 460404 4228
rect 465388 4172 465444 4228
rect 468748 4172 468804 4228
rect 472108 4172 472164 4228
rect 474012 4172 474068 4228
rect 475468 4172 475524 4228
rect 477148 4172 477204 4228
rect 478828 4172 478884 4228
rect 480508 4172 480564 4228
rect 482188 4172 482244 4228
rect 487340 4172 487396 4228
rect 488908 4172 488964 4228
rect 492268 4172 492324 4228
rect 493948 4172 494004 4228
rect 495628 4172 495684 4228
rect 497644 4172 497700 4228
rect 501340 4172 501396 4228
rect 504028 4172 504084 4228
rect 505708 4172 505764 4228
rect 508284 4172 508340 4228
rect 509068 4172 509124 4228
rect 510748 4172 510804 4228
rect 515900 4172 515956 4228
rect 517468 4172 517524 4228
rect 520828 4172 520884 4228
rect 522508 4172 522564 4228
rect 525868 4172 525924 4228
rect 531132 4172 531188 4228
rect 532588 4172 532644 4228
rect 534268 4172 534324 4228
rect 537628 4172 537684 4228
rect 539308 4172 539364 4228
rect 544460 4172 544516 4228
rect 549388 4172 549444 4228
rect 554428 4172 554484 4228
rect 561148 4172 561204 4228
rect 564508 4172 564564 4228
rect 566188 4172 566244 4228
rect 573020 4172 573076 4228
rect 574588 4172 574644 4228
rect 576268 4172 576324 4228
rect 53116 4060 53172 4116
rect 54124 4060 54180 4116
rect 68124 4060 68180 4116
rect 68908 4060 68964 4116
rect 70140 4060 70196 4116
rect 72268 4060 72324 4116
rect 73724 4060 73780 4116
rect 40908 3724 40964 3780
rect 74172 3948 74228 4004
rect 79548 3948 79604 4004
rect 91420 3948 91476 4004
rect 61628 3836 61684 3892
rect 79996 3836 80052 3892
rect 80668 3836 80724 3892
rect 43148 3724 43204 3780
rect 44268 3724 44324 3780
rect 44716 3724 44772 3780
rect 44940 3724 44996 3780
rect 45612 3724 45668 3780
rect 46508 3724 46564 3780
rect 46844 3724 46900 3780
rect 47628 3724 47684 3780
rect 48188 3724 48244 3780
rect 48524 3724 48580 3780
rect 48972 3724 49028 3780
rect 49196 3724 49252 3780
rect 49868 3724 49924 3780
rect 50316 3724 50372 3780
rect 50540 3724 50596 3780
rect 50988 3724 51044 3780
rect 51212 3724 51268 3780
rect 51772 3724 51828 3780
rect 52332 3724 52388 3780
rect 53228 3724 53284 3780
rect 53452 3724 53508 3780
rect 53900 3724 53956 3780
rect 54124 3724 54180 3780
rect 54348 3724 54404 3780
rect 55244 3724 55300 3780
rect 55692 3724 55748 3780
rect 56700 3724 56756 3780
rect 56924 3724 56980 3780
rect 57260 3724 57316 3780
rect 57708 3724 57764 3780
rect 57932 3724 57988 3780
rect 58380 3724 58436 3780
rect 59052 3724 59108 3780
rect 59276 3724 59332 3780
rect 59500 3724 59556 3780
rect 59724 3724 59780 3780
rect 60172 3724 60228 3780
rect 60396 3724 60452 3780
rect 60844 3724 60900 3780
rect 61068 3724 61124 3780
rect 61292 3724 61348 3780
rect 61740 3724 61796 3780
rect 62860 3724 62916 3780
rect 63644 3724 63700 3780
rect 63980 3724 64036 3780
rect 64204 3724 64260 3780
rect 64428 3724 64484 3780
rect 65100 3724 65156 3780
rect 65436 3724 65492 3780
rect 65996 3724 66052 3780
rect 66332 3724 66388 3780
rect 66668 3724 66724 3780
rect 67788 3724 67844 3780
rect 68460 3724 68516 3780
rect 68908 3724 68964 3780
rect 69132 3724 69188 3780
rect 69468 3724 69524 3780
rect 70140 3724 70196 3780
rect 70364 3724 70420 3780
rect 71596 3724 71652 3780
rect 71932 3724 71988 3780
rect 72268 3724 72324 3780
rect 72492 3724 72548 3780
rect 72716 3724 72772 3780
rect 73164 3724 73220 3780
rect 73500 3724 73556 3780
rect 73836 3724 73892 3780
rect 74508 3724 74564 3780
rect 75180 3724 75236 3780
rect 75404 3724 75460 3780
rect 75852 3724 75908 3780
rect 76076 3724 76132 3780
rect 76972 3724 77028 3780
rect 77644 3724 77700 3780
rect 78876 3724 78932 3780
rect 79436 3724 79492 3780
rect 80556 3724 80612 3780
rect 80780 3724 80836 3780
rect 81228 3724 81284 3780
rect 82012 3724 82068 3780
rect 82572 3724 82628 3780
rect 82796 3724 82852 3780
rect 83020 3724 83076 3780
rect 83692 3724 83748 3780
rect 84140 3724 84196 3780
rect 84588 3724 84644 3780
rect 85484 3724 85540 3780
rect 87276 3836 87332 3892
rect 88956 3836 89012 3892
rect 92988 3836 93044 3892
rect 93324 3836 93380 3892
rect 85932 3724 85988 3780
rect 86156 3724 86212 3780
rect 86828 3724 86884 3780
rect 87164 3724 87220 3780
rect 87724 3724 87780 3780
rect 87948 3724 88004 3780
rect 88844 3724 88900 3780
rect 89068 3724 89124 3780
rect 89292 3724 89348 3780
rect 89516 3724 89572 3780
rect 89740 3724 89796 3780
rect 90412 3724 90468 3780
rect 90860 3724 90916 3780
rect 91308 3724 91364 3780
rect 92092 3724 92148 3780
rect 93660 3724 93716 3780
rect 94220 3724 94276 3780
rect 95452 3724 95508 3780
rect 96012 3724 96068 3780
rect 96236 3724 96292 3780
rect 96460 3724 96516 3780
rect 97244 3724 97300 3780
rect 98588 3724 98644 3780
rect 99372 3724 99428 3780
rect 99596 3724 99652 3780
rect 99820 3724 99876 3780
rect 100156 3724 100212 3780
rect 100604 3724 100660 3780
rect 102396 3724 102452 3780
rect 63308 3612 63364 3668
rect 63756 3612 63812 3668
rect 64876 3612 64932 3668
rect 65324 3612 65380 3668
rect 66220 3612 66276 3668
rect 66444 3612 66500 3668
rect 68796 3612 68852 3668
rect 69916 3612 69972 3668
rect 71708 3612 71764 3668
rect 73612 3612 73668 3668
rect 75292 3612 75348 3668
rect 76748 3612 76804 3668
rect 80108 3612 80164 3668
rect 81900 3612 81956 3668
rect 82124 3612 82180 3668
rect 82908 3612 82964 3668
rect 83804 3612 83860 3668
rect 85372 3612 85428 3668
rect 209356 3612 209412 3668
rect 46396 3500 46452 3556
rect 46732 3500 46788 3556
rect 48412 3500 48468 3556
rect 50204 3500 50260 3556
rect 51996 3500 52052 3556
rect 53564 3500 53620 3556
rect 55356 3500 55412 3556
rect 55580 3500 55636 3556
rect 57484 3500 57540 3556
rect 60284 3500 60340 3556
rect 62076 3500 62132 3556
rect 68572 3500 68628 3556
rect 77084 3500 77140 3556
rect 79884 3500 79940 3556
rect 81452 3500 81508 3556
rect 84812 3500 84868 3556
rect 104188 3500 104244 3556
rect 106540 3500 106596 3556
rect 107548 3500 107604 3556
rect 109228 3500 109284 3556
rect 110908 3500 110964 3556
rect 116060 3500 116116 3556
rect 119308 3500 119364 3556
rect 121100 3500 121156 3556
rect 257068 3500 257124 3556
rect 468300 3500 468356 3556
rect 46284 3388 46340 3444
rect 46956 3388 47012 3444
rect 48300 3388 48356 3444
rect 50092 3388 50148 3444
rect 51884 3388 51940 3444
rect 54572 3388 54628 3444
rect 72044 3388 72100 3444
rect 86716 3388 86772 3444
rect 88732 3388 88788 3444
rect 90636 3388 90692 3444
rect 92316 3388 92372 3444
rect 93100 3388 93156 3444
rect 93436 3388 93492 3444
rect 95676 3388 95732 3444
rect 97356 3388 97412 3444
rect 98700 3388 98756 3444
rect 100492 3388 100548 3444
rect 102060 3388 102116 3444
rect 114268 3388 114324 3444
rect 193228 3388 193284 3444
rect 268380 3388 268436 3444
rect 308364 3388 308420 3444
rect 409276 3388 409332 3444
rect 414988 3388 415044 3444
rect 462588 3388 462644 3444
rect 563500 3388 563556 3444
rect 42476 3276 42532 3332
rect 45836 3276 45892 3332
rect 52556 3276 52612 3332
rect 56140 3276 56196 3332
rect 57596 3276 57652 3332
rect 58492 3276 58548 3332
rect 61852 3276 61908 3332
rect 63196 3276 63252 3332
rect 63980 3276 64036 3332
rect 81676 3276 81732 3332
rect 86604 3276 86660 3332
rect 92204 3276 92260 3332
rect 92876 3276 92932 3332
rect 95564 3276 95620 3332
rect 97132 3276 97188 3332
rect 98812 3276 98868 3332
rect 123452 3276 123508 3332
rect 60508 3164 60564 3220
rect 63532 3164 63588 3220
rect 68684 3164 68740 3220
rect 69804 3164 69860 3220
rect 74732 3164 74788 3220
rect 75068 3164 75124 3220
rect 78428 3164 78484 3220
rect 93772 3164 93828 3220
rect 94444 3164 94500 3220
rect 98924 3164 98980 3220
rect 43820 3052 43876 3108
rect 56588 3052 56644 3108
rect 63420 3052 63476 3108
rect 66668 3052 66724 3108
rect 68348 3052 68404 3108
rect 76860 3052 76916 3108
rect 85036 2940 85092 2996
rect 95228 2940 95284 2996
rect 74172 2828 74228 2884
rect 79772 2828 79828 2884
rect 83580 2828 83636 2884
rect 87500 2828 87556 2884
rect 68124 2716 68180 2772
rect 74844 2716 74900 2772
rect 80444 2716 80500 2772
rect 95900 2716 95956 2772
rect 99036 2716 99092 2772
rect 62972 2604 63028 2660
rect 63196 2604 63252 2660
rect 64764 2604 64820 2660
rect 77980 2604 78036 2660
rect 91532 2604 91588 2660
rect 93212 2604 93268 2660
rect 95228 2604 95284 2660
rect 78652 2492 78708 2548
rect 96348 2492 96404 2548
rect 121772 2492 121828 2548
rect 63196 2380 63252 2436
rect 46284 2268 46340 2324
rect 53116 2268 53172 2324
rect 57148 2268 57204 2324
rect 58940 2268 58996 2324
rect 60508 2268 60564 2324
rect 63980 2268 64036 2324
rect 49868 2156 49924 2212
rect 117964 2044 118020 2100
rect 197932 1932 197988 1988
rect 93996 1820 94052 1876
rect 542556 1820 542612 1876
rect 80556 1708 80612 1764
rect 85932 1708 85988 1764
rect 89404 1708 89460 1764
rect 557788 1708 557844 1764
rect 569548 1708 569604 1764
rect 48076 1596 48132 1652
rect 53452 1596 53508 1652
rect 58156 1596 58212 1652
rect 61516 1596 61572 1652
rect 61964 1596 62020 1652
rect 74956 1596 75012 1652
rect 76300 1596 76356 1652
rect 83244 1596 83300 1652
rect 88172 1596 88228 1652
rect 90748 1596 90804 1652
rect 95340 1596 95396 1652
rect 98476 1596 98532 1652
rect 99148 1596 99204 1652
rect 100492 1596 100548 1652
rect 49868 1484 49924 1540
rect 62412 1484 62468 1540
rect 65772 1484 65828 1540
rect 85932 1484 85988 1540
rect 95004 1484 95060 1540
rect 31948 1372 32004 1428
rect 46620 1372 46676 1428
rect 48636 1372 48692 1428
rect 54012 1372 54068 1428
rect 77308 1372 77364 1428
rect 93996 1372 94052 1428
rect 79660 1260 79716 1316
rect 81788 1260 81844 1316
rect 87276 1260 87332 1316
rect 80108 1148 80164 1204
rect 93884 1148 93940 1204
rect 80556 1036 80612 1092
rect 90972 1036 91028 1092
rect 62188 812 62244 868
rect 80108 812 80164 868
rect 83020 812 83076 868
rect 31892 700 31948 756
rect 84700 700 84756 756
rect 211260 588 211316 644
rect 53788 364 53844 420
rect 78540 476 78596 532
rect 94892 476 94948 532
rect 84924 252 84980 308
<< metal4 >>
rect -1916 598172 -1296 598268
rect -1916 598116 -1820 598172
rect -1764 598116 -1696 598172
rect -1640 598116 -1572 598172
rect -1516 598116 -1448 598172
rect -1392 598116 -1296 598172
rect -1916 598048 -1296 598116
rect -1916 597992 -1820 598048
rect -1764 597992 -1696 598048
rect -1640 597992 -1572 598048
rect -1516 597992 -1448 598048
rect -1392 597992 -1296 598048
rect -1916 597924 -1296 597992
rect -1916 597868 -1820 597924
rect -1764 597868 -1696 597924
rect -1640 597868 -1572 597924
rect -1516 597868 -1448 597924
rect -1392 597868 -1296 597924
rect -1916 597800 -1296 597868
rect -1916 597744 -1820 597800
rect -1764 597744 -1696 597800
rect -1640 597744 -1572 597800
rect -1516 597744 -1448 597800
rect -1392 597744 -1296 597800
rect -1916 586350 -1296 597744
rect -1916 586294 -1820 586350
rect -1764 586294 -1696 586350
rect -1640 586294 -1572 586350
rect -1516 586294 -1448 586350
rect -1392 586294 -1296 586350
rect -1916 586226 -1296 586294
rect -1916 586170 -1820 586226
rect -1764 586170 -1696 586226
rect -1640 586170 -1572 586226
rect -1516 586170 -1448 586226
rect -1392 586170 -1296 586226
rect -1916 586102 -1296 586170
rect -1916 586046 -1820 586102
rect -1764 586046 -1696 586102
rect -1640 586046 -1572 586102
rect -1516 586046 -1448 586102
rect -1392 586046 -1296 586102
rect -1916 585978 -1296 586046
rect -1916 585922 -1820 585978
rect -1764 585922 -1696 585978
rect -1640 585922 -1572 585978
rect -1516 585922 -1448 585978
rect -1392 585922 -1296 585978
rect -1916 568350 -1296 585922
rect -1916 568294 -1820 568350
rect -1764 568294 -1696 568350
rect -1640 568294 -1572 568350
rect -1516 568294 -1448 568350
rect -1392 568294 -1296 568350
rect -1916 568226 -1296 568294
rect -1916 568170 -1820 568226
rect -1764 568170 -1696 568226
rect -1640 568170 -1572 568226
rect -1516 568170 -1448 568226
rect -1392 568170 -1296 568226
rect -1916 568102 -1296 568170
rect -1916 568046 -1820 568102
rect -1764 568046 -1696 568102
rect -1640 568046 -1572 568102
rect -1516 568046 -1448 568102
rect -1392 568046 -1296 568102
rect -1916 567978 -1296 568046
rect -1916 567922 -1820 567978
rect -1764 567922 -1696 567978
rect -1640 567922 -1572 567978
rect -1516 567922 -1448 567978
rect -1392 567922 -1296 567978
rect -1916 550350 -1296 567922
rect -1916 550294 -1820 550350
rect -1764 550294 -1696 550350
rect -1640 550294 -1572 550350
rect -1516 550294 -1448 550350
rect -1392 550294 -1296 550350
rect -1916 550226 -1296 550294
rect -1916 550170 -1820 550226
rect -1764 550170 -1696 550226
rect -1640 550170 -1572 550226
rect -1516 550170 -1448 550226
rect -1392 550170 -1296 550226
rect -1916 550102 -1296 550170
rect -1916 550046 -1820 550102
rect -1764 550046 -1696 550102
rect -1640 550046 -1572 550102
rect -1516 550046 -1448 550102
rect -1392 550046 -1296 550102
rect -1916 549978 -1296 550046
rect -1916 549922 -1820 549978
rect -1764 549922 -1696 549978
rect -1640 549922 -1572 549978
rect -1516 549922 -1448 549978
rect -1392 549922 -1296 549978
rect -1916 532350 -1296 549922
rect -1916 532294 -1820 532350
rect -1764 532294 -1696 532350
rect -1640 532294 -1572 532350
rect -1516 532294 -1448 532350
rect -1392 532294 -1296 532350
rect -1916 532226 -1296 532294
rect -1916 532170 -1820 532226
rect -1764 532170 -1696 532226
rect -1640 532170 -1572 532226
rect -1516 532170 -1448 532226
rect -1392 532170 -1296 532226
rect -1916 532102 -1296 532170
rect -1916 532046 -1820 532102
rect -1764 532046 -1696 532102
rect -1640 532046 -1572 532102
rect -1516 532046 -1448 532102
rect -1392 532046 -1296 532102
rect -1916 531978 -1296 532046
rect -1916 531922 -1820 531978
rect -1764 531922 -1696 531978
rect -1640 531922 -1572 531978
rect -1516 531922 -1448 531978
rect -1392 531922 -1296 531978
rect -1916 514350 -1296 531922
rect -1916 514294 -1820 514350
rect -1764 514294 -1696 514350
rect -1640 514294 -1572 514350
rect -1516 514294 -1448 514350
rect -1392 514294 -1296 514350
rect -1916 514226 -1296 514294
rect -1916 514170 -1820 514226
rect -1764 514170 -1696 514226
rect -1640 514170 -1572 514226
rect -1516 514170 -1448 514226
rect -1392 514170 -1296 514226
rect -1916 514102 -1296 514170
rect -1916 514046 -1820 514102
rect -1764 514046 -1696 514102
rect -1640 514046 -1572 514102
rect -1516 514046 -1448 514102
rect -1392 514046 -1296 514102
rect -1916 513978 -1296 514046
rect -1916 513922 -1820 513978
rect -1764 513922 -1696 513978
rect -1640 513922 -1572 513978
rect -1516 513922 -1448 513978
rect -1392 513922 -1296 513978
rect -1916 496350 -1296 513922
rect -1916 496294 -1820 496350
rect -1764 496294 -1696 496350
rect -1640 496294 -1572 496350
rect -1516 496294 -1448 496350
rect -1392 496294 -1296 496350
rect -1916 496226 -1296 496294
rect -1916 496170 -1820 496226
rect -1764 496170 -1696 496226
rect -1640 496170 -1572 496226
rect -1516 496170 -1448 496226
rect -1392 496170 -1296 496226
rect -1916 496102 -1296 496170
rect -1916 496046 -1820 496102
rect -1764 496046 -1696 496102
rect -1640 496046 -1572 496102
rect -1516 496046 -1448 496102
rect -1392 496046 -1296 496102
rect -1916 495978 -1296 496046
rect -1916 495922 -1820 495978
rect -1764 495922 -1696 495978
rect -1640 495922 -1572 495978
rect -1516 495922 -1448 495978
rect -1392 495922 -1296 495978
rect -1916 478350 -1296 495922
rect -1916 478294 -1820 478350
rect -1764 478294 -1696 478350
rect -1640 478294 -1572 478350
rect -1516 478294 -1448 478350
rect -1392 478294 -1296 478350
rect -1916 478226 -1296 478294
rect -1916 478170 -1820 478226
rect -1764 478170 -1696 478226
rect -1640 478170 -1572 478226
rect -1516 478170 -1448 478226
rect -1392 478170 -1296 478226
rect -1916 478102 -1296 478170
rect -1916 478046 -1820 478102
rect -1764 478046 -1696 478102
rect -1640 478046 -1572 478102
rect -1516 478046 -1448 478102
rect -1392 478046 -1296 478102
rect -1916 477978 -1296 478046
rect -1916 477922 -1820 477978
rect -1764 477922 -1696 477978
rect -1640 477922 -1572 477978
rect -1516 477922 -1448 477978
rect -1392 477922 -1296 477978
rect -1916 460350 -1296 477922
rect -1916 460294 -1820 460350
rect -1764 460294 -1696 460350
rect -1640 460294 -1572 460350
rect -1516 460294 -1448 460350
rect -1392 460294 -1296 460350
rect -1916 460226 -1296 460294
rect -1916 460170 -1820 460226
rect -1764 460170 -1696 460226
rect -1640 460170 -1572 460226
rect -1516 460170 -1448 460226
rect -1392 460170 -1296 460226
rect -1916 460102 -1296 460170
rect -1916 460046 -1820 460102
rect -1764 460046 -1696 460102
rect -1640 460046 -1572 460102
rect -1516 460046 -1448 460102
rect -1392 460046 -1296 460102
rect -1916 459978 -1296 460046
rect -1916 459922 -1820 459978
rect -1764 459922 -1696 459978
rect -1640 459922 -1572 459978
rect -1516 459922 -1448 459978
rect -1392 459922 -1296 459978
rect -1916 442350 -1296 459922
rect -1916 442294 -1820 442350
rect -1764 442294 -1696 442350
rect -1640 442294 -1572 442350
rect -1516 442294 -1448 442350
rect -1392 442294 -1296 442350
rect -1916 442226 -1296 442294
rect -1916 442170 -1820 442226
rect -1764 442170 -1696 442226
rect -1640 442170 -1572 442226
rect -1516 442170 -1448 442226
rect -1392 442170 -1296 442226
rect -1916 442102 -1296 442170
rect -1916 442046 -1820 442102
rect -1764 442046 -1696 442102
rect -1640 442046 -1572 442102
rect -1516 442046 -1448 442102
rect -1392 442046 -1296 442102
rect -1916 441978 -1296 442046
rect -1916 441922 -1820 441978
rect -1764 441922 -1696 441978
rect -1640 441922 -1572 441978
rect -1516 441922 -1448 441978
rect -1392 441922 -1296 441978
rect -1916 424350 -1296 441922
rect -1916 424294 -1820 424350
rect -1764 424294 -1696 424350
rect -1640 424294 -1572 424350
rect -1516 424294 -1448 424350
rect -1392 424294 -1296 424350
rect -1916 424226 -1296 424294
rect -1916 424170 -1820 424226
rect -1764 424170 -1696 424226
rect -1640 424170 -1572 424226
rect -1516 424170 -1448 424226
rect -1392 424170 -1296 424226
rect -1916 424102 -1296 424170
rect -1916 424046 -1820 424102
rect -1764 424046 -1696 424102
rect -1640 424046 -1572 424102
rect -1516 424046 -1448 424102
rect -1392 424046 -1296 424102
rect -1916 423978 -1296 424046
rect -1916 423922 -1820 423978
rect -1764 423922 -1696 423978
rect -1640 423922 -1572 423978
rect -1516 423922 -1448 423978
rect -1392 423922 -1296 423978
rect -1916 406350 -1296 423922
rect -1916 406294 -1820 406350
rect -1764 406294 -1696 406350
rect -1640 406294 -1572 406350
rect -1516 406294 -1448 406350
rect -1392 406294 -1296 406350
rect -1916 406226 -1296 406294
rect -1916 406170 -1820 406226
rect -1764 406170 -1696 406226
rect -1640 406170 -1572 406226
rect -1516 406170 -1448 406226
rect -1392 406170 -1296 406226
rect -1916 406102 -1296 406170
rect -1916 406046 -1820 406102
rect -1764 406046 -1696 406102
rect -1640 406046 -1572 406102
rect -1516 406046 -1448 406102
rect -1392 406046 -1296 406102
rect -1916 405978 -1296 406046
rect -1916 405922 -1820 405978
rect -1764 405922 -1696 405978
rect -1640 405922 -1572 405978
rect -1516 405922 -1448 405978
rect -1392 405922 -1296 405978
rect -1916 388350 -1296 405922
rect -1916 388294 -1820 388350
rect -1764 388294 -1696 388350
rect -1640 388294 -1572 388350
rect -1516 388294 -1448 388350
rect -1392 388294 -1296 388350
rect -1916 388226 -1296 388294
rect -1916 388170 -1820 388226
rect -1764 388170 -1696 388226
rect -1640 388170 -1572 388226
rect -1516 388170 -1448 388226
rect -1392 388170 -1296 388226
rect -1916 388102 -1296 388170
rect -1916 388046 -1820 388102
rect -1764 388046 -1696 388102
rect -1640 388046 -1572 388102
rect -1516 388046 -1448 388102
rect -1392 388046 -1296 388102
rect -1916 387978 -1296 388046
rect -1916 387922 -1820 387978
rect -1764 387922 -1696 387978
rect -1640 387922 -1572 387978
rect -1516 387922 -1448 387978
rect -1392 387922 -1296 387978
rect -1916 370350 -1296 387922
rect -1916 370294 -1820 370350
rect -1764 370294 -1696 370350
rect -1640 370294 -1572 370350
rect -1516 370294 -1448 370350
rect -1392 370294 -1296 370350
rect -1916 370226 -1296 370294
rect -1916 370170 -1820 370226
rect -1764 370170 -1696 370226
rect -1640 370170 -1572 370226
rect -1516 370170 -1448 370226
rect -1392 370170 -1296 370226
rect -1916 370102 -1296 370170
rect -1916 370046 -1820 370102
rect -1764 370046 -1696 370102
rect -1640 370046 -1572 370102
rect -1516 370046 -1448 370102
rect -1392 370046 -1296 370102
rect -1916 369978 -1296 370046
rect -1916 369922 -1820 369978
rect -1764 369922 -1696 369978
rect -1640 369922 -1572 369978
rect -1516 369922 -1448 369978
rect -1392 369922 -1296 369978
rect -1916 352350 -1296 369922
rect -1916 352294 -1820 352350
rect -1764 352294 -1696 352350
rect -1640 352294 -1572 352350
rect -1516 352294 -1448 352350
rect -1392 352294 -1296 352350
rect -1916 352226 -1296 352294
rect -1916 352170 -1820 352226
rect -1764 352170 -1696 352226
rect -1640 352170 -1572 352226
rect -1516 352170 -1448 352226
rect -1392 352170 -1296 352226
rect -1916 352102 -1296 352170
rect -1916 352046 -1820 352102
rect -1764 352046 -1696 352102
rect -1640 352046 -1572 352102
rect -1516 352046 -1448 352102
rect -1392 352046 -1296 352102
rect -1916 351978 -1296 352046
rect -1916 351922 -1820 351978
rect -1764 351922 -1696 351978
rect -1640 351922 -1572 351978
rect -1516 351922 -1448 351978
rect -1392 351922 -1296 351978
rect -1916 334350 -1296 351922
rect -1916 334294 -1820 334350
rect -1764 334294 -1696 334350
rect -1640 334294 -1572 334350
rect -1516 334294 -1448 334350
rect -1392 334294 -1296 334350
rect -1916 334226 -1296 334294
rect -1916 334170 -1820 334226
rect -1764 334170 -1696 334226
rect -1640 334170 -1572 334226
rect -1516 334170 -1448 334226
rect -1392 334170 -1296 334226
rect -1916 334102 -1296 334170
rect -1916 334046 -1820 334102
rect -1764 334046 -1696 334102
rect -1640 334046 -1572 334102
rect -1516 334046 -1448 334102
rect -1392 334046 -1296 334102
rect -1916 333978 -1296 334046
rect -1916 333922 -1820 333978
rect -1764 333922 -1696 333978
rect -1640 333922 -1572 333978
rect -1516 333922 -1448 333978
rect -1392 333922 -1296 333978
rect -1916 316350 -1296 333922
rect -1916 316294 -1820 316350
rect -1764 316294 -1696 316350
rect -1640 316294 -1572 316350
rect -1516 316294 -1448 316350
rect -1392 316294 -1296 316350
rect -1916 316226 -1296 316294
rect -1916 316170 -1820 316226
rect -1764 316170 -1696 316226
rect -1640 316170 -1572 316226
rect -1516 316170 -1448 316226
rect -1392 316170 -1296 316226
rect -1916 316102 -1296 316170
rect -1916 316046 -1820 316102
rect -1764 316046 -1696 316102
rect -1640 316046 -1572 316102
rect -1516 316046 -1448 316102
rect -1392 316046 -1296 316102
rect -1916 315978 -1296 316046
rect -1916 315922 -1820 315978
rect -1764 315922 -1696 315978
rect -1640 315922 -1572 315978
rect -1516 315922 -1448 315978
rect -1392 315922 -1296 315978
rect -1916 298350 -1296 315922
rect -1916 298294 -1820 298350
rect -1764 298294 -1696 298350
rect -1640 298294 -1572 298350
rect -1516 298294 -1448 298350
rect -1392 298294 -1296 298350
rect -1916 298226 -1296 298294
rect -1916 298170 -1820 298226
rect -1764 298170 -1696 298226
rect -1640 298170 -1572 298226
rect -1516 298170 -1448 298226
rect -1392 298170 -1296 298226
rect -1916 298102 -1296 298170
rect -1916 298046 -1820 298102
rect -1764 298046 -1696 298102
rect -1640 298046 -1572 298102
rect -1516 298046 -1448 298102
rect -1392 298046 -1296 298102
rect -1916 297978 -1296 298046
rect -1916 297922 -1820 297978
rect -1764 297922 -1696 297978
rect -1640 297922 -1572 297978
rect -1516 297922 -1448 297978
rect -1392 297922 -1296 297978
rect -1916 280350 -1296 297922
rect -1916 280294 -1820 280350
rect -1764 280294 -1696 280350
rect -1640 280294 -1572 280350
rect -1516 280294 -1448 280350
rect -1392 280294 -1296 280350
rect -1916 280226 -1296 280294
rect -1916 280170 -1820 280226
rect -1764 280170 -1696 280226
rect -1640 280170 -1572 280226
rect -1516 280170 -1448 280226
rect -1392 280170 -1296 280226
rect -1916 280102 -1296 280170
rect -1916 280046 -1820 280102
rect -1764 280046 -1696 280102
rect -1640 280046 -1572 280102
rect -1516 280046 -1448 280102
rect -1392 280046 -1296 280102
rect -1916 279978 -1296 280046
rect -1916 279922 -1820 279978
rect -1764 279922 -1696 279978
rect -1640 279922 -1572 279978
rect -1516 279922 -1448 279978
rect -1392 279922 -1296 279978
rect -1916 262350 -1296 279922
rect -1916 262294 -1820 262350
rect -1764 262294 -1696 262350
rect -1640 262294 -1572 262350
rect -1516 262294 -1448 262350
rect -1392 262294 -1296 262350
rect -1916 262226 -1296 262294
rect -1916 262170 -1820 262226
rect -1764 262170 -1696 262226
rect -1640 262170 -1572 262226
rect -1516 262170 -1448 262226
rect -1392 262170 -1296 262226
rect -1916 262102 -1296 262170
rect -1916 262046 -1820 262102
rect -1764 262046 -1696 262102
rect -1640 262046 -1572 262102
rect -1516 262046 -1448 262102
rect -1392 262046 -1296 262102
rect -1916 261978 -1296 262046
rect -1916 261922 -1820 261978
rect -1764 261922 -1696 261978
rect -1640 261922 -1572 261978
rect -1516 261922 -1448 261978
rect -1392 261922 -1296 261978
rect -1916 244350 -1296 261922
rect -1916 244294 -1820 244350
rect -1764 244294 -1696 244350
rect -1640 244294 -1572 244350
rect -1516 244294 -1448 244350
rect -1392 244294 -1296 244350
rect -1916 244226 -1296 244294
rect -1916 244170 -1820 244226
rect -1764 244170 -1696 244226
rect -1640 244170 -1572 244226
rect -1516 244170 -1448 244226
rect -1392 244170 -1296 244226
rect -1916 244102 -1296 244170
rect -1916 244046 -1820 244102
rect -1764 244046 -1696 244102
rect -1640 244046 -1572 244102
rect -1516 244046 -1448 244102
rect -1392 244046 -1296 244102
rect -1916 243978 -1296 244046
rect -1916 243922 -1820 243978
rect -1764 243922 -1696 243978
rect -1640 243922 -1572 243978
rect -1516 243922 -1448 243978
rect -1392 243922 -1296 243978
rect -1916 226350 -1296 243922
rect -1916 226294 -1820 226350
rect -1764 226294 -1696 226350
rect -1640 226294 -1572 226350
rect -1516 226294 -1448 226350
rect -1392 226294 -1296 226350
rect -1916 226226 -1296 226294
rect -1916 226170 -1820 226226
rect -1764 226170 -1696 226226
rect -1640 226170 -1572 226226
rect -1516 226170 -1448 226226
rect -1392 226170 -1296 226226
rect -1916 226102 -1296 226170
rect -1916 226046 -1820 226102
rect -1764 226046 -1696 226102
rect -1640 226046 -1572 226102
rect -1516 226046 -1448 226102
rect -1392 226046 -1296 226102
rect -1916 225978 -1296 226046
rect -1916 225922 -1820 225978
rect -1764 225922 -1696 225978
rect -1640 225922 -1572 225978
rect -1516 225922 -1448 225978
rect -1392 225922 -1296 225978
rect -1916 208350 -1296 225922
rect -1916 208294 -1820 208350
rect -1764 208294 -1696 208350
rect -1640 208294 -1572 208350
rect -1516 208294 -1448 208350
rect -1392 208294 -1296 208350
rect -1916 208226 -1296 208294
rect -1916 208170 -1820 208226
rect -1764 208170 -1696 208226
rect -1640 208170 -1572 208226
rect -1516 208170 -1448 208226
rect -1392 208170 -1296 208226
rect -1916 208102 -1296 208170
rect -1916 208046 -1820 208102
rect -1764 208046 -1696 208102
rect -1640 208046 -1572 208102
rect -1516 208046 -1448 208102
rect -1392 208046 -1296 208102
rect -1916 207978 -1296 208046
rect -1916 207922 -1820 207978
rect -1764 207922 -1696 207978
rect -1640 207922 -1572 207978
rect -1516 207922 -1448 207978
rect -1392 207922 -1296 207978
rect -1916 190350 -1296 207922
rect -1916 190294 -1820 190350
rect -1764 190294 -1696 190350
rect -1640 190294 -1572 190350
rect -1516 190294 -1448 190350
rect -1392 190294 -1296 190350
rect -1916 190226 -1296 190294
rect -1916 190170 -1820 190226
rect -1764 190170 -1696 190226
rect -1640 190170 -1572 190226
rect -1516 190170 -1448 190226
rect -1392 190170 -1296 190226
rect -1916 190102 -1296 190170
rect -1916 190046 -1820 190102
rect -1764 190046 -1696 190102
rect -1640 190046 -1572 190102
rect -1516 190046 -1448 190102
rect -1392 190046 -1296 190102
rect -1916 189978 -1296 190046
rect -1916 189922 -1820 189978
rect -1764 189922 -1696 189978
rect -1640 189922 -1572 189978
rect -1516 189922 -1448 189978
rect -1392 189922 -1296 189978
rect -1916 172350 -1296 189922
rect -1916 172294 -1820 172350
rect -1764 172294 -1696 172350
rect -1640 172294 -1572 172350
rect -1516 172294 -1448 172350
rect -1392 172294 -1296 172350
rect -1916 172226 -1296 172294
rect -1916 172170 -1820 172226
rect -1764 172170 -1696 172226
rect -1640 172170 -1572 172226
rect -1516 172170 -1448 172226
rect -1392 172170 -1296 172226
rect -1916 172102 -1296 172170
rect -1916 172046 -1820 172102
rect -1764 172046 -1696 172102
rect -1640 172046 -1572 172102
rect -1516 172046 -1448 172102
rect -1392 172046 -1296 172102
rect -1916 171978 -1296 172046
rect -1916 171922 -1820 171978
rect -1764 171922 -1696 171978
rect -1640 171922 -1572 171978
rect -1516 171922 -1448 171978
rect -1392 171922 -1296 171978
rect -1916 154350 -1296 171922
rect -1916 154294 -1820 154350
rect -1764 154294 -1696 154350
rect -1640 154294 -1572 154350
rect -1516 154294 -1448 154350
rect -1392 154294 -1296 154350
rect -1916 154226 -1296 154294
rect -1916 154170 -1820 154226
rect -1764 154170 -1696 154226
rect -1640 154170 -1572 154226
rect -1516 154170 -1448 154226
rect -1392 154170 -1296 154226
rect -1916 154102 -1296 154170
rect -1916 154046 -1820 154102
rect -1764 154046 -1696 154102
rect -1640 154046 -1572 154102
rect -1516 154046 -1448 154102
rect -1392 154046 -1296 154102
rect -1916 153978 -1296 154046
rect -1916 153922 -1820 153978
rect -1764 153922 -1696 153978
rect -1640 153922 -1572 153978
rect -1516 153922 -1448 153978
rect -1392 153922 -1296 153978
rect -1916 136350 -1296 153922
rect -1916 136294 -1820 136350
rect -1764 136294 -1696 136350
rect -1640 136294 -1572 136350
rect -1516 136294 -1448 136350
rect -1392 136294 -1296 136350
rect -1916 136226 -1296 136294
rect -1916 136170 -1820 136226
rect -1764 136170 -1696 136226
rect -1640 136170 -1572 136226
rect -1516 136170 -1448 136226
rect -1392 136170 -1296 136226
rect -1916 136102 -1296 136170
rect -1916 136046 -1820 136102
rect -1764 136046 -1696 136102
rect -1640 136046 -1572 136102
rect -1516 136046 -1448 136102
rect -1392 136046 -1296 136102
rect -1916 135978 -1296 136046
rect -1916 135922 -1820 135978
rect -1764 135922 -1696 135978
rect -1640 135922 -1572 135978
rect -1516 135922 -1448 135978
rect -1392 135922 -1296 135978
rect -1916 118350 -1296 135922
rect -1916 118294 -1820 118350
rect -1764 118294 -1696 118350
rect -1640 118294 -1572 118350
rect -1516 118294 -1448 118350
rect -1392 118294 -1296 118350
rect -1916 118226 -1296 118294
rect -1916 118170 -1820 118226
rect -1764 118170 -1696 118226
rect -1640 118170 -1572 118226
rect -1516 118170 -1448 118226
rect -1392 118170 -1296 118226
rect -1916 118102 -1296 118170
rect -1916 118046 -1820 118102
rect -1764 118046 -1696 118102
rect -1640 118046 -1572 118102
rect -1516 118046 -1448 118102
rect -1392 118046 -1296 118102
rect -1916 117978 -1296 118046
rect -1916 117922 -1820 117978
rect -1764 117922 -1696 117978
rect -1640 117922 -1572 117978
rect -1516 117922 -1448 117978
rect -1392 117922 -1296 117978
rect -1916 100350 -1296 117922
rect -1916 100294 -1820 100350
rect -1764 100294 -1696 100350
rect -1640 100294 -1572 100350
rect -1516 100294 -1448 100350
rect -1392 100294 -1296 100350
rect -1916 100226 -1296 100294
rect -1916 100170 -1820 100226
rect -1764 100170 -1696 100226
rect -1640 100170 -1572 100226
rect -1516 100170 -1448 100226
rect -1392 100170 -1296 100226
rect -1916 100102 -1296 100170
rect -1916 100046 -1820 100102
rect -1764 100046 -1696 100102
rect -1640 100046 -1572 100102
rect -1516 100046 -1448 100102
rect -1392 100046 -1296 100102
rect -1916 99978 -1296 100046
rect -1916 99922 -1820 99978
rect -1764 99922 -1696 99978
rect -1640 99922 -1572 99978
rect -1516 99922 -1448 99978
rect -1392 99922 -1296 99978
rect -1916 82350 -1296 99922
rect -1916 82294 -1820 82350
rect -1764 82294 -1696 82350
rect -1640 82294 -1572 82350
rect -1516 82294 -1448 82350
rect -1392 82294 -1296 82350
rect -1916 82226 -1296 82294
rect -1916 82170 -1820 82226
rect -1764 82170 -1696 82226
rect -1640 82170 -1572 82226
rect -1516 82170 -1448 82226
rect -1392 82170 -1296 82226
rect -1916 82102 -1296 82170
rect -1916 82046 -1820 82102
rect -1764 82046 -1696 82102
rect -1640 82046 -1572 82102
rect -1516 82046 -1448 82102
rect -1392 82046 -1296 82102
rect -1916 81978 -1296 82046
rect -1916 81922 -1820 81978
rect -1764 81922 -1696 81978
rect -1640 81922 -1572 81978
rect -1516 81922 -1448 81978
rect -1392 81922 -1296 81978
rect -1916 64350 -1296 81922
rect -1916 64294 -1820 64350
rect -1764 64294 -1696 64350
rect -1640 64294 -1572 64350
rect -1516 64294 -1448 64350
rect -1392 64294 -1296 64350
rect -1916 64226 -1296 64294
rect -1916 64170 -1820 64226
rect -1764 64170 -1696 64226
rect -1640 64170 -1572 64226
rect -1516 64170 -1448 64226
rect -1392 64170 -1296 64226
rect -1916 64102 -1296 64170
rect -1916 64046 -1820 64102
rect -1764 64046 -1696 64102
rect -1640 64046 -1572 64102
rect -1516 64046 -1448 64102
rect -1392 64046 -1296 64102
rect -1916 63978 -1296 64046
rect -1916 63922 -1820 63978
rect -1764 63922 -1696 63978
rect -1640 63922 -1572 63978
rect -1516 63922 -1448 63978
rect -1392 63922 -1296 63978
rect -1916 46350 -1296 63922
rect -1916 46294 -1820 46350
rect -1764 46294 -1696 46350
rect -1640 46294 -1572 46350
rect -1516 46294 -1448 46350
rect -1392 46294 -1296 46350
rect -1916 46226 -1296 46294
rect -1916 46170 -1820 46226
rect -1764 46170 -1696 46226
rect -1640 46170 -1572 46226
rect -1516 46170 -1448 46226
rect -1392 46170 -1296 46226
rect -1916 46102 -1296 46170
rect -1916 46046 -1820 46102
rect -1764 46046 -1696 46102
rect -1640 46046 -1572 46102
rect -1516 46046 -1448 46102
rect -1392 46046 -1296 46102
rect -1916 45978 -1296 46046
rect -1916 45922 -1820 45978
rect -1764 45922 -1696 45978
rect -1640 45922 -1572 45978
rect -1516 45922 -1448 45978
rect -1392 45922 -1296 45978
rect -1916 28350 -1296 45922
rect -1916 28294 -1820 28350
rect -1764 28294 -1696 28350
rect -1640 28294 -1572 28350
rect -1516 28294 -1448 28350
rect -1392 28294 -1296 28350
rect -1916 28226 -1296 28294
rect -1916 28170 -1820 28226
rect -1764 28170 -1696 28226
rect -1640 28170 -1572 28226
rect -1516 28170 -1448 28226
rect -1392 28170 -1296 28226
rect -1916 28102 -1296 28170
rect -1916 28046 -1820 28102
rect -1764 28046 -1696 28102
rect -1640 28046 -1572 28102
rect -1516 28046 -1448 28102
rect -1392 28046 -1296 28102
rect -1916 27978 -1296 28046
rect -1916 27922 -1820 27978
rect -1764 27922 -1696 27978
rect -1640 27922 -1572 27978
rect -1516 27922 -1448 27978
rect -1392 27922 -1296 27978
rect -1916 10350 -1296 27922
rect -1916 10294 -1820 10350
rect -1764 10294 -1696 10350
rect -1640 10294 -1572 10350
rect -1516 10294 -1448 10350
rect -1392 10294 -1296 10350
rect -1916 10226 -1296 10294
rect -1916 10170 -1820 10226
rect -1764 10170 -1696 10226
rect -1640 10170 -1572 10226
rect -1516 10170 -1448 10226
rect -1392 10170 -1296 10226
rect -1916 10102 -1296 10170
rect -1916 10046 -1820 10102
rect -1764 10046 -1696 10102
rect -1640 10046 -1572 10102
rect -1516 10046 -1448 10102
rect -1392 10046 -1296 10102
rect -1916 9978 -1296 10046
rect -1916 9922 -1820 9978
rect -1764 9922 -1696 9978
rect -1640 9922 -1572 9978
rect -1516 9922 -1448 9978
rect -1392 9922 -1296 9978
rect -1916 -1120 -1296 9922
rect -956 597212 -336 597308
rect -956 597156 -860 597212
rect -804 597156 -736 597212
rect -680 597156 -612 597212
rect -556 597156 -488 597212
rect -432 597156 -336 597212
rect -956 597088 -336 597156
rect -956 597032 -860 597088
rect -804 597032 -736 597088
rect -680 597032 -612 597088
rect -556 597032 -488 597088
rect -432 597032 -336 597088
rect -956 596964 -336 597032
rect -956 596908 -860 596964
rect -804 596908 -736 596964
rect -680 596908 -612 596964
rect -556 596908 -488 596964
rect -432 596908 -336 596964
rect -956 596840 -336 596908
rect -956 596784 -860 596840
rect -804 596784 -736 596840
rect -680 596784 -612 596840
rect -556 596784 -488 596840
rect -432 596784 -336 596840
rect -956 580350 -336 596784
rect 5418 597212 6038 598268
rect 5418 597156 5514 597212
rect 5570 597156 5638 597212
rect 5694 597156 5762 597212
rect 5818 597156 5886 597212
rect 5942 597156 6038 597212
rect 5418 597088 6038 597156
rect 5418 597032 5514 597088
rect 5570 597032 5638 597088
rect 5694 597032 5762 597088
rect 5818 597032 5886 597088
rect 5942 597032 6038 597088
rect 5418 596964 6038 597032
rect 5418 596908 5514 596964
rect 5570 596908 5638 596964
rect 5694 596908 5762 596964
rect 5818 596908 5886 596964
rect 5942 596908 6038 596964
rect 5418 596840 6038 596908
rect 5418 596784 5514 596840
rect 5570 596784 5638 596840
rect 5694 596784 5762 596840
rect 5818 596784 5886 596840
rect 5942 596784 6038 596840
rect -956 580294 -860 580350
rect -804 580294 -736 580350
rect -680 580294 -612 580350
rect -556 580294 -488 580350
rect -432 580294 -336 580350
rect -956 580226 -336 580294
rect -956 580170 -860 580226
rect -804 580170 -736 580226
rect -680 580170 -612 580226
rect -556 580170 -488 580226
rect -432 580170 -336 580226
rect -956 580102 -336 580170
rect -956 580046 -860 580102
rect -804 580046 -736 580102
rect -680 580046 -612 580102
rect -556 580046 -488 580102
rect -432 580046 -336 580102
rect -956 579978 -336 580046
rect -956 579922 -860 579978
rect -804 579922 -736 579978
rect -680 579922 -612 579978
rect -556 579922 -488 579978
rect -432 579922 -336 579978
rect -956 562350 -336 579922
rect 3388 587188 3444 587198
rect 3388 576118 3444 587132
rect -956 562294 -860 562350
rect -804 562294 -736 562350
rect -680 562294 -612 562350
rect -556 562294 -488 562350
rect -432 562294 -336 562350
rect -956 562226 -336 562294
rect -956 562170 -860 562226
rect -804 562170 -736 562226
rect -680 562170 -612 562226
rect -556 562170 -488 562226
rect -432 562170 -336 562226
rect -956 562102 -336 562170
rect -956 562046 -860 562102
rect -804 562046 -736 562102
rect -680 562046 -612 562102
rect -556 562046 -488 562102
rect -432 562046 -336 562102
rect -956 561978 -336 562046
rect -956 561922 -860 561978
rect -804 561922 -736 561978
rect -680 561922 -612 561978
rect -556 561922 -488 561978
rect -432 561922 -336 561978
rect -956 544350 -336 561922
rect 3276 576062 3444 576118
rect 5418 580350 6038 596784
rect 5418 580294 5514 580350
rect 5570 580294 5638 580350
rect 5694 580294 5762 580350
rect 5818 580294 5886 580350
rect 5942 580294 6038 580350
rect 5418 580226 6038 580294
rect 5418 580170 5514 580226
rect 5570 580170 5638 580226
rect 5694 580170 5762 580226
rect 5818 580170 5886 580226
rect 5942 580170 6038 580226
rect 5418 580102 6038 580170
rect 5418 580046 5514 580102
rect 5570 580046 5638 580102
rect 5694 580046 5762 580102
rect 5818 580046 5886 580102
rect 5942 580046 6038 580102
rect 5418 579978 6038 580046
rect 5418 579922 5514 579978
rect 5570 579922 5638 579978
rect 5694 579922 5762 579978
rect 5818 579922 5886 579978
rect 5942 579922 6038 579978
rect -956 544294 -860 544350
rect -804 544294 -736 544350
rect -680 544294 -612 544350
rect -556 544294 -488 544350
rect -432 544294 -336 544350
rect -956 544226 -336 544294
rect -956 544170 -860 544226
rect -804 544170 -736 544226
rect -680 544170 -612 544226
rect -556 544170 -488 544226
rect -432 544170 -336 544226
rect -956 544102 -336 544170
rect -956 544046 -860 544102
rect -804 544046 -736 544102
rect -680 544046 -612 544102
rect -556 544046 -488 544102
rect -432 544046 -336 544102
rect -956 543978 -336 544046
rect -956 543922 -860 543978
rect -804 543922 -736 543978
rect -680 543922 -612 543978
rect -556 543922 -488 543978
rect -432 543922 -336 543978
rect -956 526350 -336 543922
rect -956 526294 -860 526350
rect -804 526294 -736 526350
rect -680 526294 -612 526350
rect -556 526294 -488 526350
rect -432 526294 -336 526350
rect -956 526226 -336 526294
rect -956 526170 -860 526226
rect -804 526170 -736 526226
rect -680 526170 -612 526226
rect -556 526170 -488 526226
rect -432 526170 -336 526226
rect -956 526102 -336 526170
rect -956 526046 -860 526102
rect -804 526046 -736 526102
rect -680 526046 -612 526102
rect -556 526046 -488 526102
rect -432 526046 -336 526102
rect -956 525978 -336 526046
rect -956 525922 -860 525978
rect -804 525922 -736 525978
rect -680 525922 -612 525978
rect -556 525922 -488 525978
rect -432 525922 -336 525978
rect -956 508350 -336 525922
rect -956 508294 -860 508350
rect -804 508294 -736 508350
rect -680 508294 -612 508350
rect -556 508294 -488 508350
rect -432 508294 -336 508350
rect -956 508226 -336 508294
rect -956 508170 -860 508226
rect -804 508170 -736 508226
rect -680 508170 -612 508226
rect -556 508170 -488 508226
rect -432 508170 -336 508226
rect -956 508102 -336 508170
rect -956 508046 -860 508102
rect -804 508046 -736 508102
rect -680 508046 -612 508102
rect -556 508046 -488 508102
rect -432 508046 -336 508102
rect -956 507978 -336 508046
rect -956 507922 -860 507978
rect -804 507922 -736 507978
rect -680 507922 -612 507978
rect -556 507922 -488 507978
rect -432 507922 -336 507978
rect -956 490350 -336 507922
rect -956 490294 -860 490350
rect -804 490294 -736 490350
rect -680 490294 -612 490350
rect -556 490294 -488 490350
rect -432 490294 -336 490350
rect -956 490226 -336 490294
rect -956 490170 -860 490226
rect -804 490170 -736 490226
rect -680 490170 -612 490226
rect -556 490170 -488 490226
rect -432 490170 -336 490226
rect -956 490102 -336 490170
rect -956 490046 -860 490102
rect -804 490046 -736 490102
rect -680 490046 -612 490102
rect -556 490046 -488 490102
rect -432 490046 -336 490102
rect -956 489978 -336 490046
rect -956 489922 -860 489978
rect -804 489922 -736 489978
rect -680 489922 -612 489978
rect -556 489922 -488 489978
rect -432 489922 -336 489978
rect -956 472350 -336 489922
rect -956 472294 -860 472350
rect -804 472294 -736 472350
rect -680 472294 -612 472350
rect -556 472294 -488 472350
rect -432 472294 -336 472350
rect -956 472226 -336 472294
rect -956 472170 -860 472226
rect -804 472170 -736 472226
rect -680 472170 -612 472226
rect -556 472170 -488 472226
rect -432 472170 -336 472226
rect -956 472102 -336 472170
rect -956 472046 -860 472102
rect -804 472046 -736 472102
rect -680 472046 -612 472102
rect -556 472046 -488 472102
rect -432 472046 -336 472102
rect -956 471978 -336 472046
rect -956 471922 -860 471978
rect -804 471922 -736 471978
rect -680 471922 -612 471978
rect -556 471922 -488 471978
rect -432 471922 -336 471978
rect -956 454350 -336 471922
rect -956 454294 -860 454350
rect -804 454294 -736 454350
rect -680 454294 -612 454350
rect -556 454294 -488 454350
rect -432 454294 -336 454350
rect -956 454226 -336 454294
rect -956 454170 -860 454226
rect -804 454170 -736 454226
rect -680 454170 -612 454226
rect -556 454170 -488 454226
rect -432 454170 -336 454226
rect -956 454102 -336 454170
rect -956 454046 -860 454102
rect -804 454046 -736 454102
rect -680 454046 -612 454102
rect -556 454046 -488 454102
rect -432 454046 -336 454102
rect -956 453978 -336 454046
rect -956 453922 -860 453978
rect -804 453922 -736 453978
rect -680 453922 -612 453978
rect -556 453922 -488 453978
rect -432 453922 -336 453978
rect -956 436350 -336 453922
rect -956 436294 -860 436350
rect -804 436294 -736 436350
rect -680 436294 -612 436350
rect -556 436294 -488 436350
rect -432 436294 -336 436350
rect -956 436226 -336 436294
rect -956 436170 -860 436226
rect -804 436170 -736 436226
rect -680 436170 -612 436226
rect -556 436170 -488 436226
rect -432 436170 -336 436226
rect -956 436102 -336 436170
rect -956 436046 -860 436102
rect -804 436046 -736 436102
rect -680 436046 -612 436102
rect -556 436046 -488 436102
rect -432 436046 -336 436102
rect -956 435978 -336 436046
rect -956 435922 -860 435978
rect -804 435922 -736 435978
rect -680 435922 -612 435978
rect -556 435922 -488 435978
rect -432 435922 -336 435978
rect -956 418350 -336 435922
rect -956 418294 -860 418350
rect -804 418294 -736 418350
rect -680 418294 -612 418350
rect -556 418294 -488 418350
rect -432 418294 -336 418350
rect -956 418226 -336 418294
rect -956 418170 -860 418226
rect -804 418170 -736 418226
rect -680 418170 -612 418226
rect -556 418170 -488 418226
rect -432 418170 -336 418226
rect -956 418102 -336 418170
rect -956 418046 -860 418102
rect -804 418046 -736 418102
rect -680 418046 -612 418102
rect -556 418046 -488 418102
rect -432 418046 -336 418102
rect -956 417978 -336 418046
rect -956 417922 -860 417978
rect -804 417922 -736 417978
rect -680 417922 -612 417978
rect -556 417922 -488 417978
rect -432 417922 -336 417978
rect -956 400350 -336 417922
rect -956 400294 -860 400350
rect -804 400294 -736 400350
rect -680 400294 -612 400350
rect -556 400294 -488 400350
rect -432 400294 -336 400350
rect -956 400226 -336 400294
rect -956 400170 -860 400226
rect -804 400170 -736 400226
rect -680 400170 -612 400226
rect -556 400170 -488 400226
rect -432 400170 -336 400226
rect -956 400102 -336 400170
rect -956 400046 -860 400102
rect -804 400046 -736 400102
rect -680 400046 -612 400102
rect -556 400046 -488 400102
rect -432 400046 -336 400102
rect -956 399978 -336 400046
rect -956 399922 -860 399978
rect -804 399922 -736 399978
rect -680 399922 -612 399978
rect -556 399922 -488 399978
rect -432 399922 -336 399978
rect -956 382350 -336 399922
rect -956 382294 -860 382350
rect -804 382294 -736 382350
rect -680 382294 -612 382350
rect -556 382294 -488 382350
rect -432 382294 -336 382350
rect -956 382226 -336 382294
rect -956 382170 -860 382226
rect -804 382170 -736 382226
rect -680 382170 -612 382226
rect -556 382170 -488 382226
rect -432 382170 -336 382226
rect -956 382102 -336 382170
rect -956 382046 -860 382102
rect -804 382046 -736 382102
rect -680 382046 -612 382102
rect -556 382046 -488 382102
rect -432 382046 -336 382102
rect -956 381978 -336 382046
rect -956 381922 -860 381978
rect -804 381922 -736 381978
rect -680 381922 -612 381978
rect -556 381922 -488 381978
rect -432 381922 -336 381978
rect -956 364350 -336 381922
rect -956 364294 -860 364350
rect -804 364294 -736 364350
rect -680 364294 -612 364350
rect -556 364294 -488 364350
rect -432 364294 -336 364350
rect -956 364226 -336 364294
rect -956 364170 -860 364226
rect -804 364170 -736 364226
rect -680 364170 -612 364226
rect -556 364170 -488 364226
rect -432 364170 -336 364226
rect -956 364102 -336 364170
rect -956 364046 -860 364102
rect -804 364046 -736 364102
rect -680 364046 -612 364102
rect -556 364046 -488 364102
rect -432 364046 -336 364102
rect -956 363978 -336 364046
rect -956 363922 -860 363978
rect -804 363922 -736 363978
rect -680 363922 -612 363978
rect -556 363922 -488 363978
rect -432 363922 -336 363978
rect -956 346350 -336 363922
rect -956 346294 -860 346350
rect -804 346294 -736 346350
rect -680 346294 -612 346350
rect -556 346294 -488 346350
rect -432 346294 -336 346350
rect -956 346226 -336 346294
rect -956 346170 -860 346226
rect -804 346170 -736 346226
rect -680 346170 -612 346226
rect -556 346170 -488 346226
rect -432 346170 -336 346226
rect -956 346102 -336 346170
rect -956 346046 -860 346102
rect -804 346046 -736 346102
rect -680 346046 -612 346102
rect -556 346046 -488 346102
rect -432 346046 -336 346102
rect -956 345978 -336 346046
rect -956 345922 -860 345978
rect -804 345922 -736 345978
rect -680 345922 -612 345978
rect -556 345922 -488 345978
rect -432 345922 -336 345978
rect -956 328350 -336 345922
rect -956 328294 -860 328350
rect -804 328294 -736 328350
rect -680 328294 -612 328350
rect -556 328294 -488 328350
rect -432 328294 -336 328350
rect -956 328226 -336 328294
rect -956 328170 -860 328226
rect -804 328170 -736 328226
rect -680 328170 -612 328226
rect -556 328170 -488 328226
rect -432 328170 -336 328226
rect -956 328102 -336 328170
rect -956 328046 -860 328102
rect -804 328046 -736 328102
rect -680 328046 -612 328102
rect -556 328046 -488 328102
rect -432 328046 -336 328102
rect -956 327978 -336 328046
rect -956 327922 -860 327978
rect -804 327922 -736 327978
rect -680 327922 -612 327978
rect -556 327922 -488 327978
rect -432 327922 -336 327978
rect -956 310350 -336 327922
rect -956 310294 -860 310350
rect -804 310294 -736 310350
rect -680 310294 -612 310350
rect -556 310294 -488 310350
rect -432 310294 -336 310350
rect -956 310226 -336 310294
rect -956 310170 -860 310226
rect -804 310170 -736 310226
rect -680 310170 -612 310226
rect -556 310170 -488 310226
rect -432 310170 -336 310226
rect -956 310102 -336 310170
rect -956 310046 -860 310102
rect -804 310046 -736 310102
rect -680 310046 -612 310102
rect -556 310046 -488 310102
rect -432 310046 -336 310102
rect -956 309978 -336 310046
rect -956 309922 -860 309978
rect -804 309922 -736 309978
rect -680 309922 -612 309978
rect -556 309922 -488 309978
rect -432 309922 -336 309978
rect -956 292350 -336 309922
rect -956 292294 -860 292350
rect -804 292294 -736 292350
rect -680 292294 -612 292350
rect -556 292294 -488 292350
rect -432 292294 -336 292350
rect -956 292226 -336 292294
rect -956 292170 -860 292226
rect -804 292170 -736 292226
rect -680 292170 -612 292226
rect -556 292170 -488 292226
rect -432 292170 -336 292226
rect -956 292102 -336 292170
rect -956 292046 -860 292102
rect -804 292046 -736 292102
rect -680 292046 -612 292102
rect -556 292046 -488 292102
rect -432 292046 -336 292102
rect -956 291978 -336 292046
rect -956 291922 -860 291978
rect -804 291922 -736 291978
rect -680 291922 -612 291978
rect -556 291922 -488 291978
rect -432 291922 -336 291978
rect -956 274350 -336 291922
rect -956 274294 -860 274350
rect -804 274294 -736 274350
rect -680 274294 -612 274350
rect -556 274294 -488 274350
rect -432 274294 -336 274350
rect -956 274226 -336 274294
rect -956 274170 -860 274226
rect -804 274170 -736 274226
rect -680 274170 -612 274226
rect -556 274170 -488 274226
rect -432 274170 -336 274226
rect -956 274102 -336 274170
rect -956 274046 -860 274102
rect -804 274046 -736 274102
rect -680 274046 -612 274102
rect -556 274046 -488 274102
rect -432 274046 -336 274102
rect -956 273978 -336 274046
rect -956 273922 -860 273978
rect -804 273922 -736 273978
rect -680 273922 -612 273978
rect -556 273922 -488 273978
rect -432 273922 -336 273978
rect -956 256350 -336 273922
rect -956 256294 -860 256350
rect -804 256294 -736 256350
rect -680 256294 -612 256350
rect -556 256294 -488 256350
rect -432 256294 -336 256350
rect -956 256226 -336 256294
rect -956 256170 -860 256226
rect -804 256170 -736 256226
rect -680 256170 -612 256226
rect -556 256170 -488 256226
rect -432 256170 -336 256226
rect -956 256102 -336 256170
rect -956 256046 -860 256102
rect -804 256046 -736 256102
rect -680 256046 -612 256102
rect -556 256046 -488 256102
rect -432 256046 -336 256102
rect -956 255978 -336 256046
rect -956 255922 -860 255978
rect -804 255922 -736 255978
rect -680 255922 -612 255978
rect -556 255922 -488 255978
rect -432 255922 -336 255978
rect -956 238350 -336 255922
rect -956 238294 -860 238350
rect -804 238294 -736 238350
rect -680 238294 -612 238350
rect -556 238294 -488 238350
rect -432 238294 -336 238350
rect -956 238226 -336 238294
rect -956 238170 -860 238226
rect -804 238170 -736 238226
rect -680 238170 -612 238226
rect -556 238170 -488 238226
rect -432 238170 -336 238226
rect -956 238102 -336 238170
rect -956 238046 -860 238102
rect -804 238046 -736 238102
rect -680 238046 -612 238102
rect -556 238046 -488 238102
rect -432 238046 -336 238102
rect -956 237978 -336 238046
rect -956 237922 -860 237978
rect -804 237922 -736 237978
rect -680 237922 -612 237978
rect -556 237922 -488 237978
rect -432 237922 -336 237978
rect -956 220350 -336 237922
rect -956 220294 -860 220350
rect -804 220294 -736 220350
rect -680 220294 -612 220350
rect -556 220294 -488 220350
rect -432 220294 -336 220350
rect -956 220226 -336 220294
rect -956 220170 -860 220226
rect -804 220170 -736 220226
rect -680 220170 -612 220226
rect -556 220170 -488 220226
rect -432 220170 -336 220226
rect -956 220102 -336 220170
rect -956 220046 -860 220102
rect -804 220046 -736 220102
rect -680 220046 -612 220102
rect -556 220046 -488 220102
rect -432 220046 -336 220102
rect -956 219978 -336 220046
rect -956 219922 -860 219978
rect -804 219922 -736 219978
rect -680 219922 -612 219978
rect -556 219922 -488 219978
rect -432 219922 -336 219978
rect -956 202350 -336 219922
rect -956 202294 -860 202350
rect -804 202294 -736 202350
rect -680 202294 -612 202350
rect -556 202294 -488 202350
rect -432 202294 -336 202350
rect -956 202226 -336 202294
rect -956 202170 -860 202226
rect -804 202170 -736 202226
rect -680 202170 -612 202226
rect -556 202170 -488 202226
rect -432 202170 -336 202226
rect -956 202102 -336 202170
rect -956 202046 -860 202102
rect -804 202046 -736 202102
rect -680 202046 -612 202102
rect -556 202046 -488 202102
rect -432 202046 -336 202102
rect -956 201978 -336 202046
rect -956 201922 -860 201978
rect -804 201922 -736 201978
rect -680 201922 -612 201978
rect -556 201922 -488 201978
rect -432 201922 -336 201978
rect -956 184350 -336 201922
rect -956 184294 -860 184350
rect -804 184294 -736 184350
rect -680 184294 -612 184350
rect -556 184294 -488 184350
rect -432 184294 -336 184350
rect -956 184226 -336 184294
rect -956 184170 -860 184226
rect -804 184170 -736 184226
rect -680 184170 -612 184226
rect -556 184170 -488 184226
rect -432 184170 -336 184226
rect -956 184102 -336 184170
rect -956 184046 -860 184102
rect -804 184046 -736 184102
rect -680 184046 -612 184102
rect -556 184046 -488 184102
rect -432 184046 -336 184102
rect -956 183978 -336 184046
rect -956 183922 -860 183978
rect -804 183922 -736 183978
rect -680 183922 -612 183978
rect -556 183922 -488 183978
rect -432 183922 -336 183978
rect -956 166350 -336 183922
rect -956 166294 -860 166350
rect -804 166294 -736 166350
rect -680 166294 -612 166350
rect -556 166294 -488 166350
rect -432 166294 -336 166350
rect -956 166226 -336 166294
rect -956 166170 -860 166226
rect -804 166170 -736 166226
rect -680 166170 -612 166226
rect -556 166170 -488 166226
rect -432 166170 -336 166226
rect -956 166102 -336 166170
rect -956 166046 -860 166102
rect -804 166046 -736 166102
rect -680 166046 -612 166102
rect -556 166046 -488 166102
rect -432 166046 -336 166102
rect -956 165978 -336 166046
rect -956 165922 -860 165978
rect -804 165922 -736 165978
rect -680 165922 -612 165978
rect -556 165922 -488 165978
rect -432 165922 -336 165978
rect -956 148350 -336 165922
rect -956 148294 -860 148350
rect -804 148294 -736 148350
rect -680 148294 -612 148350
rect -556 148294 -488 148350
rect -432 148294 -336 148350
rect -956 148226 -336 148294
rect -956 148170 -860 148226
rect -804 148170 -736 148226
rect -680 148170 -612 148226
rect -556 148170 -488 148226
rect -432 148170 -336 148226
rect -956 148102 -336 148170
rect -956 148046 -860 148102
rect -804 148046 -736 148102
rect -680 148046 -612 148102
rect -556 148046 -488 148102
rect -432 148046 -336 148102
rect -956 147978 -336 148046
rect -956 147922 -860 147978
rect -804 147922 -736 147978
rect -680 147922 -612 147978
rect -556 147922 -488 147978
rect -432 147922 -336 147978
rect -956 130350 -336 147922
rect -956 130294 -860 130350
rect -804 130294 -736 130350
rect -680 130294 -612 130350
rect -556 130294 -488 130350
rect -432 130294 -336 130350
rect -956 130226 -336 130294
rect -956 130170 -860 130226
rect -804 130170 -736 130226
rect -680 130170 -612 130226
rect -556 130170 -488 130226
rect -432 130170 -336 130226
rect -956 130102 -336 130170
rect -956 130046 -860 130102
rect -804 130046 -736 130102
rect -680 130046 -612 130102
rect -556 130046 -488 130102
rect -432 130046 -336 130102
rect -956 129978 -336 130046
rect -956 129922 -860 129978
rect -804 129922 -736 129978
rect -680 129922 -612 129978
rect -556 129922 -488 129978
rect -432 129922 -336 129978
rect -956 112350 -336 129922
rect -956 112294 -860 112350
rect -804 112294 -736 112350
rect -680 112294 -612 112350
rect -556 112294 -488 112350
rect -432 112294 -336 112350
rect -956 112226 -336 112294
rect -956 112170 -860 112226
rect -804 112170 -736 112226
rect -680 112170 -612 112226
rect -556 112170 -488 112226
rect -432 112170 -336 112226
rect -956 112102 -336 112170
rect -956 112046 -860 112102
rect -804 112046 -736 112102
rect -680 112046 -612 112102
rect -556 112046 -488 112102
rect -432 112046 -336 112102
rect -956 111978 -336 112046
rect -956 111922 -860 111978
rect -804 111922 -736 111978
rect -680 111922 -612 111978
rect -556 111922 -488 111978
rect -432 111922 -336 111978
rect -956 94350 -336 111922
rect -956 94294 -860 94350
rect -804 94294 -736 94350
rect -680 94294 -612 94350
rect -556 94294 -488 94350
rect -432 94294 -336 94350
rect -956 94226 -336 94294
rect -956 94170 -860 94226
rect -804 94170 -736 94226
rect -680 94170 -612 94226
rect -556 94170 -488 94226
rect -432 94170 -336 94226
rect -956 94102 -336 94170
rect -956 94046 -860 94102
rect -804 94046 -736 94102
rect -680 94046 -612 94102
rect -556 94046 -488 94102
rect -432 94046 -336 94102
rect -956 93978 -336 94046
rect -956 93922 -860 93978
rect -804 93922 -736 93978
rect -680 93922 -612 93978
rect -556 93922 -488 93978
rect -432 93922 -336 93978
rect -956 76350 -336 93922
rect -956 76294 -860 76350
rect -804 76294 -736 76350
rect -680 76294 -612 76350
rect -556 76294 -488 76350
rect -432 76294 -336 76350
rect -956 76226 -336 76294
rect -956 76170 -860 76226
rect -804 76170 -736 76226
rect -680 76170 -612 76226
rect -556 76170 -488 76226
rect -432 76170 -336 76226
rect -956 76102 -336 76170
rect -956 76046 -860 76102
rect -804 76046 -736 76102
rect -680 76046 -612 76102
rect -556 76046 -488 76102
rect -432 76046 -336 76102
rect -956 75978 -336 76046
rect -956 75922 -860 75978
rect -804 75922 -736 75978
rect -680 75922 -612 75978
rect -556 75922 -488 75978
rect -432 75922 -336 75978
rect -956 58350 -336 75922
rect -956 58294 -860 58350
rect -804 58294 -736 58350
rect -680 58294 -612 58350
rect -556 58294 -488 58350
rect -432 58294 -336 58350
rect -956 58226 -336 58294
rect -956 58170 -860 58226
rect -804 58170 -736 58226
rect -680 58170 -612 58226
rect -556 58170 -488 58226
rect -432 58170 -336 58226
rect -956 58102 -336 58170
rect -956 58046 -860 58102
rect -804 58046 -736 58102
rect -680 58046 -612 58102
rect -556 58046 -488 58102
rect -432 58046 -336 58102
rect -956 57978 -336 58046
rect -956 57922 -860 57978
rect -804 57922 -736 57978
rect -680 57922 -612 57978
rect -556 57922 -488 57978
rect -432 57922 -336 57978
rect -956 40350 -336 57922
rect -956 40294 -860 40350
rect -804 40294 -736 40350
rect -680 40294 -612 40350
rect -556 40294 -488 40350
rect -432 40294 -336 40350
rect -956 40226 -336 40294
rect -956 40170 -860 40226
rect -804 40170 -736 40226
rect -680 40170 -612 40226
rect -556 40170 -488 40226
rect -432 40170 -336 40226
rect -956 40102 -336 40170
rect -956 40046 -860 40102
rect -804 40046 -736 40102
rect -680 40046 -612 40102
rect -556 40046 -488 40102
rect -432 40046 -336 40102
rect -956 39978 -336 40046
rect -956 39922 -860 39978
rect -804 39922 -736 39978
rect -680 39922 -612 39978
rect -556 39922 -488 39978
rect -432 39922 -336 39978
rect -956 22350 -336 39922
rect 28 544740 84 544750
rect 28 25060 84 544684
rect 3164 523348 3220 523358
rect 2492 502516 2548 502526
rect 28 24994 84 25004
rect 140 474180 196 474190
rect -956 22294 -860 22350
rect -804 22294 -736 22350
rect -680 22294 -612 22350
rect -556 22294 -488 22350
rect -432 22294 -336 22350
rect -956 22226 -336 22294
rect -956 22170 -860 22226
rect -804 22170 -736 22226
rect -680 22170 -612 22226
rect -556 22170 -488 22226
rect -432 22170 -336 22226
rect -956 22102 -336 22170
rect -956 22046 -860 22102
rect -804 22046 -736 22102
rect -680 22046 -612 22102
rect -556 22046 -488 22102
rect -432 22046 -336 22102
rect -956 21978 -336 22046
rect -956 21922 -860 21978
rect -804 21922 -736 21978
rect -680 21922 -612 21978
rect -556 21922 -488 21978
rect -432 21922 -336 21978
rect -956 4350 -336 21922
rect 140 20580 196 474124
rect 140 20514 196 20524
rect 252 417732 308 417742
rect 252 16996 308 417676
rect 588 333172 644 333182
rect 588 314188 644 333116
rect 252 16930 308 16940
rect 364 314132 644 314188
rect 364 11620 420 314132
rect 2492 22372 2548 502460
rect 2492 22306 2548 22316
rect 2604 375508 2660 375518
rect 2604 14308 2660 375452
rect 2604 14242 2660 14252
rect 2716 347284 2772 347294
rect 2716 12516 2772 347228
rect 3052 80038 3108 80048
rect 3052 32228 3108 79982
rect 3164 54628 3220 523292
rect 3164 54562 3220 54572
rect 3052 32162 3108 32172
rect 3276 27748 3332 576062
rect 5418 562350 6038 579922
rect 5418 562294 5514 562350
rect 5570 562294 5638 562350
rect 5694 562294 5762 562350
rect 5818 562294 5886 562350
rect 5942 562294 6038 562350
rect 5418 562226 6038 562294
rect 5418 562170 5514 562226
rect 5570 562170 5638 562226
rect 5694 562170 5762 562226
rect 5818 562170 5886 562226
rect 5942 562170 6038 562226
rect 5418 562102 6038 562170
rect 5418 562046 5514 562102
rect 5570 562046 5638 562102
rect 5694 562046 5762 562102
rect 5818 562046 5886 562102
rect 5942 562046 6038 562102
rect 5418 561978 6038 562046
rect 5418 561922 5514 561978
rect 5570 561922 5638 561978
rect 5694 561922 5762 561978
rect 5818 561922 5886 561978
rect 5942 561922 6038 561978
rect 5418 544350 6038 561922
rect 5418 544294 5514 544350
rect 5570 544294 5638 544350
rect 5694 544294 5762 544350
rect 5818 544294 5886 544350
rect 5942 544294 6038 544350
rect 5418 544226 6038 544294
rect 5418 544170 5514 544226
rect 5570 544170 5638 544226
rect 5694 544170 5762 544226
rect 5818 544170 5886 544226
rect 5942 544170 6038 544226
rect 5418 544102 6038 544170
rect 5418 544046 5514 544102
rect 5570 544046 5638 544102
rect 5694 544046 5762 544102
rect 5818 544046 5886 544102
rect 5942 544046 6038 544102
rect 5418 543978 6038 544046
rect 5418 543922 5514 543978
rect 5570 543922 5638 543978
rect 5694 543922 5762 543978
rect 5818 543922 5886 543978
rect 5942 543922 6038 543978
rect 5418 526350 6038 543922
rect 5418 526294 5514 526350
rect 5570 526294 5638 526350
rect 5694 526294 5762 526350
rect 5818 526294 5886 526350
rect 5942 526294 6038 526350
rect 5418 526226 6038 526294
rect 5418 526170 5514 526226
rect 5570 526170 5638 526226
rect 5694 526170 5762 526226
rect 5818 526170 5886 526226
rect 5942 526170 6038 526226
rect 5418 526102 6038 526170
rect 5418 526046 5514 526102
rect 5570 526046 5638 526102
rect 5694 526046 5762 526102
rect 5818 526046 5886 526102
rect 5942 526046 6038 526102
rect 5418 525978 6038 526046
rect 5418 525922 5514 525978
rect 5570 525922 5638 525978
rect 5694 525922 5762 525978
rect 5818 525922 5886 525978
rect 5942 525922 6038 525978
rect 5418 508350 6038 525922
rect 5418 508294 5514 508350
rect 5570 508294 5638 508350
rect 5694 508294 5762 508350
rect 5818 508294 5886 508350
rect 5942 508294 6038 508350
rect 5418 508226 6038 508294
rect 5418 508170 5514 508226
rect 5570 508170 5638 508226
rect 5694 508170 5762 508226
rect 5818 508170 5886 508226
rect 5942 508170 6038 508226
rect 5418 508102 6038 508170
rect 5418 508046 5514 508102
rect 5570 508046 5638 508102
rect 5694 508046 5762 508102
rect 5818 508046 5886 508102
rect 5942 508046 6038 508102
rect 5418 507978 6038 508046
rect 5418 507922 5514 507978
rect 5570 507922 5638 507978
rect 5694 507922 5762 507978
rect 5818 507922 5886 507978
rect 5942 507922 6038 507978
rect 5418 490350 6038 507922
rect 5418 490294 5514 490350
rect 5570 490294 5638 490350
rect 5694 490294 5762 490350
rect 5818 490294 5886 490350
rect 5942 490294 6038 490350
rect 5418 490226 6038 490294
rect 5418 490170 5514 490226
rect 5570 490170 5638 490226
rect 5694 490170 5762 490226
rect 5818 490170 5886 490226
rect 5942 490170 6038 490226
rect 5418 490102 6038 490170
rect 5418 490046 5514 490102
rect 5570 490046 5638 490102
rect 5694 490046 5762 490102
rect 5818 490046 5886 490102
rect 5942 490046 6038 490102
rect 5418 489978 6038 490046
rect 5418 489922 5514 489978
rect 5570 489922 5638 489978
rect 5694 489922 5762 489978
rect 5818 489922 5886 489978
rect 5942 489922 6038 489978
rect 5418 472350 6038 489922
rect 9138 598172 9758 598268
rect 9138 598116 9234 598172
rect 9290 598116 9358 598172
rect 9414 598116 9482 598172
rect 9538 598116 9606 598172
rect 9662 598116 9758 598172
rect 9138 598048 9758 598116
rect 9138 597992 9234 598048
rect 9290 597992 9358 598048
rect 9414 597992 9482 598048
rect 9538 597992 9606 598048
rect 9662 597992 9758 598048
rect 9138 597924 9758 597992
rect 9138 597868 9234 597924
rect 9290 597868 9358 597924
rect 9414 597868 9482 597924
rect 9538 597868 9606 597924
rect 9662 597868 9758 597924
rect 9138 597800 9758 597868
rect 9138 597744 9234 597800
rect 9290 597744 9358 597800
rect 9414 597744 9482 597800
rect 9538 597744 9606 597800
rect 9662 597744 9758 597800
rect 9138 586350 9758 597744
rect 36138 597212 36758 598268
rect 36138 597156 36234 597212
rect 36290 597156 36358 597212
rect 36414 597156 36482 597212
rect 36538 597156 36606 597212
rect 36662 597156 36758 597212
rect 36138 597088 36758 597156
rect 36138 597032 36234 597088
rect 36290 597032 36358 597088
rect 36414 597032 36482 597088
rect 36538 597032 36606 597088
rect 36662 597032 36758 597088
rect 36138 596964 36758 597032
rect 36138 596908 36234 596964
rect 36290 596908 36358 596964
rect 36414 596908 36482 596964
rect 36538 596908 36606 596964
rect 36662 596908 36758 596964
rect 36138 596840 36758 596908
rect 36138 596784 36234 596840
rect 36290 596784 36358 596840
rect 36414 596784 36482 596840
rect 36538 596784 36606 596840
rect 36662 596784 36758 596840
rect 27692 590660 27748 590670
rect 9138 586294 9234 586350
rect 9290 586294 9358 586350
rect 9414 586294 9482 586350
rect 9538 586294 9606 586350
rect 9662 586294 9758 586350
rect 9138 586226 9758 586294
rect 9138 586170 9234 586226
rect 9290 586170 9358 586226
rect 9414 586170 9482 586226
rect 9538 586170 9606 586226
rect 9662 586170 9758 586226
rect 9138 586102 9758 586170
rect 9138 586046 9234 586102
rect 9290 586046 9358 586102
rect 9414 586046 9482 586102
rect 9538 586046 9606 586102
rect 9662 586046 9758 586102
rect 9138 585978 9758 586046
rect 9138 585922 9234 585978
rect 9290 585922 9358 585978
rect 9414 585922 9482 585978
rect 9538 585922 9606 585978
rect 9662 585922 9758 585978
rect 9138 568350 9758 585922
rect 26012 588644 26068 588654
rect 22652 582148 22708 582158
rect 19292 578788 19348 578798
rect 17612 575428 17668 575438
rect 9138 568294 9234 568350
rect 9290 568294 9358 568350
rect 9414 568294 9482 568350
rect 9538 568294 9606 568350
rect 9662 568294 9758 568350
rect 9138 568226 9758 568294
rect 9138 568170 9234 568226
rect 9290 568170 9358 568226
rect 9414 568170 9482 568226
rect 9538 568170 9606 568226
rect 9662 568170 9758 568226
rect 9138 568102 9758 568170
rect 9138 568046 9234 568102
rect 9290 568046 9358 568102
rect 9414 568046 9482 568102
rect 9538 568046 9606 568102
rect 9662 568046 9758 568102
rect 9138 567978 9758 568046
rect 9138 567922 9234 567978
rect 9290 567922 9358 567978
rect 9414 567922 9482 567978
rect 9538 567922 9606 567978
rect 9662 567922 9758 567978
rect 9138 550350 9758 567922
rect 12012 573076 12068 573086
rect 9138 550294 9234 550350
rect 9290 550294 9358 550350
rect 9414 550294 9482 550350
rect 9538 550294 9606 550350
rect 9662 550294 9758 550350
rect 9138 550226 9758 550294
rect 9138 550170 9234 550226
rect 9290 550170 9358 550226
rect 9414 550170 9482 550226
rect 9538 550170 9606 550226
rect 9662 550170 9758 550226
rect 9138 550102 9758 550170
rect 9138 550046 9234 550102
rect 9290 550046 9358 550102
rect 9414 550046 9482 550102
rect 9538 550046 9606 550102
rect 9662 550046 9758 550102
rect 9138 549978 9758 550046
rect 9138 549922 9234 549978
rect 9290 549922 9358 549978
rect 9414 549922 9482 549978
rect 9538 549922 9606 549978
rect 9662 549922 9758 549978
rect 9138 532350 9758 549922
rect 9138 532294 9234 532350
rect 9290 532294 9358 532350
rect 9414 532294 9482 532350
rect 9538 532294 9606 532350
rect 9662 532294 9758 532350
rect 9138 532226 9758 532294
rect 9138 532170 9234 532226
rect 9290 532170 9358 532226
rect 9414 532170 9482 532226
rect 9538 532170 9606 532226
rect 9662 532170 9758 532226
rect 9138 532102 9758 532170
rect 9138 532046 9234 532102
rect 9290 532046 9358 532102
rect 9414 532046 9482 532102
rect 9538 532046 9606 532102
rect 9662 532046 9758 532102
rect 9138 531978 9758 532046
rect 9138 531922 9234 531978
rect 9290 531922 9358 531978
rect 9414 531922 9482 531978
rect 9538 531922 9606 531978
rect 9662 531922 9758 531978
rect 9138 514350 9758 531922
rect 9138 514294 9234 514350
rect 9290 514294 9358 514350
rect 9414 514294 9482 514350
rect 9538 514294 9606 514350
rect 9662 514294 9758 514350
rect 9138 514226 9758 514294
rect 9138 514170 9234 514226
rect 9290 514170 9358 514226
rect 9414 514170 9482 514226
rect 9538 514170 9606 514226
rect 9662 514170 9758 514226
rect 9138 514102 9758 514170
rect 9138 514046 9234 514102
rect 9290 514046 9358 514102
rect 9414 514046 9482 514102
rect 9538 514046 9606 514102
rect 9662 514046 9758 514102
rect 9138 513978 9758 514046
rect 9138 513922 9234 513978
rect 9290 513922 9358 513978
rect 9414 513922 9482 513978
rect 9538 513922 9606 513978
rect 9662 513922 9758 513978
rect 9138 496350 9758 513922
rect 9138 496294 9234 496350
rect 9290 496294 9358 496350
rect 9414 496294 9482 496350
rect 9538 496294 9606 496350
rect 9662 496294 9758 496350
rect 9138 496226 9758 496294
rect 9138 496170 9234 496226
rect 9290 496170 9358 496226
rect 9414 496170 9482 496226
rect 9538 496170 9606 496226
rect 9662 496170 9758 496226
rect 9138 496102 9758 496170
rect 9138 496046 9234 496102
rect 9290 496046 9358 496102
rect 9414 496046 9482 496102
rect 9538 496046 9606 496102
rect 9662 496046 9758 496102
rect 9138 495978 9758 496046
rect 9138 495922 9234 495978
rect 9290 495922 9358 495978
rect 9414 495922 9482 495978
rect 9538 495922 9606 495978
rect 9662 495922 9758 495978
rect 5418 472294 5514 472350
rect 5570 472294 5638 472350
rect 5694 472294 5762 472350
rect 5818 472294 5886 472350
rect 5942 472294 6038 472350
rect 5418 472226 6038 472294
rect 5418 472170 5514 472226
rect 5570 472170 5638 472226
rect 5694 472170 5762 472226
rect 5818 472170 5886 472226
rect 5942 472170 6038 472226
rect 5418 472102 6038 472170
rect 5418 472046 5514 472102
rect 5570 472046 5638 472102
rect 5694 472046 5762 472102
rect 5818 472046 5886 472102
rect 5942 472046 6038 472102
rect 5418 471978 6038 472046
rect 5418 471922 5514 471978
rect 5570 471922 5638 471978
rect 5694 471922 5762 471978
rect 5818 471922 5886 471978
rect 5942 471922 6038 471978
rect 5418 454350 6038 471922
rect 8316 482916 8372 482926
rect 5418 454294 5514 454350
rect 5570 454294 5638 454350
rect 5694 454294 5762 454350
rect 5818 454294 5886 454350
rect 5942 454294 6038 454350
rect 5418 454226 6038 454294
rect 5418 454170 5514 454226
rect 5570 454170 5638 454226
rect 5694 454170 5762 454226
rect 5818 454170 5886 454226
rect 5942 454170 6038 454226
rect 5418 454102 6038 454170
rect 5418 454046 5514 454102
rect 5570 454046 5638 454102
rect 5694 454046 5762 454102
rect 5818 454046 5886 454102
rect 5942 454046 6038 454102
rect 5418 453978 6038 454046
rect 5418 453922 5514 453978
rect 5570 453922 5638 453978
rect 5694 453922 5762 453978
rect 5818 453922 5886 453978
rect 5942 453922 6038 453978
rect 4620 446068 4676 446078
rect 3276 27682 3332 27692
rect 4172 431956 4228 431966
rect 4172 17892 4228 431900
rect 4172 17826 4228 17836
rect 4284 389620 4340 389630
rect 4284 15204 4340 389564
rect 4284 15138 4340 15148
rect 4396 304948 4452 304958
rect 2716 12450 2772 12460
rect 364 11554 420 11564
rect 4396 9828 4452 304892
rect 4620 304164 4676 446012
rect 5418 436350 6038 453922
rect 5418 436294 5514 436350
rect 5570 436294 5638 436350
rect 5694 436294 5762 436350
rect 5818 436294 5886 436350
rect 5942 436294 6038 436350
rect 5418 436226 6038 436294
rect 5418 436170 5514 436226
rect 5570 436170 5638 436226
rect 5694 436170 5762 436226
rect 5818 436170 5886 436226
rect 5942 436170 6038 436226
rect 5418 436102 6038 436170
rect 5418 436046 5514 436102
rect 5570 436046 5638 436102
rect 5694 436046 5762 436102
rect 5818 436046 5886 436102
rect 5942 436046 6038 436102
rect 5418 435978 6038 436046
rect 5418 435922 5514 435978
rect 5570 435922 5638 435978
rect 5694 435922 5762 435978
rect 5818 435922 5886 435978
rect 5942 435922 6038 435978
rect 5418 418350 6038 435922
rect 5418 418294 5514 418350
rect 5570 418294 5638 418350
rect 5694 418294 5762 418350
rect 5818 418294 5886 418350
rect 5942 418294 6038 418350
rect 5418 418226 6038 418294
rect 5418 418170 5514 418226
rect 5570 418170 5638 418226
rect 5694 418170 5762 418226
rect 5818 418170 5886 418226
rect 5942 418170 6038 418226
rect 5418 418102 6038 418170
rect 5418 418046 5514 418102
rect 5570 418046 5638 418102
rect 5694 418046 5762 418102
rect 5818 418046 5886 418102
rect 5942 418046 6038 418102
rect 5418 417978 6038 418046
rect 5418 417922 5514 417978
rect 5570 417922 5638 417978
rect 5694 417922 5762 417978
rect 5818 417922 5886 417978
rect 5942 417922 6038 417978
rect 5418 400350 6038 417922
rect 5418 400294 5514 400350
rect 5570 400294 5638 400350
rect 5694 400294 5762 400350
rect 5818 400294 5886 400350
rect 5942 400294 6038 400350
rect 5418 400226 6038 400294
rect 5418 400170 5514 400226
rect 5570 400170 5638 400226
rect 5694 400170 5762 400226
rect 5818 400170 5886 400226
rect 5942 400170 6038 400226
rect 5418 400102 6038 400170
rect 5418 400046 5514 400102
rect 5570 400046 5638 400102
rect 5694 400046 5762 400102
rect 5818 400046 5886 400102
rect 5942 400046 6038 400102
rect 5418 399978 6038 400046
rect 5418 399922 5514 399978
rect 5570 399922 5638 399978
rect 5694 399922 5762 399978
rect 5818 399922 5886 399978
rect 5942 399922 6038 399978
rect 5418 382350 6038 399922
rect 5418 382294 5514 382350
rect 5570 382294 5638 382350
rect 5694 382294 5762 382350
rect 5818 382294 5886 382350
rect 5942 382294 6038 382350
rect 5418 382226 6038 382294
rect 5418 382170 5514 382226
rect 5570 382170 5638 382226
rect 5694 382170 5762 382226
rect 5818 382170 5886 382226
rect 5942 382170 6038 382226
rect 5418 382102 6038 382170
rect 5418 382046 5514 382102
rect 5570 382046 5638 382102
rect 5694 382046 5762 382102
rect 5818 382046 5886 382102
rect 5942 382046 6038 382102
rect 5418 381978 6038 382046
rect 5418 381922 5514 381978
rect 5570 381922 5638 381978
rect 5694 381922 5762 381978
rect 5818 381922 5886 381978
rect 5942 381922 6038 381978
rect 5418 364350 6038 381922
rect 5418 364294 5514 364350
rect 5570 364294 5638 364350
rect 5694 364294 5762 364350
rect 5818 364294 5886 364350
rect 5942 364294 6038 364350
rect 5418 364226 6038 364294
rect 5418 364170 5514 364226
rect 5570 364170 5638 364226
rect 5694 364170 5762 364226
rect 5818 364170 5886 364226
rect 5942 364170 6038 364226
rect 5418 364102 6038 364170
rect 5418 364046 5514 364102
rect 5570 364046 5638 364102
rect 5694 364046 5762 364102
rect 5818 364046 5886 364102
rect 5942 364046 6038 364102
rect 5418 363978 6038 364046
rect 5418 363922 5514 363978
rect 5570 363922 5638 363978
rect 5694 363922 5762 363978
rect 5818 363922 5886 363978
rect 5942 363922 6038 363978
rect 4620 304098 4676 304108
rect 4732 361396 4788 361406
rect 4396 9762 4452 9772
rect 4508 276724 4564 276734
rect 4508 8036 4564 276668
rect 4732 275604 4788 361340
rect 4732 275538 4788 275548
rect 5418 346350 6038 363922
rect 5418 346294 5514 346350
rect 5570 346294 5638 346350
rect 5694 346294 5762 346350
rect 5818 346294 5886 346350
rect 5942 346294 6038 346350
rect 5418 346226 6038 346294
rect 5418 346170 5514 346226
rect 5570 346170 5638 346226
rect 5694 346170 5762 346226
rect 5818 346170 5886 346226
rect 5942 346170 6038 346226
rect 5418 346102 6038 346170
rect 5418 346046 5514 346102
rect 5570 346046 5638 346102
rect 5694 346046 5762 346102
rect 5818 346046 5886 346102
rect 5942 346046 6038 346102
rect 5418 345978 6038 346046
rect 5418 345922 5514 345978
rect 5570 345922 5638 345978
rect 5694 345922 5762 345978
rect 5818 345922 5886 345978
rect 5942 345922 6038 345978
rect 5418 328350 6038 345922
rect 5418 328294 5514 328350
rect 5570 328294 5638 328350
rect 5694 328294 5762 328350
rect 5818 328294 5886 328350
rect 5942 328294 6038 328350
rect 5418 328226 6038 328294
rect 5418 328170 5514 328226
rect 5570 328170 5638 328226
rect 5694 328170 5762 328226
rect 5818 328170 5886 328226
rect 5942 328170 6038 328226
rect 5418 328102 6038 328170
rect 5418 328046 5514 328102
rect 5570 328046 5638 328102
rect 5694 328046 5762 328102
rect 5818 328046 5886 328102
rect 5942 328046 6038 328102
rect 5418 327978 6038 328046
rect 5418 327922 5514 327978
rect 5570 327922 5638 327978
rect 5694 327922 5762 327978
rect 5818 327922 5886 327978
rect 5942 327922 6038 327978
rect 5418 310350 6038 327922
rect 5418 310294 5514 310350
rect 5570 310294 5638 310350
rect 5694 310294 5762 310350
rect 5818 310294 5886 310350
rect 5942 310294 6038 310350
rect 5418 310226 6038 310294
rect 5418 310170 5514 310226
rect 5570 310170 5638 310226
rect 5694 310170 5762 310226
rect 5818 310170 5886 310226
rect 5942 310170 6038 310226
rect 5418 310102 6038 310170
rect 5418 310046 5514 310102
rect 5570 310046 5638 310102
rect 5694 310046 5762 310102
rect 5818 310046 5886 310102
rect 5942 310046 6038 310102
rect 5418 309978 6038 310046
rect 5418 309922 5514 309978
rect 5570 309922 5638 309978
rect 5694 309922 5762 309978
rect 5818 309922 5886 309978
rect 5942 309922 6038 309978
rect 5418 292350 6038 309922
rect 5418 292294 5514 292350
rect 5570 292294 5638 292350
rect 5694 292294 5762 292350
rect 5818 292294 5886 292350
rect 5942 292294 6038 292350
rect 5418 292226 6038 292294
rect 5418 292170 5514 292226
rect 5570 292170 5638 292226
rect 5694 292170 5762 292226
rect 5818 292170 5886 292226
rect 5942 292170 6038 292226
rect 5418 292102 6038 292170
rect 5418 292046 5514 292102
rect 5570 292046 5638 292102
rect 5694 292046 5762 292102
rect 5818 292046 5886 292102
rect 5942 292046 6038 292102
rect 5418 291978 6038 292046
rect 5418 291922 5514 291978
rect 5570 291922 5638 291978
rect 5694 291922 5762 291978
rect 5818 291922 5886 291978
rect 5942 291922 6038 291978
rect 5418 274350 6038 291922
rect 7532 460180 7588 460190
rect 5418 274294 5514 274350
rect 5570 274294 5638 274350
rect 5694 274294 5762 274350
rect 5818 274294 5886 274350
rect 5942 274294 6038 274350
rect 5418 274226 6038 274294
rect 5418 274170 5514 274226
rect 5570 274170 5638 274226
rect 5694 274170 5762 274226
rect 5818 274170 5886 274226
rect 5942 274170 6038 274226
rect 5418 274102 6038 274170
rect 5418 274046 5514 274102
rect 5570 274046 5638 274102
rect 5694 274046 5762 274102
rect 5818 274046 5886 274102
rect 5942 274046 6038 274102
rect 5418 273978 6038 274046
rect 5418 273922 5514 273978
rect 5570 273922 5638 273978
rect 5694 273922 5762 273978
rect 5818 273922 5886 273978
rect 5942 273922 6038 273978
rect 4620 262612 4676 262622
rect 4620 33572 4676 262556
rect 4620 33506 4676 33516
rect 5418 256350 6038 273922
rect 5418 256294 5514 256350
rect 5570 256294 5638 256350
rect 5694 256294 5762 256350
rect 5818 256294 5886 256350
rect 5942 256294 6038 256350
rect 5418 256226 6038 256294
rect 5418 256170 5514 256226
rect 5570 256170 5638 256226
rect 5694 256170 5762 256226
rect 5818 256170 5886 256226
rect 5942 256170 6038 256226
rect 5418 256102 6038 256170
rect 5418 256046 5514 256102
rect 5570 256046 5638 256102
rect 5694 256046 5762 256102
rect 5818 256046 5886 256102
rect 5942 256046 6038 256102
rect 5418 255978 6038 256046
rect 5418 255922 5514 255978
rect 5570 255922 5638 255978
rect 5694 255922 5762 255978
rect 5818 255922 5886 255978
rect 5942 255922 6038 255978
rect 5418 238350 6038 255922
rect 5418 238294 5514 238350
rect 5570 238294 5638 238350
rect 5694 238294 5762 238350
rect 5818 238294 5886 238350
rect 5942 238294 6038 238350
rect 5418 238226 6038 238294
rect 5418 238170 5514 238226
rect 5570 238170 5638 238226
rect 5694 238170 5762 238226
rect 5818 238170 5886 238226
rect 5942 238170 6038 238226
rect 5418 238102 6038 238170
rect 5418 238046 5514 238102
rect 5570 238046 5638 238102
rect 5694 238046 5762 238102
rect 5818 238046 5886 238102
rect 5942 238046 6038 238102
rect 5418 237978 6038 238046
rect 5418 237922 5514 237978
rect 5570 237922 5638 237978
rect 5694 237922 5762 237978
rect 5818 237922 5886 237978
rect 5942 237922 6038 237978
rect 5418 220350 6038 237922
rect 5418 220294 5514 220350
rect 5570 220294 5638 220350
rect 5694 220294 5762 220350
rect 5818 220294 5886 220350
rect 5942 220294 6038 220350
rect 5418 220226 6038 220294
rect 5418 220170 5514 220226
rect 5570 220170 5638 220226
rect 5694 220170 5762 220226
rect 5818 220170 5886 220226
rect 5942 220170 6038 220226
rect 5418 220102 6038 220170
rect 5418 220046 5514 220102
rect 5570 220046 5638 220102
rect 5694 220046 5762 220102
rect 5818 220046 5886 220102
rect 5942 220046 6038 220102
rect 5418 219978 6038 220046
rect 5418 219922 5514 219978
rect 5570 219922 5638 219978
rect 5694 219922 5762 219978
rect 5818 219922 5886 219978
rect 5942 219922 6038 219978
rect 5418 202350 6038 219922
rect 5418 202294 5514 202350
rect 5570 202294 5638 202350
rect 5694 202294 5762 202350
rect 5818 202294 5886 202350
rect 5942 202294 6038 202350
rect 5418 202226 6038 202294
rect 5418 202170 5514 202226
rect 5570 202170 5638 202226
rect 5694 202170 5762 202226
rect 5818 202170 5886 202226
rect 5942 202170 6038 202226
rect 5418 202102 6038 202170
rect 5418 202046 5514 202102
rect 5570 202046 5638 202102
rect 5694 202046 5762 202102
rect 5818 202046 5886 202102
rect 5942 202046 6038 202102
rect 5418 201978 6038 202046
rect 5418 201922 5514 201978
rect 5570 201922 5638 201978
rect 5694 201922 5762 201978
rect 5818 201922 5886 201978
rect 5942 201922 6038 201978
rect 5418 184350 6038 201922
rect 5418 184294 5514 184350
rect 5570 184294 5638 184350
rect 5694 184294 5762 184350
rect 5818 184294 5886 184350
rect 5942 184294 6038 184350
rect 5418 184226 6038 184294
rect 5418 184170 5514 184226
rect 5570 184170 5638 184226
rect 5694 184170 5762 184226
rect 5818 184170 5886 184226
rect 5942 184170 6038 184226
rect 5418 184102 6038 184170
rect 5418 184046 5514 184102
rect 5570 184046 5638 184102
rect 5694 184046 5762 184102
rect 5818 184046 5886 184102
rect 5942 184046 6038 184102
rect 5418 183978 6038 184046
rect 5418 183922 5514 183978
rect 5570 183922 5638 183978
rect 5694 183922 5762 183978
rect 5818 183922 5886 183978
rect 5942 183922 6038 183978
rect 5418 166350 6038 183922
rect 5418 166294 5514 166350
rect 5570 166294 5638 166350
rect 5694 166294 5762 166350
rect 5818 166294 5886 166350
rect 5942 166294 6038 166350
rect 5418 166226 6038 166294
rect 5418 166170 5514 166226
rect 5570 166170 5638 166226
rect 5694 166170 5762 166226
rect 5818 166170 5886 166226
rect 5942 166170 6038 166226
rect 5418 166102 6038 166170
rect 5418 166046 5514 166102
rect 5570 166046 5638 166102
rect 5694 166046 5762 166102
rect 5818 166046 5886 166102
rect 5942 166046 6038 166102
rect 5418 165978 6038 166046
rect 5418 165922 5514 165978
rect 5570 165922 5638 165978
rect 5694 165922 5762 165978
rect 5818 165922 5886 165978
rect 5942 165922 6038 165978
rect 5418 148350 6038 165922
rect 5418 148294 5514 148350
rect 5570 148294 5638 148350
rect 5694 148294 5762 148350
rect 5818 148294 5886 148350
rect 5942 148294 6038 148350
rect 5418 148226 6038 148294
rect 5418 148170 5514 148226
rect 5570 148170 5638 148226
rect 5694 148170 5762 148226
rect 5818 148170 5886 148226
rect 5942 148170 6038 148226
rect 5418 148102 6038 148170
rect 5418 148046 5514 148102
rect 5570 148046 5638 148102
rect 5694 148046 5762 148102
rect 5818 148046 5886 148102
rect 5942 148046 6038 148102
rect 5418 147978 6038 148046
rect 5418 147922 5514 147978
rect 5570 147922 5638 147978
rect 5694 147922 5762 147978
rect 5818 147922 5886 147978
rect 5942 147922 6038 147978
rect 5418 130350 6038 147922
rect 5418 130294 5514 130350
rect 5570 130294 5638 130350
rect 5694 130294 5762 130350
rect 5818 130294 5886 130350
rect 5942 130294 6038 130350
rect 5418 130226 6038 130294
rect 5418 130170 5514 130226
rect 5570 130170 5638 130226
rect 5694 130170 5762 130226
rect 5818 130170 5886 130226
rect 5942 130170 6038 130226
rect 5418 130102 6038 130170
rect 5418 130046 5514 130102
rect 5570 130046 5638 130102
rect 5694 130046 5762 130102
rect 5818 130046 5886 130102
rect 5942 130046 6038 130102
rect 5418 129978 6038 130046
rect 5418 129922 5514 129978
rect 5570 129922 5638 129978
rect 5694 129922 5762 129978
rect 5818 129922 5886 129978
rect 5942 129922 6038 129978
rect 5418 112350 6038 129922
rect 5418 112294 5514 112350
rect 5570 112294 5638 112350
rect 5694 112294 5762 112350
rect 5818 112294 5886 112350
rect 5942 112294 6038 112350
rect 5418 112226 6038 112294
rect 5418 112170 5514 112226
rect 5570 112170 5638 112226
rect 5694 112170 5762 112226
rect 5818 112170 5886 112226
rect 5942 112170 6038 112226
rect 5418 112102 6038 112170
rect 5418 112046 5514 112102
rect 5570 112046 5638 112102
rect 5694 112046 5762 112102
rect 5818 112046 5886 112102
rect 5942 112046 6038 112102
rect 5418 111978 6038 112046
rect 5418 111922 5514 111978
rect 5570 111922 5638 111978
rect 5694 111922 5762 111978
rect 5818 111922 5886 111978
rect 5942 111922 6038 111978
rect 5418 94350 6038 111922
rect 5418 94294 5514 94350
rect 5570 94294 5638 94350
rect 5694 94294 5762 94350
rect 5818 94294 5886 94350
rect 5942 94294 6038 94350
rect 5418 94226 6038 94294
rect 5418 94170 5514 94226
rect 5570 94170 5638 94226
rect 5694 94170 5762 94226
rect 5818 94170 5886 94226
rect 5942 94170 6038 94226
rect 5418 94102 6038 94170
rect 5418 94046 5514 94102
rect 5570 94046 5638 94102
rect 5694 94046 5762 94102
rect 5818 94046 5886 94102
rect 5942 94046 6038 94102
rect 5418 93978 6038 94046
rect 5418 93922 5514 93978
rect 5570 93922 5638 93978
rect 5694 93922 5762 93978
rect 5818 93922 5886 93978
rect 5942 93922 6038 93978
rect 5418 76350 6038 93922
rect 5418 76294 5514 76350
rect 5570 76294 5638 76350
rect 5694 76294 5762 76350
rect 5818 76294 5886 76350
rect 5942 76294 6038 76350
rect 5418 76226 6038 76294
rect 5418 76170 5514 76226
rect 5570 76170 5638 76226
rect 5694 76170 5762 76226
rect 5818 76170 5886 76226
rect 5942 76170 6038 76226
rect 5418 76102 6038 76170
rect 5418 76046 5514 76102
rect 5570 76046 5638 76102
rect 5694 76046 5762 76102
rect 5818 76046 5886 76102
rect 5942 76046 6038 76102
rect 5418 75978 6038 76046
rect 5418 75922 5514 75978
rect 5570 75922 5638 75978
rect 5694 75922 5762 75978
rect 5818 75922 5886 75978
rect 5942 75922 6038 75978
rect 5418 58350 6038 75922
rect 5418 58294 5514 58350
rect 5570 58294 5638 58350
rect 5694 58294 5762 58350
rect 5818 58294 5886 58350
rect 5942 58294 6038 58350
rect 5418 58226 6038 58294
rect 5418 58170 5514 58226
rect 5570 58170 5638 58226
rect 5694 58170 5762 58226
rect 5818 58170 5886 58226
rect 5942 58170 6038 58226
rect 5418 58102 6038 58170
rect 5418 58046 5514 58102
rect 5570 58046 5638 58102
rect 5694 58046 5762 58102
rect 5818 58046 5886 58102
rect 5942 58046 6038 58102
rect 5418 57978 6038 58046
rect 5418 57922 5514 57978
rect 5570 57922 5638 57978
rect 5694 57922 5762 57978
rect 5818 57922 5886 57978
rect 5942 57922 6038 57978
rect 5418 40350 6038 57922
rect 5418 40294 5514 40350
rect 5570 40294 5638 40350
rect 5694 40294 5762 40350
rect 5818 40294 5886 40350
rect 5942 40294 6038 40350
rect 5418 40226 6038 40294
rect 5418 40170 5514 40226
rect 5570 40170 5638 40226
rect 5694 40170 5762 40226
rect 5818 40170 5886 40226
rect 5942 40170 6038 40226
rect 5418 40102 6038 40170
rect 5418 40046 5514 40102
rect 5570 40046 5638 40102
rect 5694 40046 5762 40102
rect 5818 40046 5886 40102
rect 5942 40046 6038 40102
rect 5418 39978 6038 40046
rect 5418 39922 5514 39978
rect 5570 39922 5638 39978
rect 5694 39922 5762 39978
rect 5818 39922 5886 39978
rect 5942 39922 6038 39978
rect 4508 7970 4564 7980
rect 5418 22350 6038 39922
rect 5418 22294 5514 22350
rect 5570 22294 5638 22350
rect 5694 22294 5762 22350
rect 5818 22294 5886 22350
rect 5942 22294 6038 22350
rect 5418 22226 6038 22294
rect 5418 22170 5514 22226
rect 5570 22170 5638 22226
rect 5694 22170 5762 22226
rect 5818 22170 5886 22226
rect 5942 22170 6038 22226
rect 5418 22102 6038 22170
rect 5418 22046 5514 22102
rect 5570 22046 5638 22102
rect 5694 22046 5762 22102
rect 5818 22046 5886 22102
rect 5942 22046 6038 22102
rect 5418 21978 6038 22046
rect 5418 21922 5514 21978
rect 5570 21922 5638 21978
rect 5694 21922 5762 21978
rect 5818 21922 5886 21978
rect 5942 21922 6038 21978
rect -956 4294 -860 4350
rect -804 4294 -736 4350
rect -680 4294 -612 4350
rect -556 4294 -488 4350
rect -432 4294 -336 4350
rect -956 4226 -336 4294
rect -956 4170 -860 4226
rect -804 4170 -736 4226
rect -680 4170 -612 4226
rect -556 4170 -488 4226
rect -432 4170 -336 4226
rect -956 4102 -336 4170
rect -956 4046 -860 4102
rect -804 4046 -736 4102
rect -680 4046 -612 4102
rect -556 4046 -488 4102
rect -432 4046 -336 4102
rect -956 3978 -336 4046
rect -956 3922 -860 3978
rect -804 3922 -736 3978
rect -680 3922 -612 3978
rect -556 3922 -488 3978
rect -432 3922 -336 3978
rect -956 -160 -336 3922
rect -956 -216 -860 -160
rect -804 -216 -736 -160
rect -680 -216 -612 -160
rect -556 -216 -488 -160
rect -432 -216 -336 -160
rect -956 -284 -336 -216
rect -956 -340 -860 -284
rect -804 -340 -736 -284
rect -680 -340 -612 -284
rect -556 -340 -488 -284
rect -432 -340 -336 -284
rect -956 -408 -336 -340
rect -956 -464 -860 -408
rect -804 -464 -736 -408
rect -680 -464 -612 -408
rect -556 -464 -488 -408
rect -432 -464 -336 -408
rect -956 -532 -336 -464
rect -956 -588 -860 -532
rect -804 -588 -736 -532
rect -680 -588 -612 -532
rect -556 -588 -488 -532
rect -432 -588 -336 -532
rect -956 -684 -336 -588
rect 5418 4350 6038 21922
rect 6188 275604 6244 275614
rect 6188 13412 6244 275548
rect 6524 79858 6580 79868
rect 6524 42084 6580 79802
rect 6524 42018 6580 42028
rect 6636 78238 6692 78248
rect 6636 40292 6692 78182
rect 6636 40226 6692 40236
rect 7532 19684 7588 460124
rect 8204 403620 8260 403630
rect 7532 19618 7588 19628
rect 7644 290836 7700 290846
rect 6188 13346 6244 13356
rect 7644 8932 7700 290780
rect 8092 78418 8148 78428
rect 7980 74998 8036 75008
rect 7980 34916 8036 74942
rect 7980 34850 8036 34860
rect 7644 8866 7700 8876
rect 7756 33572 7812 33582
rect 7756 7140 7812 33516
rect 8092 33124 8148 78362
rect 8204 65380 8260 403564
rect 8204 65314 8260 65324
rect 8316 60004 8372 482860
rect 9138 478350 9758 495922
rect 9138 478294 9234 478350
rect 9290 478294 9358 478350
rect 9414 478294 9482 478350
rect 9538 478294 9606 478350
rect 9662 478294 9758 478350
rect 9138 478226 9758 478294
rect 9138 478170 9234 478226
rect 9290 478170 9358 478226
rect 9414 478170 9482 478226
rect 9538 478170 9606 478226
rect 9662 478170 9758 478226
rect 9138 478102 9758 478170
rect 9138 478046 9234 478102
rect 9290 478046 9358 478102
rect 9414 478046 9482 478102
rect 9538 478046 9606 478102
rect 9662 478046 9758 478102
rect 9138 477978 9758 478046
rect 9138 477922 9234 477978
rect 9290 477922 9358 477978
rect 9414 477922 9482 477978
rect 9538 477922 9606 477978
rect 9662 477922 9758 477978
rect 9138 460350 9758 477922
rect 9138 460294 9234 460350
rect 9290 460294 9358 460350
rect 9414 460294 9482 460350
rect 9538 460294 9606 460350
rect 9662 460294 9758 460350
rect 9138 460226 9758 460294
rect 9138 460170 9234 460226
rect 9290 460170 9358 460226
rect 9414 460170 9482 460226
rect 9538 460170 9606 460226
rect 9662 460170 9758 460226
rect 9138 460102 9758 460170
rect 9138 460046 9234 460102
rect 9290 460046 9358 460102
rect 9414 460046 9482 460102
rect 9538 460046 9606 460102
rect 9662 460046 9758 460102
rect 9138 459978 9758 460046
rect 9138 459922 9234 459978
rect 9290 459922 9358 459978
rect 9414 459922 9482 459978
rect 9538 459922 9606 459978
rect 9662 459922 9758 459978
rect 9138 442350 9758 459922
rect 9138 442294 9234 442350
rect 9290 442294 9358 442350
rect 9414 442294 9482 442350
rect 9538 442294 9606 442350
rect 9662 442294 9758 442350
rect 9138 442226 9758 442294
rect 9138 442170 9234 442226
rect 9290 442170 9358 442226
rect 9414 442170 9482 442226
rect 9538 442170 9606 442226
rect 9662 442170 9758 442226
rect 9138 442102 9758 442170
rect 9138 442046 9234 442102
rect 9290 442046 9358 442102
rect 9414 442046 9482 442102
rect 9538 442046 9606 442102
rect 9662 442046 9758 442102
rect 9138 441978 9758 442046
rect 9138 441922 9234 441978
rect 9290 441922 9358 441978
rect 9414 441922 9482 441978
rect 9538 441922 9606 441978
rect 9662 441922 9758 441978
rect 9138 424350 9758 441922
rect 9138 424294 9234 424350
rect 9290 424294 9358 424350
rect 9414 424294 9482 424350
rect 9538 424294 9606 424350
rect 9662 424294 9758 424350
rect 9138 424226 9758 424294
rect 9138 424170 9234 424226
rect 9290 424170 9358 424226
rect 9414 424170 9482 424226
rect 9538 424170 9606 424226
rect 9662 424170 9758 424226
rect 9138 424102 9758 424170
rect 9138 424046 9234 424102
rect 9290 424046 9358 424102
rect 9414 424046 9482 424102
rect 9538 424046 9606 424102
rect 9662 424046 9758 424102
rect 9138 423978 9758 424046
rect 9138 423922 9234 423978
rect 9290 423922 9358 423978
rect 9414 423922 9482 423978
rect 9538 423922 9606 423978
rect 9662 423922 9758 423978
rect 9138 406350 9758 423922
rect 9138 406294 9234 406350
rect 9290 406294 9358 406350
rect 9414 406294 9482 406350
rect 9538 406294 9606 406350
rect 9662 406294 9758 406350
rect 9138 406226 9758 406294
rect 9138 406170 9234 406226
rect 9290 406170 9358 406226
rect 9414 406170 9482 406226
rect 9538 406170 9606 406226
rect 9662 406170 9758 406226
rect 9138 406102 9758 406170
rect 9138 406046 9234 406102
rect 9290 406046 9358 406102
rect 9414 406046 9482 406102
rect 9538 406046 9606 406102
rect 9662 406046 9758 406102
rect 9138 405978 9758 406046
rect 9138 405922 9234 405978
rect 9290 405922 9358 405978
rect 9414 405922 9482 405978
rect 9538 405922 9606 405978
rect 9662 405922 9758 405978
rect 9138 388350 9758 405922
rect 9138 388294 9234 388350
rect 9290 388294 9358 388350
rect 9414 388294 9482 388350
rect 9538 388294 9606 388350
rect 9662 388294 9758 388350
rect 9138 388226 9758 388294
rect 9138 388170 9234 388226
rect 9290 388170 9358 388226
rect 9414 388170 9482 388226
rect 9538 388170 9606 388226
rect 9662 388170 9758 388226
rect 9138 388102 9758 388170
rect 9138 388046 9234 388102
rect 9290 388046 9358 388102
rect 9414 388046 9482 388102
rect 9538 388046 9606 388102
rect 9662 388046 9758 388102
rect 9138 387978 9758 388046
rect 9138 387922 9234 387978
rect 9290 387922 9358 387978
rect 9414 387922 9482 387978
rect 9538 387922 9606 387978
rect 9662 387922 9758 387978
rect 9138 370350 9758 387922
rect 9138 370294 9234 370350
rect 9290 370294 9358 370350
rect 9414 370294 9482 370350
rect 9538 370294 9606 370350
rect 9662 370294 9758 370350
rect 9138 370226 9758 370294
rect 9138 370170 9234 370226
rect 9290 370170 9358 370226
rect 9414 370170 9482 370226
rect 9538 370170 9606 370226
rect 9662 370170 9758 370226
rect 9138 370102 9758 370170
rect 9138 370046 9234 370102
rect 9290 370046 9358 370102
rect 9414 370046 9482 370102
rect 9538 370046 9606 370102
rect 9662 370046 9758 370102
rect 9138 369978 9758 370046
rect 9138 369922 9234 369978
rect 9290 369922 9358 369978
rect 9414 369922 9482 369978
rect 9538 369922 9606 369978
rect 9662 369922 9758 369978
rect 9138 352350 9758 369922
rect 9138 352294 9234 352350
rect 9290 352294 9358 352350
rect 9414 352294 9482 352350
rect 9538 352294 9606 352350
rect 9662 352294 9758 352350
rect 9138 352226 9758 352294
rect 9138 352170 9234 352226
rect 9290 352170 9358 352226
rect 9414 352170 9482 352226
rect 9538 352170 9606 352226
rect 9662 352170 9758 352226
rect 9138 352102 9758 352170
rect 9138 352046 9234 352102
rect 9290 352046 9358 352102
rect 9414 352046 9482 352102
rect 9538 352046 9606 352102
rect 9662 352046 9758 352102
rect 9138 351978 9758 352046
rect 9138 351922 9234 351978
rect 9290 351922 9358 351978
rect 9414 351922 9482 351978
rect 9538 351922 9606 351978
rect 9662 351922 9758 351978
rect 9138 334350 9758 351922
rect 9138 334294 9234 334350
rect 9290 334294 9358 334350
rect 9414 334294 9482 334350
rect 9538 334294 9606 334350
rect 9662 334294 9758 334350
rect 9138 334226 9758 334294
rect 9138 334170 9234 334226
rect 9290 334170 9358 334226
rect 9414 334170 9482 334226
rect 9538 334170 9606 334226
rect 9662 334170 9758 334226
rect 9138 334102 9758 334170
rect 9138 334046 9234 334102
rect 9290 334046 9358 334102
rect 9414 334046 9482 334102
rect 9538 334046 9606 334102
rect 9662 334046 9758 334102
rect 9138 333978 9758 334046
rect 9138 333922 9234 333978
rect 9290 333922 9358 333978
rect 9414 333922 9482 333978
rect 9538 333922 9606 333978
rect 9662 333922 9758 333978
rect 9138 316350 9758 333922
rect 9138 316294 9234 316350
rect 9290 316294 9358 316350
rect 9414 316294 9482 316350
rect 9538 316294 9606 316350
rect 9662 316294 9758 316350
rect 9138 316226 9758 316294
rect 9138 316170 9234 316226
rect 9290 316170 9358 316226
rect 9414 316170 9482 316226
rect 9538 316170 9606 316226
rect 9662 316170 9758 316226
rect 9138 316102 9758 316170
rect 9138 316046 9234 316102
rect 9290 316046 9358 316102
rect 9414 316046 9482 316102
rect 9538 316046 9606 316102
rect 9662 316046 9758 316102
rect 9138 315978 9758 316046
rect 9138 315922 9234 315978
rect 9290 315922 9358 315978
rect 9414 315922 9482 315978
rect 9538 315922 9606 315978
rect 9662 315922 9758 315978
rect 9138 298350 9758 315922
rect 9138 298294 9234 298350
rect 9290 298294 9358 298350
rect 9414 298294 9482 298350
rect 9538 298294 9606 298350
rect 9662 298294 9758 298350
rect 9138 298226 9758 298294
rect 9138 298170 9234 298226
rect 9290 298170 9358 298226
rect 9414 298170 9482 298226
rect 9538 298170 9606 298226
rect 9662 298170 9758 298226
rect 9138 298102 9758 298170
rect 9138 298046 9234 298102
rect 9290 298046 9358 298102
rect 9414 298046 9482 298102
rect 9538 298046 9606 298102
rect 9662 298046 9758 298102
rect 9138 297978 9758 298046
rect 9138 297922 9234 297978
rect 9290 297922 9358 297978
rect 9414 297922 9482 297978
rect 9538 297922 9606 297978
rect 9662 297922 9758 297978
rect 9138 280350 9758 297922
rect 9138 280294 9234 280350
rect 9290 280294 9358 280350
rect 9414 280294 9482 280350
rect 9538 280294 9606 280350
rect 9662 280294 9758 280350
rect 9138 280226 9758 280294
rect 9138 280170 9234 280226
rect 9290 280170 9358 280226
rect 9414 280170 9482 280226
rect 9538 280170 9606 280226
rect 9662 280170 9758 280226
rect 9138 280102 9758 280170
rect 9138 280046 9234 280102
rect 9290 280046 9358 280102
rect 9414 280046 9482 280102
rect 9538 280046 9606 280102
rect 9662 280046 9758 280102
rect 9138 279978 9758 280046
rect 9138 279922 9234 279978
rect 9290 279922 9358 279978
rect 9414 279922 9482 279978
rect 9538 279922 9606 279978
rect 9662 279922 9758 279978
rect 9138 262350 9758 279922
rect 9138 262294 9234 262350
rect 9290 262294 9358 262350
rect 9414 262294 9482 262350
rect 9538 262294 9606 262350
rect 9662 262294 9758 262350
rect 9138 262226 9758 262294
rect 9138 262170 9234 262226
rect 9290 262170 9358 262226
rect 9414 262170 9482 262226
rect 9538 262170 9606 262226
rect 9662 262170 9758 262226
rect 9138 262102 9758 262170
rect 9138 262046 9234 262102
rect 9290 262046 9358 262102
rect 9414 262046 9482 262102
rect 9538 262046 9606 262102
rect 9662 262046 9758 262102
rect 9138 261978 9758 262046
rect 9138 261922 9234 261978
rect 9290 261922 9358 261978
rect 9414 261922 9482 261978
rect 9538 261922 9606 261978
rect 9662 261922 9758 261978
rect 9138 244350 9758 261922
rect 9138 244294 9234 244350
rect 9290 244294 9358 244350
rect 9414 244294 9482 244350
rect 9538 244294 9606 244350
rect 9662 244294 9758 244350
rect 9138 244226 9758 244294
rect 9138 244170 9234 244226
rect 9290 244170 9358 244226
rect 9414 244170 9482 244226
rect 9538 244170 9606 244226
rect 9662 244170 9758 244226
rect 9138 244102 9758 244170
rect 9138 244046 9234 244102
rect 9290 244046 9358 244102
rect 9414 244046 9482 244102
rect 9538 244046 9606 244102
rect 9662 244046 9758 244102
rect 9138 243978 9758 244046
rect 9138 243922 9234 243978
rect 9290 243922 9358 243978
rect 9414 243922 9482 243978
rect 9538 243922 9606 243978
rect 9662 243922 9758 243978
rect 9138 226350 9758 243922
rect 9138 226294 9234 226350
rect 9290 226294 9358 226350
rect 9414 226294 9482 226350
rect 9538 226294 9606 226350
rect 9662 226294 9758 226350
rect 9138 226226 9758 226294
rect 9138 226170 9234 226226
rect 9290 226170 9358 226226
rect 9414 226170 9482 226226
rect 9538 226170 9606 226226
rect 9662 226170 9758 226226
rect 9138 226102 9758 226170
rect 9138 226046 9234 226102
rect 9290 226046 9358 226102
rect 9414 226046 9482 226102
rect 9538 226046 9606 226102
rect 9662 226046 9758 226102
rect 9138 225978 9758 226046
rect 9138 225922 9234 225978
rect 9290 225922 9358 225978
rect 9414 225922 9482 225978
rect 9538 225922 9606 225978
rect 9662 225922 9758 225978
rect 9138 208350 9758 225922
rect 9138 208294 9234 208350
rect 9290 208294 9358 208350
rect 9414 208294 9482 208350
rect 9538 208294 9606 208350
rect 9662 208294 9758 208350
rect 9138 208226 9758 208294
rect 9138 208170 9234 208226
rect 9290 208170 9358 208226
rect 9414 208170 9482 208226
rect 9538 208170 9606 208226
rect 9662 208170 9758 208226
rect 9138 208102 9758 208170
rect 9138 208046 9234 208102
rect 9290 208046 9358 208102
rect 9414 208046 9482 208102
rect 9538 208046 9606 208102
rect 9662 208046 9758 208102
rect 9138 207978 9758 208046
rect 9138 207922 9234 207978
rect 9290 207922 9358 207978
rect 9414 207922 9482 207978
rect 9538 207922 9606 207978
rect 9662 207922 9758 207978
rect 9138 190350 9758 207922
rect 9138 190294 9234 190350
rect 9290 190294 9358 190350
rect 9414 190294 9482 190350
rect 9538 190294 9606 190350
rect 9662 190294 9758 190350
rect 9138 190226 9758 190294
rect 9138 190170 9234 190226
rect 9290 190170 9358 190226
rect 9414 190170 9482 190226
rect 9538 190170 9606 190226
rect 9662 190170 9758 190226
rect 9138 190102 9758 190170
rect 9138 190046 9234 190102
rect 9290 190046 9358 190102
rect 9414 190046 9482 190102
rect 9538 190046 9606 190102
rect 9662 190046 9758 190102
rect 9138 189978 9758 190046
rect 9138 189922 9234 189978
rect 9290 189922 9358 189978
rect 9414 189922 9482 189978
rect 9538 189922 9606 189978
rect 9662 189922 9758 189978
rect 9138 172350 9758 189922
rect 9138 172294 9234 172350
rect 9290 172294 9358 172350
rect 9414 172294 9482 172350
rect 9538 172294 9606 172350
rect 9662 172294 9758 172350
rect 9138 172226 9758 172294
rect 9138 172170 9234 172226
rect 9290 172170 9358 172226
rect 9414 172170 9482 172226
rect 9538 172170 9606 172226
rect 9662 172170 9758 172226
rect 9138 172102 9758 172170
rect 9138 172046 9234 172102
rect 9290 172046 9358 172102
rect 9414 172046 9482 172102
rect 9538 172046 9606 172102
rect 9662 172046 9758 172102
rect 9138 171978 9758 172046
rect 9138 171922 9234 171978
rect 9290 171922 9358 171978
rect 9414 171922 9482 171978
rect 9538 171922 9606 171978
rect 9662 171922 9758 171978
rect 9138 154350 9758 171922
rect 9138 154294 9234 154350
rect 9290 154294 9358 154350
rect 9414 154294 9482 154350
rect 9538 154294 9606 154350
rect 9662 154294 9758 154350
rect 9138 154226 9758 154294
rect 9138 154170 9234 154226
rect 9290 154170 9358 154226
rect 9414 154170 9482 154226
rect 9538 154170 9606 154226
rect 9662 154170 9758 154226
rect 9138 154102 9758 154170
rect 9138 154046 9234 154102
rect 9290 154046 9358 154102
rect 9414 154046 9482 154102
rect 9538 154046 9606 154102
rect 9662 154046 9758 154102
rect 9138 153978 9758 154046
rect 9138 153922 9234 153978
rect 9290 153922 9358 153978
rect 9414 153922 9482 153978
rect 9538 153922 9606 153978
rect 9662 153922 9758 153978
rect 9138 136350 9758 153922
rect 9138 136294 9234 136350
rect 9290 136294 9358 136350
rect 9414 136294 9482 136350
rect 9538 136294 9606 136350
rect 9662 136294 9758 136350
rect 9138 136226 9758 136294
rect 9138 136170 9234 136226
rect 9290 136170 9358 136226
rect 9414 136170 9482 136226
rect 9538 136170 9606 136226
rect 9662 136170 9758 136226
rect 9138 136102 9758 136170
rect 9138 136046 9234 136102
rect 9290 136046 9358 136102
rect 9414 136046 9482 136102
rect 9538 136046 9606 136102
rect 9662 136046 9758 136102
rect 9138 135978 9758 136046
rect 9138 135922 9234 135978
rect 9290 135922 9358 135978
rect 9414 135922 9482 135978
rect 9538 135922 9606 135978
rect 9662 135922 9758 135978
rect 9138 118350 9758 135922
rect 9138 118294 9234 118350
rect 9290 118294 9358 118350
rect 9414 118294 9482 118350
rect 9538 118294 9606 118350
rect 9662 118294 9758 118350
rect 9138 118226 9758 118294
rect 9138 118170 9234 118226
rect 9290 118170 9358 118226
rect 9414 118170 9482 118226
rect 9538 118170 9606 118226
rect 9662 118170 9758 118226
rect 9138 118102 9758 118170
rect 9138 118046 9234 118102
rect 9290 118046 9358 118102
rect 9414 118046 9482 118102
rect 9538 118046 9606 118102
rect 9662 118046 9758 118102
rect 9138 117978 9758 118046
rect 9138 117922 9234 117978
rect 9290 117922 9358 117978
rect 9414 117922 9482 117978
rect 9538 117922 9606 117978
rect 9662 117922 9758 117978
rect 8652 105028 8708 105038
rect 8316 59938 8372 59948
rect 8540 72996 8596 73006
rect 8092 33058 8148 33068
rect 8540 16100 8596 72940
rect 8652 68068 8708 104972
rect 9138 100350 9758 117922
rect 9138 100294 9234 100350
rect 9290 100294 9358 100350
rect 9414 100294 9482 100350
rect 9538 100294 9606 100350
rect 9662 100294 9758 100350
rect 9138 100226 9758 100294
rect 9138 100170 9234 100226
rect 9290 100170 9358 100226
rect 9414 100170 9482 100226
rect 9538 100170 9606 100226
rect 9662 100170 9758 100226
rect 9138 100102 9758 100170
rect 9138 100046 9234 100102
rect 9290 100046 9358 100102
rect 9414 100046 9482 100102
rect 9538 100046 9606 100102
rect 9662 100046 9758 100102
rect 9138 99978 9758 100046
rect 9138 99922 9234 99978
rect 9290 99922 9358 99978
rect 9414 99922 9482 99978
rect 9538 99922 9606 99978
rect 9662 99922 9758 99978
rect 9138 82350 9758 99922
rect 9138 82294 9234 82350
rect 9290 82294 9358 82350
rect 9414 82294 9482 82350
rect 9538 82294 9606 82350
rect 9662 82294 9758 82350
rect 9138 82226 9758 82294
rect 9138 82170 9234 82226
rect 9290 82170 9358 82226
rect 9414 82170 9482 82226
rect 9538 82170 9606 82226
rect 9662 82170 9758 82226
rect 9138 82102 9758 82170
rect 9138 82046 9234 82102
rect 9290 82046 9358 82102
rect 9414 82046 9482 82102
rect 9538 82046 9606 82102
rect 9662 82046 9758 82102
rect 9138 81978 9758 82046
rect 9138 81922 9234 81978
rect 9290 81922 9358 81978
rect 9414 81922 9482 81978
rect 9538 81922 9606 81978
rect 9662 81922 9758 81978
rect 8652 68002 8708 68012
rect 8764 74004 8820 74014
rect 8540 16034 8596 16044
rect 8764 10724 8820 73948
rect 8988 72118 9044 72128
rect 8876 68878 8932 68888
rect 8876 21476 8932 68822
rect 8988 24164 9044 72062
rect 8988 24098 9044 24108
rect 9138 64350 9758 81922
rect 10892 558964 10948 558974
rect 9884 81508 9940 81518
rect 9884 70756 9940 81452
rect 9884 70690 9940 70700
rect 9996 74788 10052 74798
rect 9996 69860 10052 74732
rect 9996 69794 10052 69804
rect 9996 69636 10052 69646
rect 9996 67172 10052 69580
rect 9996 67106 10052 67116
rect 9138 64294 9234 64350
rect 9290 64294 9358 64350
rect 9414 64294 9482 64350
rect 9538 64294 9606 64350
rect 9662 64294 9758 64350
rect 9138 64226 9758 64294
rect 9138 64170 9234 64226
rect 9290 64170 9358 64226
rect 9414 64170 9482 64226
rect 9538 64170 9606 64226
rect 9662 64170 9758 64226
rect 9138 64102 9758 64170
rect 9138 64046 9234 64102
rect 9290 64046 9358 64102
rect 9414 64046 9482 64102
rect 9538 64046 9606 64102
rect 9662 64046 9758 64102
rect 9138 63978 9758 64046
rect 9138 63922 9234 63978
rect 9290 63922 9358 63978
rect 9414 63922 9482 63978
rect 9538 63922 9606 63978
rect 9662 63922 9758 63978
rect 9138 46350 9758 63922
rect 9996 65604 10052 65614
rect 9996 60900 10052 65548
rect 9996 60834 10052 60844
rect 9138 46294 9234 46350
rect 9290 46294 9358 46350
rect 9414 46294 9482 46350
rect 9538 46294 9606 46350
rect 9662 46294 9758 46350
rect 9138 46226 9758 46294
rect 9138 46170 9234 46226
rect 9290 46170 9358 46226
rect 9414 46170 9482 46226
rect 9538 46170 9606 46226
rect 9662 46170 9758 46226
rect 9138 46102 9758 46170
rect 9138 46046 9234 46102
rect 9290 46046 9358 46102
rect 9414 46046 9482 46102
rect 9538 46046 9606 46102
rect 9662 46046 9758 46102
rect 9138 45978 9758 46046
rect 9138 45922 9234 45978
rect 9290 45922 9358 45978
rect 9414 45922 9482 45978
rect 9538 45922 9606 45978
rect 9662 45922 9758 45978
rect 9138 28350 9758 45922
rect 9996 49618 10052 49628
rect 9996 44772 10052 49562
rect 9996 44706 10052 44716
rect 9138 28294 9234 28350
rect 9290 28294 9358 28350
rect 9414 28294 9482 28350
rect 9538 28294 9606 28350
rect 9662 28294 9758 28350
rect 9138 28226 9758 28294
rect 9138 28170 9234 28226
rect 9290 28170 9358 28226
rect 9414 28170 9482 28226
rect 9538 28170 9606 28226
rect 9662 28170 9758 28226
rect 9138 28102 9758 28170
rect 9138 28046 9234 28102
rect 9290 28046 9358 28102
rect 9414 28046 9482 28102
rect 9538 28046 9606 28102
rect 9662 28046 9758 28102
rect 9138 27978 9758 28046
rect 9138 27922 9234 27978
rect 9290 27922 9358 27978
rect 9414 27922 9482 27978
rect 9538 27922 9606 27978
rect 9662 27922 9758 27978
rect 8876 21410 8932 21420
rect 8764 10658 8820 10668
rect 7756 7074 7812 7084
rect 9138 10350 9758 27922
rect 10892 25956 10948 558908
rect 11900 516628 11956 516638
rect 11676 430164 11732 430174
rect 10892 25890 10948 25900
rect 11004 304164 11060 304174
rect 11004 18788 11060 304108
rect 11676 78988 11732 430108
rect 11340 78932 11732 78988
rect 11788 319060 11844 319070
rect 11340 63588 11396 78932
rect 11340 63522 11396 63532
rect 11452 78058 11508 78068
rect 11452 57316 11508 78002
rect 11452 57250 11508 57260
rect 11564 74818 11620 74828
rect 11564 35812 11620 74762
rect 11788 74004 11844 319004
rect 11788 73938 11844 73948
rect 11564 35746 11620 35756
rect 11900 26578 11956 516572
rect 12012 67228 12068 573020
rect 15148 530740 15204 530750
rect 14252 509348 14308 509358
rect 13468 488404 13524 488414
rect 12684 69058 12740 69068
rect 12684 68964 12740 69002
rect 12684 68898 12740 68908
rect 13468 68878 13524 488348
rect 13580 403732 13636 403742
rect 13580 72996 13636 403676
rect 13580 72930 13636 72940
rect 13468 68812 13524 68822
rect 12012 67172 12180 67228
rect 12124 31948 12180 67172
rect 12684 67078 12740 67088
rect 12572 67022 12684 67078
rect 12572 66948 12628 67022
rect 12684 67012 12740 67022
rect 12572 66882 12628 66892
rect 12460 65458 12516 65468
rect 12460 65044 12516 65402
rect 12460 64978 12516 64988
rect 12460 63658 12516 63668
rect 12460 63364 12516 63602
rect 12460 63298 12516 63308
rect 12684 62038 12740 62048
rect 12684 61796 12740 61982
rect 12684 61730 12740 61740
rect 12684 60778 12740 60788
rect 12572 60722 12684 60778
rect 12460 60418 12516 60428
rect 12460 59668 12516 60362
rect 12460 59602 12516 59612
rect 12572 58772 12628 60722
rect 12684 60712 12740 60722
rect 14252 60778 14308 509292
rect 15148 72118 15204 530684
rect 15148 72052 15204 72062
rect 15932 350756 15988 350766
rect 15932 69058 15988 350700
rect 15932 68992 15988 69002
rect 14252 60712 14308 60722
rect 12572 58706 12628 58716
rect 16448 58350 16768 58384
rect 16448 58294 16518 58350
rect 16574 58294 16642 58350
rect 16698 58294 16768 58350
rect 16448 58226 16768 58294
rect 16448 58170 16518 58226
rect 16574 58170 16642 58226
rect 16698 58170 16768 58226
rect 16448 58102 16768 58170
rect 16448 58046 16518 58102
rect 16574 58046 16642 58102
rect 16698 58046 16768 58102
rect 16448 57978 16768 58046
rect 16448 57922 16518 57978
rect 16574 57922 16642 57978
rect 16698 57922 16768 57978
rect 16448 57888 16768 57922
rect 12348 56998 12404 57008
rect 12348 56196 12404 56942
rect 12348 56130 12404 56140
rect 12348 54658 12404 54668
rect 12348 53508 12404 54602
rect 12684 53758 12740 53768
rect 17612 53758 17668 575372
rect 17612 53692 17668 53702
rect 12684 53664 12740 53676
rect 12348 53442 12404 53452
rect 12348 51958 12404 51968
rect 12348 51716 12404 51902
rect 12348 51650 12404 51660
rect 12684 48718 12740 48728
rect 12684 48356 12740 48662
rect 19292 48718 19348 578732
rect 20972 456484 21028 456494
rect 20972 62038 21028 456428
rect 21084 337540 21140 337550
rect 21084 74788 21140 337484
rect 21084 74722 21140 74732
rect 20972 61972 21028 61982
rect 22652 51958 22708 582092
rect 24332 548996 24388 549006
rect 24332 56998 24388 548940
rect 24332 56932 24388 56942
rect 26012 54658 26068 588588
rect 26012 54592 26068 54602
rect 22652 51892 22708 51902
rect 27692 49618 27748 590604
rect 36138 580350 36758 596784
rect 36138 580294 36234 580350
rect 36290 580294 36358 580350
rect 36414 580294 36482 580350
rect 36538 580294 36606 580350
rect 36662 580294 36758 580350
rect 36138 580226 36758 580294
rect 36138 580170 36234 580226
rect 36290 580170 36358 580226
rect 36414 580170 36482 580226
rect 36538 580170 36606 580226
rect 36662 580170 36758 580226
rect 36138 580102 36758 580170
rect 36138 580046 36234 580102
rect 36290 580046 36358 580102
rect 36414 580046 36482 580102
rect 36538 580046 36606 580102
rect 36662 580046 36758 580102
rect 36138 579978 36758 580046
rect 36138 579922 36234 579978
rect 36290 579922 36358 579978
rect 36414 579922 36482 579978
rect 36538 579922 36606 579978
rect 36662 579922 36758 579978
rect 36138 562350 36758 579922
rect 36138 562294 36234 562350
rect 36290 562294 36358 562350
rect 36414 562294 36482 562350
rect 36538 562294 36606 562350
rect 36662 562294 36758 562350
rect 36138 562226 36758 562294
rect 36138 562170 36234 562226
rect 36290 562170 36358 562226
rect 36414 562170 36482 562226
rect 36538 562170 36606 562226
rect 36662 562170 36758 562226
rect 36138 562102 36758 562170
rect 36138 562046 36234 562102
rect 36290 562046 36358 562102
rect 36414 562046 36482 562102
rect 36538 562046 36606 562102
rect 36662 562046 36758 562102
rect 36138 561978 36758 562046
rect 36138 561922 36234 561978
rect 36290 561922 36358 561978
rect 36414 561922 36482 561978
rect 36538 561922 36606 561978
rect 36662 561922 36758 561978
rect 36138 544350 36758 561922
rect 36138 544294 36234 544350
rect 36290 544294 36358 544350
rect 36414 544294 36482 544350
rect 36538 544294 36606 544350
rect 36662 544294 36758 544350
rect 36138 544226 36758 544294
rect 36138 544170 36234 544226
rect 36290 544170 36358 544226
rect 36414 544170 36482 544226
rect 36538 544170 36606 544226
rect 36662 544170 36758 544226
rect 36138 544102 36758 544170
rect 36138 544046 36234 544102
rect 36290 544046 36358 544102
rect 36414 544046 36482 544102
rect 36538 544046 36606 544102
rect 36662 544046 36758 544102
rect 36138 543978 36758 544046
rect 36138 543922 36234 543978
rect 36290 543922 36358 543978
rect 36414 543922 36482 543978
rect 36538 543922 36606 543978
rect 36662 543922 36758 543978
rect 36138 526350 36758 543922
rect 36138 526294 36234 526350
rect 36290 526294 36358 526350
rect 36414 526294 36482 526350
rect 36538 526294 36606 526350
rect 36662 526294 36758 526350
rect 36138 526226 36758 526294
rect 36138 526170 36234 526226
rect 36290 526170 36358 526226
rect 36414 526170 36482 526226
rect 36538 526170 36606 526226
rect 36662 526170 36758 526226
rect 36138 526102 36758 526170
rect 36138 526046 36234 526102
rect 36290 526046 36358 526102
rect 36414 526046 36482 526102
rect 36538 526046 36606 526102
rect 36662 526046 36758 526102
rect 36138 525978 36758 526046
rect 36138 525922 36234 525978
rect 36290 525922 36358 525978
rect 36414 525922 36482 525978
rect 36538 525922 36606 525978
rect 36662 525922 36758 525978
rect 36138 508350 36758 525922
rect 36138 508294 36234 508350
rect 36290 508294 36358 508350
rect 36414 508294 36482 508350
rect 36538 508294 36606 508350
rect 36662 508294 36758 508350
rect 36138 508226 36758 508294
rect 36138 508170 36234 508226
rect 36290 508170 36358 508226
rect 36414 508170 36482 508226
rect 36538 508170 36606 508226
rect 36662 508170 36758 508226
rect 36138 508102 36758 508170
rect 36138 508046 36234 508102
rect 36290 508046 36358 508102
rect 36414 508046 36482 508102
rect 36538 508046 36606 508102
rect 36662 508046 36758 508102
rect 36138 507978 36758 508046
rect 36138 507922 36234 507978
rect 36290 507922 36358 507978
rect 36414 507922 36482 507978
rect 36538 507922 36606 507978
rect 36662 507922 36758 507978
rect 31052 494788 31108 494798
rect 29372 390404 29428 390414
rect 29372 67078 29428 390348
rect 29372 67012 29428 67022
rect 31052 60418 31108 494732
rect 36138 490350 36758 507922
rect 36138 490294 36234 490350
rect 36290 490294 36358 490350
rect 36414 490294 36482 490350
rect 36538 490294 36606 490350
rect 36662 490294 36758 490350
rect 36138 490226 36758 490294
rect 36138 490170 36234 490226
rect 36290 490170 36358 490226
rect 36414 490170 36482 490226
rect 36538 490170 36606 490226
rect 36662 490170 36758 490226
rect 36138 490102 36758 490170
rect 36138 490046 36234 490102
rect 36290 490046 36358 490102
rect 36414 490046 36482 490102
rect 36538 490046 36606 490102
rect 36662 490046 36758 490102
rect 36138 489978 36758 490046
rect 36138 489922 36234 489978
rect 36290 489922 36358 489978
rect 36414 489922 36482 489978
rect 36538 489922 36606 489978
rect 36662 489922 36758 489978
rect 36138 472350 36758 489922
rect 36138 472294 36234 472350
rect 36290 472294 36358 472350
rect 36414 472294 36482 472350
rect 36538 472294 36606 472350
rect 36662 472294 36758 472350
rect 36138 472226 36758 472294
rect 36138 472170 36234 472226
rect 36290 472170 36358 472226
rect 36414 472170 36482 472226
rect 36538 472170 36606 472226
rect 36662 472170 36758 472226
rect 36138 472102 36758 472170
rect 36138 472046 36234 472102
rect 36290 472046 36358 472102
rect 36414 472046 36482 472102
rect 36538 472046 36606 472102
rect 36662 472046 36758 472102
rect 36138 471978 36758 472046
rect 36138 471922 36234 471978
rect 36290 471922 36358 471978
rect 36414 471922 36482 471978
rect 36538 471922 36606 471978
rect 36662 471922 36758 471978
rect 36138 454350 36758 471922
rect 36138 454294 36234 454350
rect 36290 454294 36358 454350
rect 36414 454294 36482 454350
rect 36538 454294 36606 454350
rect 36662 454294 36758 454350
rect 36138 454226 36758 454294
rect 36138 454170 36234 454226
rect 36290 454170 36358 454226
rect 36414 454170 36482 454226
rect 36538 454170 36606 454226
rect 36662 454170 36758 454226
rect 36138 454102 36758 454170
rect 36138 454046 36234 454102
rect 36290 454046 36358 454102
rect 36414 454046 36482 454102
rect 36538 454046 36606 454102
rect 36662 454046 36758 454102
rect 36138 453978 36758 454046
rect 36138 453922 36234 453978
rect 36290 453922 36358 453978
rect 36414 453922 36482 453978
rect 36538 453922 36606 453978
rect 36662 453922 36758 453978
rect 36138 436350 36758 453922
rect 36138 436294 36234 436350
rect 36290 436294 36358 436350
rect 36414 436294 36482 436350
rect 36538 436294 36606 436350
rect 36662 436294 36758 436350
rect 36138 436226 36758 436294
rect 36138 436170 36234 436226
rect 36290 436170 36358 436226
rect 36414 436170 36482 436226
rect 36538 436170 36606 436226
rect 36662 436170 36758 436226
rect 36138 436102 36758 436170
rect 36138 436046 36234 436102
rect 36290 436046 36358 436102
rect 36414 436046 36482 436102
rect 36538 436046 36606 436102
rect 36662 436046 36758 436102
rect 36138 435978 36758 436046
rect 36138 435922 36234 435978
rect 36290 435922 36358 435978
rect 36414 435922 36482 435978
rect 36538 435922 36606 435978
rect 36662 435922 36758 435978
rect 36138 418350 36758 435922
rect 36138 418294 36234 418350
rect 36290 418294 36358 418350
rect 36414 418294 36482 418350
rect 36538 418294 36606 418350
rect 36662 418294 36758 418350
rect 36138 418226 36758 418294
rect 36138 418170 36234 418226
rect 36290 418170 36358 418226
rect 36414 418170 36482 418226
rect 36538 418170 36606 418226
rect 36662 418170 36758 418226
rect 36138 418102 36758 418170
rect 36138 418046 36234 418102
rect 36290 418046 36358 418102
rect 36414 418046 36482 418102
rect 36538 418046 36606 418102
rect 36662 418046 36758 418102
rect 36138 417978 36758 418046
rect 36138 417922 36234 417978
rect 36290 417922 36358 417978
rect 36414 417922 36482 417978
rect 36538 417922 36606 417978
rect 36662 417922 36758 417978
rect 36138 400350 36758 417922
rect 36138 400294 36234 400350
rect 36290 400294 36358 400350
rect 36414 400294 36482 400350
rect 36538 400294 36606 400350
rect 36662 400294 36758 400350
rect 36138 400226 36758 400294
rect 36138 400170 36234 400226
rect 36290 400170 36358 400226
rect 36414 400170 36482 400226
rect 36538 400170 36606 400226
rect 36662 400170 36758 400226
rect 36138 400102 36758 400170
rect 36138 400046 36234 400102
rect 36290 400046 36358 400102
rect 36414 400046 36482 400102
rect 36538 400046 36606 400102
rect 36662 400046 36758 400102
rect 36138 399978 36758 400046
rect 36138 399922 36234 399978
rect 36290 399922 36358 399978
rect 36414 399922 36482 399978
rect 36538 399922 36606 399978
rect 36662 399922 36758 399978
rect 36138 382350 36758 399922
rect 36138 382294 36234 382350
rect 36290 382294 36358 382350
rect 36414 382294 36482 382350
rect 36538 382294 36606 382350
rect 36662 382294 36758 382350
rect 36138 382226 36758 382294
rect 36138 382170 36234 382226
rect 36290 382170 36358 382226
rect 36414 382170 36482 382226
rect 36538 382170 36606 382226
rect 36662 382170 36758 382226
rect 36138 382102 36758 382170
rect 36138 382046 36234 382102
rect 36290 382046 36358 382102
rect 36414 382046 36482 382102
rect 36538 382046 36606 382102
rect 36662 382046 36758 382102
rect 36138 381978 36758 382046
rect 36138 381922 36234 381978
rect 36290 381922 36358 381978
rect 36414 381922 36482 381978
rect 36538 381922 36606 381978
rect 36662 381922 36758 381978
rect 36138 364350 36758 381922
rect 36138 364294 36234 364350
rect 36290 364294 36358 364350
rect 36414 364294 36482 364350
rect 36538 364294 36606 364350
rect 36662 364294 36758 364350
rect 36138 364226 36758 364294
rect 36138 364170 36234 364226
rect 36290 364170 36358 364226
rect 36414 364170 36482 364226
rect 36538 364170 36606 364226
rect 36662 364170 36758 364226
rect 36138 364102 36758 364170
rect 36138 364046 36234 364102
rect 36290 364046 36358 364102
rect 36414 364046 36482 364102
rect 36538 364046 36606 364102
rect 36662 364046 36758 364102
rect 36138 363978 36758 364046
rect 36138 363922 36234 363978
rect 36290 363922 36358 363978
rect 36414 363922 36482 363978
rect 36538 363922 36606 363978
rect 36662 363922 36758 363978
rect 36138 346350 36758 363922
rect 36138 346294 36234 346350
rect 36290 346294 36358 346350
rect 36414 346294 36482 346350
rect 36538 346294 36606 346350
rect 36662 346294 36758 346350
rect 36138 346226 36758 346294
rect 36138 346170 36234 346226
rect 36290 346170 36358 346226
rect 36414 346170 36482 346226
rect 36538 346170 36606 346226
rect 36662 346170 36758 346226
rect 36138 346102 36758 346170
rect 36138 346046 36234 346102
rect 36290 346046 36358 346102
rect 36414 346046 36482 346102
rect 36538 346046 36606 346102
rect 36662 346046 36758 346102
rect 36138 345978 36758 346046
rect 36138 345922 36234 345978
rect 36290 345922 36358 345978
rect 36414 345922 36482 345978
rect 36538 345922 36606 345978
rect 36662 345922 36758 345978
rect 36138 328350 36758 345922
rect 36138 328294 36234 328350
rect 36290 328294 36358 328350
rect 36414 328294 36482 328350
rect 36538 328294 36606 328350
rect 36662 328294 36758 328350
rect 36138 328226 36758 328294
rect 36138 328170 36234 328226
rect 36290 328170 36358 328226
rect 36414 328170 36482 328226
rect 36538 328170 36606 328226
rect 36662 328170 36758 328226
rect 36138 328102 36758 328170
rect 36138 328046 36234 328102
rect 36290 328046 36358 328102
rect 36414 328046 36482 328102
rect 36538 328046 36606 328102
rect 36662 328046 36758 328102
rect 36138 327978 36758 328046
rect 36138 327922 36234 327978
rect 36290 327922 36358 327978
rect 36414 327922 36482 327978
rect 36538 327922 36606 327978
rect 36662 327922 36758 327978
rect 36138 310350 36758 327922
rect 36138 310294 36234 310350
rect 36290 310294 36358 310350
rect 36414 310294 36482 310350
rect 36538 310294 36606 310350
rect 36662 310294 36758 310350
rect 36138 310226 36758 310294
rect 36138 310170 36234 310226
rect 36290 310170 36358 310226
rect 36414 310170 36482 310226
rect 36538 310170 36606 310226
rect 36662 310170 36758 310226
rect 36138 310102 36758 310170
rect 36138 310046 36234 310102
rect 36290 310046 36358 310102
rect 36414 310046 36482 310102
rect 36538 310046 36606 310102
rect 36662 310046 36758 310102
rect 36138 309978 36758 310046
rect 36138 309922 36234 309978
rect 36290 309922 36358 309978
rect 36414 309922 36482 309978
rect 36538 309922 36606 309978
rect 36662 309922 36758 309978
rect 36138 292350 36758 309922
rect 36138 292294 36234 292350
rect 36290 292294 36358 292350
rect 36414 292294 36482 292350
rect 36538 292294 36606 292350
rect 36662 292294 36758 292350
rect 36138 292226 36758 292294
rect 36138 292170 36234 292226
rect 36290 292170 36358 292226
rect 36414 292170 36482 292226
rect 36538 292170 36606 292226
rect 36662 292170 36758 292226
rect 36138 292102 36758 292170
rect 36138 292046 36234 292102
rect 36290 292046 36358 292102
rect 36414 292046 36482 292102
rect 36538 292046 36606 292102
rect 36662 292046 36758 292102
rect 36138 291978 36758 292046
rect 36138 291922 36234 291978
rect 36290 291922 36358 291978
rect 36414 291922 36482 291978
rect 36538 291922 36606 291978
rect 36662 291922 36758 291978
rect 36138 274350 36758 291922
rect 36138 274294 36234 274350
rect 36290 274294 36358 274350
rect 36414 274294 36482 274350
rect 36538 274294 36606 274350
rect 36662 274294 36758 274350
rect 36138 274226 36758 274294
rect 36138 274170 36234 274226
rect 36290 274170 36358 274226
rect 36414 274170 36482 274226
rect 36538 274170 36606 274226
rect 36662 274170 36758 274226
rect 36138 274102 36758 274170
rect 36138 274046 36234 274102
rect 36290 274046 36358 274102
rect 36414 274046 36482 274102
rect 36538 274046 36606 274102
rect 36662 274046 36758 274102
rect 36138 273978 36758 274046
rect 36138 273922 36234 273978
rect 36290 273922 36358 273978
rect 36414 273922 36482 273978
rect 36538 273922 36606 273978
rect 36662 273922 36758 273978
rect 36138 256350 36758 273922
rect 36138 256294 36234 256350
rect 36290 256294 36358 256350
rect 36414 256294 36482 256350
rect 36538 256294 36606 256350
rect 36662 256294 36758 256350
rect 36138 256226 36758 256294
rect 36138 256170 36234 256226
rect 36290 256170 36358 256226
rect 36414 256170 36482 256226
rect 36538 256170 36606 256226
rect 36662 256170 36758 256226
rect 36138 256102 36758 256170
rect 36138 256046 36234 256102
rect 36290 256046 36358 256102
rect 36414 256046 36482 256102
rect 36538 256046 36606 256102
rect 36662 256046 36758 256102
rect 36138 255978 36758 256046
rect 36138 255922 36234 255978
rect 36290 255922 36358 255978
rect 36414 255922 36482 255978
rect 36538 255922 36606 255978
rect 36662 255922 36758 255978
rect 36138 238350 36758 255922
rect 36138 238294 36234 238350
rect 36290 238294 36358 238350
rect 36414 238294 36482 238350
rect 36538 238294 36606 238350
rect 36662 238294 36758 238350
rect 36138 238226 36758 238294
rect 36138 238170 36234 238226
rect 36290 238170 36358 238226
rect 36414 238170 36482 238226
rect 36538 238170 36606 238226
rect 36662 238170 36758 238226
rect 36138 238102 36758 238170
rect 36138 238046 36234 238102
rect 36290 238046 36358 238102
rect 36414 238046 36482 238102
rect 36538 238046 36606 238102
rect 36662 238046 36758 238102
rect 36138 237978 36758 238046
rect 36138 237922 36234 237978
rect 36290 237922 36358 237978
rect 36414 237922 36482 237978
rect 36538 237922 36606 237978
rect 36662 237922 36758 237978
rect 36138 220350 36758 237922
rect 36138 220294 36234 220350
rect 36290 220294 36358 220350
rect 36414 220294 36482 220350
rect 36538 220294 36606 220350
rect 36662 220294 36758 220350
rect 36138 220226 36758 220294
rect 36138 220170 36234 220226
rect 36290 220170 36358 220226
rect 36414 220170 36482 220226
rect 36538 220170 36606 220226
rect 36662 220170 36758 220226
rect 36138 220102 36758 220170
rect 36138 220046 36234 220102
rect 36290 220046 36358 220102
rect 36414 220046 36482 220102
rect 36538 220046 36606 220102
rect 36662 220046 36758 220102
rect 36138 219978 36758 220046
rect 36138 219922 36234 219978
rect 36290 219922 36358 219978
rect 36414 219922 36482 219978
rect 36538 219922 36606 219978
rect 36662 219922 36758 219978
rect 36138 202350 36758 219922
rect 36138 202294 36234 202350
rect 36290 202294 36358 202350
rect 36414 202294 36482 202350
rect 36538 202294 36606 202350
rect 36662 202294 36758 202350
rect 36138 202226 36758 202294
rect 36138 202170 36234 202226
rect 36290 202170 36358 202226
rect 36414 202170 36482 202226
rect 36538 202170 36606 202226
rect 36662 202170 36758 202226
rect 36138 202102 36758 202170
rect 36138 202046 36234 202102
rect 36290 202046 36358 202102
rect 36414 202046 36482 202102
rect 36538 202046 36606 202102
rect 36662 202046 36758 202102
rect 36138 201978 36758 202046
rect 36138 201922 36234 201978
rect 36290 201922 36358 201978
rect 36414 201922 36482 201978
rect 36538 201922 36606 201978
rect 36662 201922 36758 201978
rect 36138 184350 36758 201922
rect 36138 184294 36234 184350
rect 36290 184294 36358 184350
rect 36414 184294 36482 184350
rect 36538 184294 36606 184350
rect 36662 184294 36758 184350
rect 36138 184226 36758 184294
rect 36138 184170 36234 184226
rect 36290 184170 36358 184226
rect 36414 184170 36482 184226
rect 36538 184170 36606 184226
rect 36662 184170 36758 184226
rect 36138 184102 36758 184170
rect 36138 184046 36234 184102
rect 36290 184046 36358 184102
rect 36414 184046 36482 184102
rect 36538 184046 36606 184102
rect 36662 184046 36758 184102
rect 36138 183978 36758 184046
rect 36138 183922 36234 183978
rect 36290 183922 36358 183978
rect 36414 183922 36482 183978
rect 36538 183922 36606 183978
rect 36662 183922 36758 183978
rect 36138 166350 36758 183922
rect 36138 166294 36234 166350
rect 36290 166294 36358 166350
rect 36414 166294 36482 166350
rect 36538 166294 36606 166350
rect 36662 166294 36758 166350
rect 36138 166226 36758 166294
rect 36138 166170 36234 166226
rect 36290 166170 36358 166226
rect 36414 166170 36482 166226
rect 36538 166170 36606 166226
rect 36662 166170 36758 166226
rect 36138 166102 36758 166170
rect 36138 166046 36234 166102
rect 36290 166046 36358 166102
rect 36414 166046 36482 166102
rect 36538 166046 36606 166102
rect 36662 166046 36758 166102
rect 36138 165978 36758 166046
rect 36138 165922 36234 165978
rect 36290 165922 36358 165978
rect 36414 165922 36482 165978
rect 36538 165922 36606 165978
rect 36662 165922 36758 165978
rect 36138 148350 36758 165922
rect 36138 148294 36234 148350
rect 36290 148294 36358 148350
rect 36414 148294 36482 148350
rect 36538 148294 36606 148350
rect 36662 148294 36758 148350
rect 36138 148226 36758 148294
rect 36138 148170 36234 148226
rect 36290 148170 36358 148226
rect 36414 148170 36482 148226
rect 36538 148170 36606 148226
rect 36662 148170 36758 148226
rect 36138 148102 36758 148170
rect 36138 148046 36234 148102
rect 36290 148046 36358 148102
rect 36414 148046 36482 148102
rect 36538 148046 36606 148102
rect 36662 148046 36758 148102
rect 36138 147978 36758 148046
rect 36138 147922 36234 147978
rect 36290 147922 36358 147978
rect 36414 147922 36482 147978
rect 36538 147922 36606 147978
rect 36662 147922 36758 147978
rect 36138 130350 36758 147922
rect 36138 130294 36234 130350
rect 36290 130294 36358 130350
rect 36414 130294 36482 130350
rect 36538 130294 36606 130350
rect 36662 130294 36758 130350
rect 36138 130226 36758 130294
rect 36138 130170 36234 130226
rect 36290 130170 36358 130226
rect 36414 130170 36482 130226
rect 36538 130170 36606 130226
rect 36662 130170 36758 130226
rect 36138 130102 36758 130170
rect 36138 130046 36234 130102
rect 36290 130046 36358 130102
rect 36414 130046 36482 130102
rect 36538 130046 36606 130102
rect 36662 130046 36758 130102
rect 36138 129978 36758 130046
rect 36138 129922 36234 129978
rect 36290 129922 36358 129978
rect 36414 129922 36482 129978
rect 36538 129922 36606 129978
rect 36662 129922 36758 129978
rect 36138 112350 36758 129922
rect 36138 112294 36234 112350
rect 36290 112294 36358 112350
rect 36414 112294 36482 112350
rect 36538 112294 36606 112350
rect 36662 112294 36758 112350
rect 36138 112226 36758 112294
rect 36138 112170 36234 112226
rect 36290 112170 36358 112226
rect 36414 112170 36482 112226
rect 36538 112170 36606 112226
rect 36662 112170 36758 112226
rect 36138 112102 36758 112170
rect 36138 112046 36234 112102
rect 36290 112046 36358 112102
rect 36414 112046 36482 112102
rect 36538 112046 36606 112102
rect 36662 112046 36758 112102
rect 36138 111978 36758 112046
rect 36138 111922 36234 111978
rect 36290 111922 36358 111978
rect 36414 111922 36482 111978
rect 36538 111922 36606 111978
rect 36662 111922 36758 111978
rect 36138 94350 36758 111922
rect 36138 94294 36234 94350
rect 36290 94294 36358 94350
rect 36414 94294 36482 94350
rect 36538 94294 36606 94350
rect 36662 94294 36758 94350
rect 36138 94226 36758 94294
rect 36138 94170 36234 94226
rect 36290 94170 36358 94226
rect 36414 94170 36482 94226
rect 36538 94170 36606 94226
rect 36662 94170 36758 94226
rect 36138 94102 36758 94170
rect 36138 94046 36234 94102
rect 36290 94046 36358 94102
rect 36414 94046 36482 94102
rect 36538 94046 36606 94102
rect 36662 94046 36758 94102
rect 36138 93978 36758 94046
rect 36138 93922 36234 93978
rect 36290 93922 36358 93978
rect 36414 93922 36482 93978
rect 36538 93922 36606 93978
rect 36662 93922 36758 93978
rect 36138 76350 36758 93922
rect 36138 76294 36234 76350
rect 36290 76294 36358 76350
rect 36414 76294 36482 76350
rect 36538 76294 36606 76350
rect 36662 76294 36758 76350
rect 36138 76226 36758 76294
rect 36138 76170 36234 76226
rect 36290 76170 36358 76226
rect 36414 76170 36482 76226
rect 36538 76170 36606 76226
rect 36662 76170 36758 76226
rect 36138 76102 36758 76170
rect 36138 76046 36234 76102
rect 36290 76046 36358 76102
rect 36414 76046 36482 76102
rect 36538 76046 36606 76102
rect 36662 76046 36758 76102
rect 36138 75978 36758 76046
rect 36138 75922 36234 75978
rect 36290 75922 36358 75978
rect 36414 75922 36482 75978
rect 36538 75922 36606 75978
rect 36662 75922 36758 75978
rect 31808 64350 32128 64384
rect 31808 64294 31878 64350
rect 31934 64294 32002 64350
rect 32058 64294 32128 64350
rect 31808 64226 32128 64294
rect 31808 64170 31878 64226
rect 31934 64170 32002 64226
rect 32058 64170 32128 64226
rect 31808 64102 32128 64170
rect 31808 64046 31878 64102
rect 31934 64046 32002 64102
rect 32058 64046 32128 64102
rect 31808 63978 32128 64046
rect 31808 63922 31878 63978
rect 31934 63922 32002 63978
rect 32058 63922 32128 63978
rect 31808 63888 32128 63922
rect 31052 60352 31108 60362
rect 27692 49552 27748 49562
rect 36138 58350 36758 75922
rect 36138 58294 36234 58350
rect 36290 58294 36358 58350
rect 36414 58294 36482 58350
rect 36538 58294 36606 58350
rect 36662 58294 36758 58350
rect 36138 58226 36758 58294
rect 36138 58170 36234 58226
rect 36290 58170 36358 58226
rect 36414 58170 36482 58226
rect 36538 58170 36606 58226
rect 36662 58170 36758 58226
rect 36138 58102 36758 58170
rect 36138 58046 36234 58102
rect 36290 58046 36358 58102
rect 36414 58046 36482 58102
rect 36538 58046 36606 58102
rect 36662 58046 36758 58102
rect 36138 57978 36758 58046
rect 36138 57922 36234 57978
rect 36290 57922 36358 57978
rect 36414 57922 36482 57978
rect 36538 57922 36606 57978
rect 36662 57922 36758 57978
rect 19292 48652 19348 48662
rect 12684 48290 12740 48300
rect 31808 46350 32128 46384
rect 31808 46294 31878 46350
rect 31934 46294 32002 46350
rect 32058 46294 32128 46350
rect 31808 46226 32128 46294
rect 31808 46170 31878 46226
rect 31934 46170 32002 46226
rect 32058 46170 32128 46226
rect 31808 46102 32128 46170
rect 31808 46046 31878 46102
rect 31934 46046 32002 46102
rect 32058 46046 32128 46102
rect 31808 45978 32128 46046
rect 31808 45922 31878 45978
rect 31934 45922 32002 45978
rect 32058 45922 32128 45978
rect 31808 45888 32128 45922
rect 16448 40350 16768 40384
rect 16448 40294 16518 40350
rect 16574 40294 16642 40350
rect 16698 40294 16768 40350
rect 16448 40226 16768 40294
rect 16448 40170 16518 40226
rect 16574 40170 16642 40226
rect 16698 40170 16768 40226
rect 16448 40102 16768 40170
rect 16448 40046 16518 40102
rect 16574 40046 16642 40102
rect 16698 40046 16768 40102
rect 16448 39978 16768 40046
rect 16448 39922 16518 39978
rect 16574 39922 16642 39978
rect 16698 39922 16768 39978
rect 16448 39888 16768 39922
rect 36138 40350 36758 57922
rect 36138 40294 36234 40350
rect 36290 40294 36358 40350
rect 36414 40294 36482 40350
rect 36538 40294 36606 40350
rect 36662 40294 36758 40350
rect 36138 40226 36758 40294
rect 36138 40170 36234 40226
rect 36290 40170 36358 40226
rect 36414 40170 36482 40226
rect 36538 40170 36606 40226
rect 36662 40170 36758 40226
rect 36138 40102 36758 40170
rect 36138 40046 36234 40102
rect 36290 40046 36358 40102
rect 36414 40046 36482 40102
rect 36538 40046 36606 40102
rect 36662 40046 36758 40102
rect 36138 39978 36758 40046
rect 36138 39922 36234 39978
rect 36290 39922 36358 39978
rect 36414 39922 36482 39978
rect 36538 39922 36606 39978
rect 36662 39922 36758 39978
rect 12012 31892 12180 31948
rect 12012 26852 12068 31892
rect 31808 28350 32128 28384
rect 31808 28294 31878 28350
rect 31934 28294 32002 28350
rect 32058 28294 32128 28350
rect 31808 28226 32128 28294
rect 31808 28170 31878 28226
rect 31934 28170 32002 28226
rect 32058 28170 32128 28226
rect 31808 28102 32128 28170
rect 31808 28046 31878 28102
rect 31934 28046 32002 28102
rect 32058 28046 32128 28102
rect 31808 27978 32128 28046
rect 31808 27922 31878 27978
rect 31934 27922 32002 27978
rect 32058 27922 32128 27978
rect 31808 27888 32128 27922
rect 12012 26786 12068 26796
rect 11900 26522 12068 26578
rect 12012 23268 12068 26522
rect 12012 23202 12068 23212
rect 16448 22350 16768 22384
rect 16448 22294 16518 22350
rect 16574 22294 16642 22350
rect 16698 22294 16768 22350
rect 16448 22226 16768 22294
rect 16448 22170 16518 22226
rect 16574 22170 16642 22226
rect 16698 22170 16768 22226
rect 16448 22102 16768 22170
rect 16448 22046 16518 22102
rect 16574 22046 16642 22102
rect 16698 22046 16768 22102
rect 16448 21978 16768 22046
rect 16448 21922 16518 21978
rect 16574 21922 16642 21978
rect 16698 21922 16768 21978
rect 16448 21888 16768 21922
rect 36138 22350 36758 39922
rect 36138 22294 36234 22350
rect 36290 22294 36358 22350
rect 36414 22294 36482 22350
rect 36538 22294 36606 22350
rect 36662 22294 36758 22350
rect 36138 22226 36758 22294
rect 36138 22170 36234 22226
rect 36290 22170 36358 22226
rect 36414 22170 36482 22226
rect 36538 22170 36606 22226
rect 36662 22170 36758 22226
rect 36138 22102 36758 22170
rect 36138 22046 36234 22102
rect 36290 22046 36358 22102
rect 36414 22046 36482 22102
rect 36538 22046 36606 22102
rect 36662 22046 36758 22102
rect 36138 21978 36758 22046
rect 36138 21922 36234 21978
rect 36290 21922 36358 21978
rect 36414 21922 36482 21978
rect 36538 21922 36606 21978
rect 36662 21922 36758 21978
rect 11004 18722 11060 18732
rect 9138 10294 9234 10350
rect 9290 10294 9358 10350
rect 9414 10294 9482 10350
rect 9538 10294 9606 10350
rect 9662 10294 9758 10350
rect 9138 10226 9758 10294
rect 9138 10170 9234 10226
rect 9290 10170 9358 10226
rect 9414 10170 9482 10226
rect 9538 10170 9606 10226
rect 9662 10170 9758 10226
rect 9138 10102 9758 10170
rect 9138 10046 9234 10102
rect 9290 10046 9358 10102
rect 9414 10046 9482 10102
rect 9538 10046 9606 10102
rect 9662 10046 9758 10102
rect 9138 9978 9758 10046
rect 9138 9922 9234 9978
rect 9290 9922 9358 9978
rect 9414 9922 9482 9978
rect 9538 9922 9606 9978
rect 9662 9922 9758 9978
rect 5418 4294 5514 4350
rect 5570 4294 5638 4350
rect 5694 4294 5762 4350
rect 5818 4294 5886 4350
rect 5942 4294 6038 4350
rect 5418 4226 6038 4294
rect 5418 4170 5514 4226
rect 5570 4170 5638 4226
rect 5694 4170 5762 4226
rect 5818 4170 5886 4226
rect 5942 4170 6038 4226
rect 5418 4102 6038 4170
rect 5418 4046 5514 4102
rect 5570 4046 5638 4102
rect 5694 4046 5762 4102
rect 5818 4046 5886 4102
rect 5942 4046 6038 4102
rect 5418 3978 6038 4046
rect 5418 3922 5514 3978
rect 5570 3922 5638 3978
rect 5694 3922 5762 3978
rect 5818 3922 5886 3978
rect 5942 3922 6038 3978
rect 5418 -160 6038 3922
rect 5418 -216 5514 -160
rect 5570 -216 5638 -160
rect 5694 -216 5762 -160
rect 5818 -216 5886 -160
rect 5942 -216 6038 -160
rect 5418 -284 6038 -216
rect 5418 -340 5514 -284
rect 5570 -340 5638 -284
rect 5694 -340 5762 -284
rect 5818 -340 5886 -284
rect 5942 -340 6038 -284
rect 5418 -408 6038 -340
rect 5418 -464 5514 -408
rect 5570 -464 5638 -408
rect 5694 -464 5762 -408
rect 5818 -464 5886 -408
rect 5942 -464 6038 -408
rect 5418 -532 6038 -464
rect 5418 -588 5514 -532
rect 5570 -588 5638 -532
rect 5694 -588 5762 -532
rect 5818 -588 5886 -532
rect 5942 -588 6038 -532
rect -1916 -1176 -1820 -1120
rect -1764 -1176 -1696 -1120
rect -1640 -1176 -1572 -1120
rect -1516 -1176 -1448 -1120
rect -1392 -1176 -1296 -1120
rect -1916 -1244 -1296 -1176
rect -1916 -1300 -1820 -1244
rect -1764 -1300 -1696 -1244
rect -1640 -1300 -1572 -1244
rect -1516 -1300 -1448 -1244
rect -1392 -1300 -1296 -1244
rect -1916 -1368 -1296 -1300
rect -1916 -1424 -1820 -1368
rect -1764 -1424 -1696 -1368
rect -1640 -1424 -1572 -1368
rect -1516 -1424 -1448 -1368
rect -1392 -1424 -1296 -1368
rect -1916 -1492 -1296 -1424
rect -1916 -1548 -1820 -1492
rect -1764 -1548 -1696 -1492
rect -1640 -1548 -1572 -1492
rect -1516 -1548 -1448 -1492
rect -1392 -1548 -1296 -1492
rect -1916 -1644 -1296 -1548
rect 5418 -1644 6038 -588
rect 9138 -1120 9758 9922
rect 31808 10350 32128 10384
rect 31808 10294 31878 10350
rect 31934 10294 32002 10350
rect 32058 10294 32128 10350
rect 31808 10226 32128 10294
rect 31808 10170 31878 10226
rect 31934 10170 32002 10226
rect 32058 10170 32128 10226
rect 31808 10102 32128 10170
rect 31808 10046 31878 10102
rect 31934 10046 32002 10102
rect 32058 10046 32128 10102
rect 31808 9978 32128 10046
rect 31808 9922 31878 9978
rect 31934 9922 32002 9978
rect 32058 9922 32128 9978
rect 31808 9888 32128 9922
rect 36138 4350 36758 21922
rect 36138 4294 36234 4350
rect 36290 4294 36358 4350
rect 36414 4294 36482 4350
rect 36538 4294 36606 4350
rect 36662 4294 36758 4350
rect 36138 4226 36758 4294
rect 36138 4170 36234 4226
rect 36290 4170 36358 4226
rect 36414 4170 36482 4226
rect 36538 4170 36606 4226
rect 36662 4170 36758 4226
rect 36138 4102 36758 4170
rect 36138 4046 36234 4102
rect 36290 4046 36358 4102
rect 36414 4046 36482 4102
rect 36538 4046 36606 4102
rect 36662 4046 36758 4102
rect 36138 3978 36758 4046
rect 36138 3922 36234 3978
rect 36290 3922 36358 3978
rect 36414 3922 36482 3978
rect 36538 3922 36606 3978
rect 36662 3922 36758 3978
rect 31948 1428 32004 1438
rect 31948 838 32004 1372
rect 31892 782 32004 838
rect 31892 756 31948 782
rect 31892 690 31948 700
rect 9138 -1176 9234 -1120
rect 9290 -1176 9358 -1120
rect 9414 -1176 9482 -1120
rect 9538 -1176 9606 -1120
rect 9662 -1176 9758 -1120
rect 9138 -1244 9758 -1176
rect 9138 -1300 9234 -1244
rect 9290 -1300 9358 -1244
rect 9414 -1300 9482 -1244
rect 9538 -1300 9606 -1244
rect 9662 -1300 9758 -1244
rect 9138 -1368 9758 -1300
rect 9138 -1424 9234 -1368
rect 9290 -1424 9358 -1368
rect 9414 -1424 9482 -1368
rect 9538 -1424 9606 -1368
rect 9662 -1424 9758 -1368
rect 9138 -1492 9758 -1424
rect 9138 -1548 9234 -1492
rect 9290 -1548 9358 -1492
rect 9414 -1548 9482 -1492
rect 9538 -1548 9606 -1492
rect 9662 -1548 9758 -1492
rect 9138 -1644 9758 -1548
rect 36138 -160 36758 3922
rect 36138 -216 36234 -160
rect 36290 -216 36358 -160
rect 36414 -216 36482 -160
rect 36538 -216 36606 -160
rect 36662 -216 36758 -160
rect 36138 -284 36758 -216
rect 36138 -340 36234 -284
rect 36290 -340 36358 -284
rect 36414 -340 36482 -284
rect 36538 -340 36606 -284
rect 36662 -340 36758 -284
rect 36138 -408 36758 -340
rect 36138 -464 36234 -408
rect 36290 -464 36358 -408
rect 36414 -464 36482 -408
rect 36538 -464 36606 -408
rect 36662 -464 36758 -408
rect 36138 -532 36758 -464
rect 36138 -588 36234 -532
rect 36290 -588 36358 -532
rect 36414 -588 36482 -532
rect 36538 -588 36606 -532
rect 36662 -588 36758 -532
rect 36138 -1644 36758 -588
rect 39858 598172 40478 598268
rect 39858 598116 39954 598172
rect 40010 598116 40078 598172
rect 40134 598116 40202 598172
rect 40258 598116 40326 598172
rect 40382 598116 40478 598172
rect 39858 598048 40478 598116
rect 39858 597992 39954 598048
rect 40010 597992 40078 598048
rect 40134 597992 40202 598048
rect 40258 597992 40326 598048
rect 40382 597992 40478 598048
rect 39858 597924 40478 597992
rect 39858 597868 39954 597924
rect 40010 597868 40078 597924
rect 40134 597868 40202 597924
rect 40258 597868 40326 597924
rect 40382 597868 40478 597924
rect 39858 597800 40478 597868
rect 39858 597744 39954 597800
rect 40010 597744 40078 597800
rect 40134 597744 40202 597800
rect 40258 597744 40326 597800
rect 40382 597744 40478 597800
rect 39858 586350 40478 597744
rect 39858 586294 39954 586350
rect 40010 586294 40078 586350
rect 40134 586294 40202 586350
rect 40258 586294 40326 586350
rect 40382 586294 40478 586350
rect 39858 586226 40478 586294
rect 39858 586170 39954 586226
rect 40010 586170 40078 586226
rect 40134 586170 40202 586226
rect 40258 586170 40326 586226
rect 40382 586170 40478 586226
rect 39858 586102 40478 586170
rect 39858 586046 39954 586102
rect 40010 586046 40078 586102
rect 40134 586046 40202 586102
rect 40258 586046 40326 586102
rect 40382 586046 40478 586102
rect 39858 585978 40478 586046
rect 39858 585922 39954 585978
rect 40010 585922 40078 585978
rect 40134 585922 40202 585978
rect 40258 585922 40326 585978
rect 40382 585922 40478 585978
rect 39858 568350 40478 585922
rect 39858 568294 39954 568350
rect 40010 568294 40078 568350
rect 40134 568294 40202 568350
rect 40258 568294 40326 568350
rect 40382 568294 40478 568350
rect 39858 568226 40478 568294
rect 39858 568170 39954 568226
rect 40010 568170 40078 568226
rect 40134 568170 40202 568226
rect 40258 568170 40326 568226
rect 40382 568170 40478 568226
rect 39858 568102 40478 568170
rect 39858 568046 39954 568102
rect 40010 568046 40078 568102
rect 40134 568046 40202 568102
rect 40258 568046 40326 568102
rect 40382 568046 40478 568102
rect 39858 567978 40478 568046
rect 39858 567922 39954 567978
rect 40010 567922 40078 567978
rect 40134 567922 40202 567978
rect 40258 567922 40326 567978
rect 40382 567922 40478 567978
rect 39858 550350 40478 567922
rect 39858 550294 39954 550350
rect 40010 550294 40078 550350
rect 40134 550294 40202 550350
rect 40258 550294 40326 550350
rect 40382 550294 40478 550350
rect 39858 550226 40478 550294
rect 39858 550170 39954 550226
rect 40010 550170 40078 550226
rect 40134 550170 40202 550226
rect 40258 550170 40326 550226
rect 40382 550170 40478 550226
rect 39858 550102 40478 550170
rect 39858 550046 39954 550102
rect 40010 550046 40078 550102
rect 40134 550046 40202 550102
rect 40258 550046 40326 550102
rect 40382 550046 40478 550102
rect 39858 549978 40478 550046
rect 39858 549922 39954 549978
rect 40010 549922 40078 549978
rect 40134 549922 40202 549978
rect 40258 549922 40326 549978
rect 40382 549922 40478 549978
rect 39858 532350 40478 549922
rect 39858 532294 39954 532350
rect 40010 532294 40078 532350
rect 40134 532294 40202 532350
rect 40258 532294 40326 532350
rect 40382 532294 40478 532350
rect 39858 532226 40478 532294
rect 39858 532170 39954 532226
rect 40010 532170 40078 532226
rect 40134 532170 40202 532226
rect 40258 532170 40326 532226
rect 40382 532170 40478 532226
rect 39858 532102 40478 532170
rect 39858 532046 39954 532102
rect 40010 532046 40078 532102
rect 40134 532046 40202 532102
rect 40258 532046 40326 532102
rect 40382 532046 40478 532102
rect 39858 531978 40478 532046
rect 39858 531922 39954 531978
rect 40010 531922 40078 531978
rect 40134 531922 40202 531978
rect 40258 531922 40326 531978
rect 40382 531922 40478 531978
rect 39858 514350 40478 531922
rect 39858 514294 39954 514350
rect 40010 514294 40078 514350
rect 40134 514294 40202 514350
rect 40258 514294 40326 514350
rect 40382 514294 40478 514350
rect 39858 514226 40478 514294
rect 39858 514170 39954 514226
rect 40010 514170 40078 514226
rect 40134 514170 40202 514226
rect 40258 514170 40326 514226
rect 40382 514170 40478 514226
rect 39858 514102 40478 514170
rect 39858 514046 39954 514102
rect 40010 514046 40078 514102
rect 40134 514046 40202 514102
rect 40258 514046 40326 514102
rect 40382 514046 40478 514102
rect 39858 513978 40478 514046
rect 39858 513922 39954 513978
rect 40010 513922 40078 513978
rect 40134 513922 40202 513978
rect 40258 513922 40326 513978
rect 40382 513922 40478 513978
rect 39858 496350 40478 513922
rect 39858 496294 39954 496350
rect 40010 496294 40078 496350
rect 40134 496294 40202 496350
rect 40258 496294 40326 496350
rect 40382 496294 40478 496350
rect 39858 496226 40478 496294
rect 39858 496170 39954 496226
rect 40010 496170 40078 496226
rect 40134 496170 40202 496226
rect 40258 496170 40326 496226
rect 40382 496170 40478 496226
rect 39858 496102 40478 496170
rect 39858 496046 39954 496102
rect 40010 496046 40078 496102
rect 40134 496046 40202 496102
rect 40258 496046 40326 496102
rect 40382 496046 40478 496102
rect 39858 495978 40478 496046
rect 39858 495922 39954 495978
rect 40010 495922 40078 495978
rect 40134 495922 40202 495978
rect 40258 495922 40326 495978
rect 40382 495922 40478 495978
rect 39858 478350 40478 495922
rect 39858 478294 39954 478350
rect 40010 478294 40078 478350
rect 40134 478294 40202 478350
rect 40258 478294 40326 478350
rect 40382 478294 40478 478350
rect 39858 478226 40478 478294
rect 39858 478170 39954 478226
rect 40010 478170 40078 478226
rect 40134 478170 40202 478226
rect 40258 478170 40326 478226
rect 40382 478170 40478 478226
rect 39858 478102 40478 478170
rect 39858 478046 39954 478102
rect 40010 478046 40078 478102
rect 40134 478046 40202 478102
rect 40258 478046 40326 478102
rect 40382 478046 40478 478102
rect 39858 477978 40478 478046
rect 39858 477922 39954 477978
rect 40010 477922 40078 477978
rect 40134 477922 40202 477978
rect 40258 477922 40326 477978
rect 40382 477922 40478 477978
rect 39858 460350 40478 477922
rect 39858 460294 39954 460350
rect 40010 460294 40078 460350
rect 40134 460294 40202 460350
rect 40258 460294 40326 460350
rect 40382 460294 40478 460350
rect 39858 460226 40478 460294
rect 39858 460170 39954 460226
rect 40010 460170 40078 460226
rect 40134 460170 40202 460226
rect 40258 460170 40326 460226
rect 40382 460170 40478 460226
rect 39858 460102 40478 460170
rect 39858 460046 39954 460102
rect 40010 460046 40078 460102
rect 40134 460046 40202 460102
rect 40258 460046 40326 460102
rect 40382 460046 40478 460102
rect 39858 459978 40478 460046
rect 39858 459922 39954 459978
rect 40010 459922 40078 459978
rect 40134 459922 40202 459978
rect 40258 459922 40326 459978
rect 40382 459922 40478 459978
rect 39858 442350 40478 459922
rect 39858 442294 39954 442350
rect 40010 442294 40078 442350
rect 40134 442294 40202 442350
rect 40258 442294 40326 442350
rect 40382 442294 40478 442350
rect 39858 442226 40478 442294
rect 39858 442170 39954 442226
rect 40010 442170 40078 442226
rect 40134 442170 40202 442226
rect 40258 442170 40326 442226
rect 40382 442170 40478 442226
rect 39858 442102 40478 442170
rect 39858 442046 39954 442102
rect 40010 442046 40078 442102
rect 40134 442046 40202 442102
rect 40258 442046 40326 442102
rect 40382 442046 40478 442102
rect 39858 441978 40478 442046
rect 39858 441922 39954 441978
rect 40010 441922 40078 441978
rect 40134 441922 40202 441978
rect 40258 441922 40326 441978
rect 40382 441922 40478 441978
rect 39858 424350 40478 441922
rect 39858 424294 39954 424350
rect 40010 424294 40078 424350
rect 40134 424294 40202 424350
rect 40258 424294 40326 424350
rect 40382 424294 40478 424350
rect 39858 424226 40478 424294
rect 39858 424170 39954 424226
rect 40010 424170 40078 424226
rect 40134 424170 40202 424226
rect 40258 424170 40326 424226
rect 40382 424170 40478 424226
rect 39858 424102 40478 424170
rect 39858 424046 39954 424102
rect 40010 424046 40078 424102
rect 40134 424046 40202 424102
rect 40258 424046 40326 424102
rect 40382 424046 40478 424102
rect 39858 423978 40478 424046
rect 39858 423922 39954 423978
rect 40010 423922 40078 423978
rect 40134 423922 40202 423978
rect 40258 423922 40326 423978
rect 40382 423922 40478 423978
rect 39858 406350 40478 423922
rect 39858 406294 39954 406350
rect 40010 406294 40078 406350
rect 40134 406294 40202 406350
rect 40258 406294 40326 406350
rect 40382 406294 40478 406350
rect 39858 406226 40478 406294
rect 39858 406170 39954 406226
rect 40010 406170 40078 406226
rect 40134 406170 40202 406226
rect 40258 406170 40326 406226
rect 40382 406170 40478 406226
rect 39858 406102 40478 406170
rect 39858 406046 39954 406102
rect 40010 406046 40078 406102
rect 40134 406046 40202 406102
rect 40258 406046 40326 406102
rect 40382 406046 40478 406102
rect 39858 405978 40478 406046
rect 39858 405922 39954 405978
rect 40010 405922 40078 405978
rect 40134 405922 40202 405978
rect 40258 405922 40326 405978
rect 40382 405922 40478 405978
rect 39858 388350 40478 405922
rect 39858 388294 39954 388350
rect 40010 388294 40078 388350
rect 40134 388294 40202 388350
rect 40258 388294 40326 388350
rect 40382 388294 40478 388350
rect 39858 388226 40478 388294
rect 39858 388170 39954 388226
rect 40010 388170 40078 388226
rect 40134 388170 40202 388226
rect 40258 388170 40326 388226
rect 40382 388170 40478 388226
rect 39858 388102 40478 388170
rect 39858 388046 39954 388102
rect 40010 388046 40078 388102
rect 40134 388046 40202 388102
rect 40258 388046 40326 388102
rect 40382 388046 40478 388102
rect 39858 387978 40478 388046
rect 39858 387922 39954 387978
rect 40010 387922 40078 387978
rect 40134 387922 40202 387978
rect 40258 387922 40326 387978
rect 40382 387922 40478 387978
rect 39858 370350 40478 387922
rect 39858 370294 39954 370350
rect 40010 370294 40078 370350
rect 40134 370294 40202 370350
rect 40258 370294 40326 370350
rect 40382 370294 40478 370350
rect 39858 370226 40478 370294
rect 39858 370170 39954 370226
rect 40010 370170 40078 370226
rect 40134 370170 40202 370226
rect 40258 370170 40326 370226
rect 40382 370170 40478 370226
rect 39858 370102 40478 370170
rect 39858 370046 39954 370102
rect 40010 370046 40078 370102
rect 40134 370046 40202 370102
rect 40258 370046 40326 370102
rect 40382 370046 40478 370102
rect 39858 369978 40478 370046
rect 39858 369922 39954 369978
rect 40010 369922 40078 369978
rect 40134 369922 40202 369978
rect 40258 369922 40326 369978
rect 40382 369922 40478 369978
rect 39858 352350 40478 369922
rect 39858 352294 39954 352350
rect 40010 352294 40078 352350
rect 40134 352294 40202 352350
rect 40258 352294 40326 352350
rect 40382 352294 40478 352350
rect 39858 352226 40478 352294
rect 39858 352170 39954 352226
rect 40010 352170 40078 352226
rect 40134 352170 40202 352226
rect 40258 352170 40326 352226
rect 40382 352170 40478 352226
rect 39858 352102 40478 352170
rect 39858 352046 39954 352102
rect 40010 352046 40078 352102
rect 40134 352046 40202 352102
rect 40258 352046 40326 352102
rect 40382 352046 40478 352102
rect 39858 351978 40478 352046
rect 39858 351922 39954 351978
rect 40010 351922 40078 351978
rect 40134 351922 40202 351978
rect 40258 351922 40326 351978
rect 40382 351922 40478 351978
rect 39858 334350 40478 351922
rect 39858 334294 39954 334350
rect 40010 334294 40078 334350
rect 40134 334294 40202 334350
rect 40258 334294 40326 334350
rect 40382 334294 40478 334350
rect 39858 334226 40478 334294
rect 39858 334170 39954 334226
rect 40010 334170 40078 334226
rect 40134 334170 40202 334226
rect 40258 334170 40326 334226
rect 40382 334170 40478 334226
rect 39858 334102 40478 334170
rect 39858 334046 39954 334102
rect 40010 334046 40078 334102
rect 40134 334046 40202 334102
rect 40258 334046 40326 334102
rect 40382 334046 40478 334102
rect 39858 333978 40478 334046
rect 39858 333922 39954 333978
rect 40010 333922 40078 333978
rect 40134 333922 40202 333978
rect 40258 333922 40326 333978
rect 40382 333922 40478 333978
rect 39858 316350 40478 333922
rect 66858 597212 67478 598268
rect 66858 597156 66954 597212
rect 67010 597156 67078 597212
rect 67134 597156 67202 597212
rect 67258 597156 67326 597212
rect 67382 597156 67478 597212
rect 66858 597088 67478 597156
rect 66858 597032 66954 597088
rect 67010 597032 67078 597088
rect 67134 597032 67202 597088
rect 67258 597032 67326 597088
rect 67382 597032 67478 597088
rect 66858 596964 67478 597032
rect 66858 596908 66954 596964
rect 67010 596908 67078 596964
rect 67134 596908 67202 596964
rect 67258 596908 67326 596964
rect 67382 596908 67478 596964
rect 66858 596840 67478 596908
rect 66858 596784 66954 596840
rect 67010 596784 67078 596840
rect 67134 596784 67202 596840
rect 67258 596784 67326 596840
rect 67382 596784 67478 596840
rect 66858 580350 67478 596784
rect 66858 580294 66954 580350
rect 67010 580294 67078 580350
rect 67134 580294 67202 580350
rect 67258 580294 67326 580350
rect 67382 580294 67478 580350
rect 66858 580226 67478 580294
rect 66858 580170 66954 580226
rect 67010 580170 67078 580226
rect 67134 580170 67202 580226
rect 67258 580170 67326 580226
rect 67382 580170 67478 580226
rect 66858 580102 67478 580170
rect 66858 580046 66954 580102
rect 67010 580046 67078 580102
rect 67134 580046 67202 580102
rect 67258 580046 67326 580102
rect 67382 580046 67478 580102
rect 66858 579978 67478 580046
rect 66858 579922 66954 579978
rect 67010 579922 67078 579978
rect 67134 579922 67202 579978
rect 67258 579922 67326 579978
rect 67382 579922 67478 579978
rect 66858 562350 67478 579922
rect 66858 562294 66954 562350
rect 67010 562294 67078 562350
rect 67134 562294 67202 562350
rect 67258 562294 67326 562350
rect 67382 562294 67478 562350
rect 66858 562226 67478 562294
rect 66858 562170 66954 562226
rect 67010 562170 67078 562226
rect 67134 562170 67202 562226
rect 67258 562170 67326 562226
rect 67382 562170 67478 562226
rect 66858 562102 67478 562170
rect 66858 562046 66954 562102
rect 67010 562046 67078 562102
rect 67134 562046 67202 562102
rect 67258 562046 67326 562102
rect 67382 562046 67478 562102
rect 66858 561978 67478 562046
rect 66858 561922 66954 561978
rect 67010 561922 67078 561978
rect 67134 561922 67202 561978
rect 67258 561922 67326 561978
rect 67382 561922 67478 561978
rect 66858 544350 67478 561922
rect 66858 544294 66954 544350
rect 67010 544294 67078 544350
rect 67134 544294 67202 544350
rect 67258 544294 67326 544350
rect 67382 544294 67478 544350
rect 66858 544226 67478 544294
rect 66858 544170 66954 544226
rect 67010 544170 67078 544226
rect 67134 544170 67202 544226
rect 67258 544170 67326 544226
rect 67382 544170 67478 544226
rect 66858 544102 67478 544170
rect 66858 544046 66954 544102
rect 67010 544046 67078 544102
rect 67134 544046 67202 544102
rect 67258 544046 67326 544102
rect 67382 544046 67478 544102
rect 66858 543978 67478 544046
rect 66858 543922 66954 543978
rect 67010 543922 67078 543978
rect 67134 543922 67202 543978
rect 67258 543922 67326 543978
rect 67382 543922 67478 543978
rect 66858 526350 67478 543922
rect 66858 526294 66954 526350
rect 67010 526294 67078 526350
rect 67134 526294 67202 526350
rect 67258 526294 67326 526350
rect 67382 526294 67478 526350
rect 66858 526226 67478 526294
rect 66858 526170 66954 526226
rect 67010 526170 67078 526226
rect 67134 526170 67202 526226
rect 67258 526170 67326 526226
rect 67382 526170 67478 526226
rect 66858 526102 67478 526170
rect 66858 526046 66954 526102
rect 67010 526046 67078 526102
rect 67134 526046 67202 526102
rect 67258 526046 67326 526102
rect 67382 526046 67478 526102
rect 66858 525978 67478 526046
rect 66858 525922 66954 525978
rect 67010 525922 67078 525978
rect 67134 525922 67202 525978
rect 67258 525922 67326 525978
rect 67382 525922 67478 525978
rect 66858 508350 67478 525922
rect 66858 508294 66954 508350
rect 67010 508294 67078 508350
rect 67134 508294 67202 508350
rect 67258 508294 67326 508350
rect 67382 508294 67478 508350
rect 66858 508226 67478 508294
rect 66858 508170 66954 508226
rect 67010 508170 67078 508226
rect 67134 508170 67202 508226
rect 67258 508170 67326 508226
rect 67382 508170 67478 508226
rect 66858 508102 67478 508170
rect 66858 508046 66954 508102
rect 67010 508046 67078 508102
rect 67134 508046 67202 508102
rect 67258 508046 67326 508102
rect 67382 508046 67478 508102
rect 66858 507978 67478 508046
rect 66858 507922 66954 507978
rect 67010 507922 67078 507978
rect 67134 507922 67202 507978
rect 67258 507922 67326 507978
rect 67382 507922 67478 507978
rect 66858 490350 67478 507922
rect 66858 490294 66954 490350
rect 67010 490294 67078 490350
rect 67134 490294 67202 490350
rect 67258 490294 67326 490350
rect 67382 490294 67478 490350
rect 66858 490226 67478 490294
rect 66858 490170 66954 490226
rect 67010 490170 67078 490226
rect 67134 490170 67202 490226
rect 67258 490170 67326 490226
rect 67382 490170 67478 490226
rect 66858 490102 67478 490170
rect 66858 490046 66954 490102
rect 67010 490046 67078 490102
rect 67134 490046 67202 490102
rect 67258 490046 67326 490102
rect 67382 490046 67478 490102
rect 66858 489978 67478 490046
rect 66858 489922 66954 489978
rect 67010 489922 67078 489978
rect 67134 489922 67202 489978
rect 67258 489922 67326 489978
rect 67382 489922 67478 489978
rect 66858 472350 67478 489922
rect 66858 472294 66954 472350
rect 67010 472294 67078 472350
rect 67134 472294 67202 472350
rect 67258 472294 67326 472350
rect 67382 472294 67478 472350
rect 66858 472226 67478 472294
rect 66858 472170 66954 472226
rect 67010 472170 67078 472226
rect 67134 472170 67202 472226
rect 67258 472170 67326 472226
rect 67382 472170 67478 472226
rect 66858 472102 67478 472170
rect 66858 472046 66954 472102
rect 67010 472046 67078 472102
rect 67134 472046 67202 472102
rect 67258 472046 67326 472102
rect 67382 472046 67478 472102
rect 66858 471978 67478 472046
rect 66858 471922 66954 471978
rect 67010 471922 67078 471978
rect 67134 471922 67202 471978
rect 67258 471922 67326 471978
rect 67382 471922 67478 471978
rect 66858 454350 67478 471922
rect 66858 454294 66954 454350
rect 67010 454294 67078 454350
rect 67134 454294 67202 454350
rect 67258 454294 67326 454350
rect 67382 454294 67478 454350
rect 66858 454226 67478 454294
rect 66858 454170 66954 454226
rect 67010 454170 67078 454226
rect 67134 454170 67202 454226
rect 67258 454170 67326 454226
rect 67382 454170 67478 454226
rect 66858 454102 67478 454170
rect 66858 454046 66954 454102
rect 67010 454046 67078 454102
rect 67134 454046 67202 454102
rect 67258 454046 67326 454102
rect 67382 454046 67478 454102
rect 66858 453978 67478 454046
rect 66858 453922 66954 453978
rect 67010 453922 67078 453978
rect 67134 453922 67202 453978
rect 67258 453922 67326 453978
rect 67382 453922 67478 453978
rect 66858 436350 67478 453922
rect 66858 436294 66954 436350
rect 67010 436294 67078 436350
rect 67134 436294 67202 436350
rect 67258 436294 67326 436350
rect 67382 436294 67478 436350
rect 66858 436226 67478 436294
rect 66858 436170 66954 436226
rect 67010 436170 67078 436226
rect 67134 436170 67202 436226
rect 67258 436170 67326 436226
rect 67382 436170 67478 436226
rect 66858 436102 67478 436170
rect 66858 436046 66954 436102
rect 67010 436046 67078 436102
rect 67134 436046 67202 436102
rect 67258 436046 67326 436102
rect 67382 436046 67478 436102
rect 66858 435978 67478 436046
rect 66858 435922 66954 435978
rect 67010 435922 67078 435978
rect 67134 435922 67202 435978
rect 67258 435922 67326 435978
rect 67382 435922 67478 435978
rect 66858 418350 67478 435922
rect 66858 418294 66954 418350
rect 67010 418294 67078 418350
rect 67134 418294 67202 418350
rect 67258 418294 67326 418350
rect 67382 418294 67478 418350
rect 66858 418226 67478 418294
rect 66858 418170 66954 418226
rect 67010 418170 67078 418226
rect 67134 418170 67202 418226
rect 67258 418170 67326 418226
rect 67382 418170 67478 418226
rect 66858 418102 67478 418170
rect 66858 418046 66954 418102
rect 67010 418046 67078 418102
rect 67134 418046 67202 418102
rect 67258 418046 67326 418102
rect 67382 418046 67478 418102
rect 66858 417978 67478 418046
rect 66858 417922 66954 417978
rect 67010 417922 67078 417978
rect 67134 417922 67202 417978
rect 67258 417922 67326 417978
rect 67382 417922 67478 417978
rect 66858 400350 67478 417922
rect 66858 400294 66954 400350
rect 67010 400294 67078 400350
rect 67134 400294 67202 400350
rect 67258 400294 67326 400350
rect 67382 400294 67478 400350
rect 66858 400226 67478 400294
rect 66858 400170 66954 400226
rect 67010 400170 67078 400226
rect 67134 400170 67202 400226
rect 67258 400170 67326 400226
rect 67382 400170 67478 400226
rect 66858 400102 67478 400170
rect 66858 400046 66954 400102
rect 67010 400046 67078 400102
rect 67134 400046 67202 400102
rect 67258 400046 67326 400102
rect 67382 400046 67478 400102
rect 66858 399978 67478 400046
rect 66858 399922 66954 399978
rect 67010 399922 67078 399978
rect 67134 399922 67202 399978
rect 67258 399922 67326 399978
rect 67382 399922 67478 399978
rect 66858 382350 67478 399922
rect 66858 382294 66954 382350
rect 67010 382294 67078 382350
rect 67134 382294 67202 382350
rect 67258 382294 67326 382350
rect 67382 382294 67478 382350
rect 66858 382226 67478 382294
rect 66858 382170 66954 382226
rect 67010 382170 67078 382226
rect 67134 382170 67202 382226
rect 67258 382170 67326 382226
rect 67382 382170 67478 382226
rect 66858 382102 67478 382170
rect 66858 382046 66954 382102
rect 67010 382046 67078 382102
rect 67134 382046 67202 382102
rect 67258 382046 67326 382102
rect 67382 382046 67478 382102
rect 66858 381978 67478 382046
rect 66858 381922 66954 381978
rect 67010 381922 67078 381978
rect 67134 381922 67202 381978
rect 67258 381922 67326 381978
rect 67382 381922 67478 381978
rect 66858 364350 67478 381922
rect 66858 364294 66954 364350
rect 67010 364294 67078 364350
rect 67134 364294 67202 364350
rect 67258 364294 67326 364350
rect 67382 364294 67478 364350
rect 66858 364226 67478 364294
rect 66858 364170 66954 364226
rect 67010 364170 67078 364226
rect 67134 364170 67202 364226
rect 67258 364170 67326 364226
rect 67382 364170 67478 364226
rect 66858 364102 67478 364170
rect 66858 364046 66954 364102
rect 67010 364046 67078 364102
rect 67134 364046 67202 364102
rect 67258 364046 67326 364102
rect 67382 364046 67478 364102
rect 66858 363978 67478 364046
rect 66858 363922 66954 363978
rect 67010 363922 67078 363978
rect 67134 363922 67202 363978
rect 67258 363922 67326 363978
rect 67382 363922 67478 363978
rect 66858 346350 67478 363922
rect 66858 346294 66954 346350
rect 67010 346294 67078 346350
rect 67134 346294 67202 346350
rect 67258 346294 67326 346350
rect 67382 346294 67478 346350
rect 66858 346226 67478 346294
rect 66858 346170 66954 346226
rect 67010 346170 67078 346226
rect 67134 346170 67202 346226
rect 67258 346170 67326 346226
rect 67382 346170 67478 346226
rect 66858 346102 67478 346170
rect 66858 346046 66954 346102
rect 67010 346046 67078 346102
rect 67134 346046 67202 346102
rect 67258 346046 67326 346102
rect 67382 346046 67478 346102
rect 66858 345978 67478 346046
rect 66858 345922 66954 345978
rect 67010 345922 67078 345978
rect 67134 345922 67202 345978
rect 67258 345922 67326 345978
rect 67382 345922 67478 345978
rect 66858 328350 67478 345922
rect 66858 328294 66954 328350
rect 67010 328294 67078 328350
rect 67134 328294 67202 328350
rect 67258 328294 67326 328350
rect 67382 328294 67478 328350
rect 66858 328226 67478 328294
rect 66858 328170 66954 328226
rect 67010 328170 67078 328226
rect 67134 328170 67202 328226
rect 67258 328170 67326 328226
rect 67382 328170 67478 328226
rect 66858 328102 67478 328170
rect 66858 328046 66954 328102
rect 67010 328046 67078 328102
rect 67134 328046 67202 328102
rect 67258 328046 67326 328102
rect 67382 328046 67478 328102
rect 66858 327978 67478 328046
rect 66858 327922 66954 327978
rect 67010 327922 67078 327978
rect 67134 327922 67202 327978
rect 67258 327922 67326 327978
rect 67382 327922 67478 327978
rect 39858 316294 39954 316350
rect 40010 316294 40078 316350
rect 40134 316294 40202 316350
rect 40258 316294 40326 316350
rect 40382 316294 40478 316350
rect 39858 316226 40478 316294
rect 39858 316170 39954 316226
rect 40010 316170 40078 316226
rect 40134 316170 40202 316226
rect 40258 316170 40326 316226
rect 40382 316170 40478 316226
rect 39858 316102 40478 316170
rect 39858 316046 39954 316102
rect 40010 316046 40078 316102
rect 40134 316046 40202 316102
rect 40258 316046 40326 316102
rect 40382 316046 40478 316102
rect 39858 315978 40478 316046
rect 39858 315922 39954 315978
rect 40010 315922 40078 315978
rect 40134 315922 40202 315978
rect 40258 315922 40326 315978
rect 40382 315922 40478 315978
rect 39858 298350 40478 315922
rect 39858 298294 39954 298350
rect 40010 298294 40078 298350
rect 40134 298294 40202 298350
rect 40258 298294 40326 298350
rect 40382 298294 40478 298350
rect 39858 298226 40478 298294
rect 39858 298170 39954 298226
rect 40010 298170 40078 298226
rect 40134 298170 40202 298226
rect 40258 298170 40326 298226
rect 40382 298170 40478 298226
rect 39858 298102 40478 298170
rect 39858 298046 39954 298102
rect 40010 298046 40078 298102
rect 40134 298046 40202 298102
rect 40258 298046 40326 298102
rect 40382 298046 40478 298102
rect 39858 297978 40478 298046
rect 39858 297922 39954 297978
rect 40010 297922 40078 297978
rect 40134 297922 40202 297978
rect 40258 297922 40326 297978
rect 40382 297922 40478 297978
rect 39858 280350 40478 297922
rect 39858 280294 39954 280350
rect 40010 280294 40078 280350
rect 40134 280294 40202 280350
rect 40258 280294 40326 280350
rect 40382 280294 40478 280350
rect 39858 280226 40478 280294
rect 39858 280170 39954 280226
rect 40010 280170 40078 280226
rect 40134 280170 40202 280226
rect 40258 280170 40326 280226
rect 40382 280170 40478 280226
rect 39858 280102 40478 280170
rect 39858 280046 39954 280102
rect 40010 280046 40078 280102
rect 40134 280046 40202 280102
rect 40258 280046 40326 280102
rect 40382 280046 40478 280102
rect 39858 279978 40478 280046
rect 39858 279922 39954 279978
rect 40010 279922 40078 279978
rect 40134 279922 40202 279978
rect 40258 279922 40326 279978
rect 40382 279922 40478 279978
rect 39858 262350 40478 279922
rect 39858 262294 39954 262350
rect 40010 262294 40078 262350
rect 40134 262294 40202 262350
rect 40258 262294 40326 262350
rect 40382 262294 40478 262350
rect 39858 262226 40478 262294
rect 39858 262170 39954 262226
rect 40010 262170 40078 262226
rect 40134 262170 40202 262226
rect 40258 262170 40326 262226
rect 40382 262170 40478 262226
rect 39858 262102 40478 262170
rect 39858 262046 39954 262102
rect 40010 262046 40078 262102
rect 40134 262046 40202 262102
rect 40258 262046 40326 262102
rect 40382 262046 40478 262102
rect 39858 261978 40478 262046
rect 39858 261922 39954 261978
rect 40010 261922 40078 261978
rect 40134 261922 40202 261978
rect 40258 261922 40326 261978
rect 40382 261922 40478 261978
rect 39858 244350 40478 261922
rect 39858 244294 39954 244350
rect 40010 244294 40078 244350
rect 40134 244294 40202 244350
rect 40258 244294 40326 244350
rect 40382 244294 40478 244350
rect 39858 244226 40478 244294
rect 39858 244170 39954 244226
rect 40010 244170 40078 244226
rect 40134 244170 40202 244226
rect 40258 244170 40326 244226
rect 40382 244170 40478 244226
rect 39858 244102 40478 244170
rect 39858 244046 39954 244102
rect 40010 244046 40078 244102
rect 40134 244046 40202 244102
rect 40258 244046 40326 244102
rect 40382 244046 40478 244102
rect 39858 243978 40478 244046
rect 39858 243922 39954 243978
rect 40010 243922 40078 243978
rect 40134 243922 40202 243978
rect 40258 243922 40326 243978
rect 40382 243922 40478 243978
rect 39858 226350 40478 243922
rect 39858 226294 39954 226350
rect 40010 226294 40078 226350
rect 40134 226294 40202 226350
rect 40258 226294 40326 226350
rect 40382 226294 40478 226350
rect 39858 226226 40478 226294
rect 39858 226170 39954 226226
rect 40010 226170 40078 226226
rect 40134 226170 40202 226226
rect 40258 226170 40326 226226
rect 40382 226170 40478 226226
rect 39858 226102 40478 226170
rect 39858 226046 39954 226102
rect 40010 226046 40078 226102
rect 40134 226046 40202 226102
rect 40258 226046 40326 226102
rect 40382 226046 40478 226102
rect 39858 225978 40478 226046
rect 39858 225922 39954 225978
rect 40010 225922 40078 225978
rect 40134 225922 40202 225978
rect 40258 225922 40326 225978
rect 40382 225922 40478 225978
rect 39858 208350 40478 225922
rect 39858 208294 39954 208350
rect 40010 208294 40078 208350
rect 40134 208294 40202 208350
rect 40258 208294 40326 208350
rect 40382 208294 40478 208350
rect 39858 208226 40478 208294
rect 39858 208170 39954 208226
rect 40010 208170 40078 208226
rect 40134 208170 40202 208226
rect 40258 208170 40326 208226
rect 40382 208170 40478 208226
rect 39858 208102 40478 208170
rect 39858 208046 39954 208102
rect 40010 208046 40078 208102
rect 40134 208046 40202 208102
rect 40258 208046 40326 208102
rect 40382 208046 40478 208102
rect 39858 207978 40478 208046
rect 39858 207922 39954 207978
rect 40010 207922 40078 207978
rect 40134 207922 40202 207978
rect 40258 207922 40326 207978
rect 40382 207922 40478 207978
rect 39858 190350 40478 207922
rect 39858 190294 39954 190350
rect 40010 190294 40078 190350
rect 40134 190294 40202 190350
rect 40258 190294 40326 190350
rect 40382 190294 40478 190350
rect 39858 190226 40478 190294
rect 39858 190170 39954 190226
rect 40010 190170 40078 190226
rect 40134 190170 40202 190226
rect 40258 190170 40326 190226
rect 40382 190170 40478 190226
rect 39858 190102 40478 190170
rect 39858 190046 39954 190102
rect 40010 190046 40078 190102
rect 40134 190046 40202 190102
rect 40258 190046 40326 190102
rect 40382 190046 40478 190102
rect 39858 189978 40478 190046
rect 39858 189922 39954 189978
rect 40010 189922 40078 189978
rect 40134 189922 40202 189978
rect 40258 189922 40326 189978
rect 40382 189922 40478 189978
rect 39858 172350 40478 189922
rect 39858 172294 39954 172350
rect 40010 172294 40078 172350
rect 40134 172294 40202 172350
rect 40258 172294 40326 172350
rect 40382 172294 40478 172350
rect 39858 172226 40478 172294
rect 39858 172170 39954 172226
rect 40010 172170 40078 172226
rect 40134 172170 40202 172226
rect 40258 172170 40326 172226
rect 40382 172170 40478 172226
rect 39858 172102 40478 172170
rect 39858 172046 39954 172102
rect 40010 172046 40078 172102
rect 40134 172046 40202 172102
rect 40258 172046 40326 172102
rect 40382 172046 40478 172102
rect 39858 171978 40478 172046
rect 39858 171922 39954 171978
rect 40010 171922 40078 171978
rect 40134 171922 40202 171978
rect 40258 171922 40326 171978
rect 40382 171922 40478 171978
rect 39858 154350 40478 171922
rect 39858 154294 39954 154350
rect 40010 154294 40078 154350
rect 40134 154294 40202 154350
rect 40258 154294 40326 154350
rect 40382 154294 40478 154350
rect 39858 154226 40478 154294
rect 39858 154170 39954 154226
rect 40010 154170 40078 154226
rect 40134 154170 40202 154226
rect 40258 154170 40326 154226
rect 40382 154170 40478 154226
rect 39858 154102 40478 154170
rect 39858 154046 39954 154102
rect 40010 154046 40078 154102
rect 40134 154046 40202 154102
rect 40258 154046 40326 154102
rect 40382 154046 40478 154102
rect 39858 153978 40478 154046
rect 39858 153922 39954 153978
rect 40010 153922 40078 153978
rect 40134 153922 40202 153978
rect 40258 153922 40326 153978
rect 40382 153922 40478 153978
rect 39858 136350 40478 153922
rect 39858 136294 39954 136350
rect 40010 136294 40078 136350
rect 40134 136294 40202 136350
rect 40258 136294 40326 136350
rect 40382 136294 40478 136350
rect 39858 136226 40478 136294
rect 39858 136170 39954 136226
rect 40010 136170 40078 136226
rect 40134 136170 40202 136226
rect 40258 136170 40326 136226
rect 40382 136170 40478 136226
rect 39858 136102 40478 136170
rect 39858 136046 39954 136102
rect 40010 136046 40078 136102
rect 40134 136046 40202 136102
rect 40258 136046 40326 136102
rect 40382 136046 40478 136102
rect 39858 135978 40478 136046
rect 39858 135922 39954 135978
rect 40010 135922 40078 135978
rect 40134 135922 40202 135978
rect 40258 135922 40326 135978
rect 40382 135922 40478 135978
rect 39858 118350 40478 135922
rect 39858 118294 39954 118350
rect 40010 118294 40078 118350
rect 40134 118294 40202 118350
rect 40258 118294 40326 118350
rect 40382 118294 40478 118350
rect 39858 118226 40478 118294
rect 39858 118170 39954 118226
rect 40010 118170 40078 118226
rect 40134 118170 40202 118226
rect 40258 118170 40326 118226
rect 40382 118170 40478 118226
rect 39858 118102 40478 118170
rect 39858 118046 39954 118102
rect 40010 118046 40078 118102
rect 40134 118046 40202 118102
rect 40258 118046 40326 118102
rect 40382 118046 40478 118102
rect 39858 117978 40478 118046
rect 39858 117922 39954 117978
rect 40010 117922 40078 117978
rect 40134 117922 40202 117978
rect 40258 117922 40326 117978
rect 40382 117922 40478 117978
rect 39858 100350 40478 117922
rect 39858 100294 39954 100350
rect 40010 100294 40078 100350
rect 40134 100294 40202 100350
rect 40258 100294 40326 100350
rect 40382 100294 40478 100350
rect 39858 100226 40478 100294
rect 39858 100170 39954 100226
rect 40010 100170 40078 100226
rect 40134 100170 40202 100226
rect 40258 100170 40326 100226
rect 40382 100170 40478 100226
rect 39858 100102 40478 100170
rect 39858 100046 39954 100102
rect 40010 100046 40078 100102
rect 40134 100046 40202 100102
rect 40258 100046 40326 100102
rect 40382 100046 40478 100102
rect 39858 99978 40478 100046
rect 39858 99922 39954 99978
rect 40010 99922 40078 99978
rect 40134 99922 40202 99978
rect 40258 99922 40326 99978
rect 40382 99922 40478 99978
rect 39858 82350 40478 99922
rect 47852 324324 47908 324334
rect 46956 82740 47012 82750
rect 39858 82294 39954 82350
rect 40010 82294 40078 82350
rect 40134 82294 40202 82350
rect 40258 82294 40326 82350
rect 40382 82294 40478 82350
rect 39858 82226 40478 82294
rect 39858 82170 39954 82226
rect 40010 82170 40078 82226
rect 40134 82170 40202 82226
rect 40258 82170 40326 82226
rect 40382 82170 40478 82226
rect 39858 82102 40478 82170
rect 39858 82046 39954 82102
rect 40010 82046 40078 82102
rect 40134 82046 40202 82102
rect 40258 82046 40326 82102
rect 40382 82046 40478 82102
rect 39858 81978 40478 82046
rect 39858 81922 39954 81978
rect 40010 81922 40078 81978
rect 40134 81922 40202 81978
rect 40258 81922 40326 81978
rect 40382 81922 40478 81978
rect 39858 64350 40478 81922
rect 39858 64294 39954 64350
rect 40010 64294 40078 64350
rect 40134 64294 40202 64350
rect 40258 64294 40326 64350
rect 40382 64294 40478 64350
rect 39858 64226 40478 64294
rect 39858 64170 39954 64226
rect 40010 64170 40078 64226
rect 40134 64170 40202 64226
rect 40258 64170 40326 64226
rect 40382 64170 40478 64226
rect 39858 64102 40478 64170
rect 39858 64046 39954 64102
rect 40010 64046 40078 64102
rect 40134 64046 40202 64102
rect 40258 64046 40326 64102
rect 40382 64046 40478 64102
rect 39858 63978 40478 64046
rect 39858 63922 39954 63978
rect 40010 63922 40078 63978
rect 40134 63922 40202 63978
rect 40258 63922 40326 63978
rect 40382 63922 40478 63978
rect 39858 46350 40478 63922
rect 39858 46294 39954 46350
rect 40010 46294 40078 46350
rect 40134 46294 40202 46350
rect 40258 46294 40326 46350
rect 40382 46294 40478 46350
rect 39858 46226 40478 46294
rect 39858 46170 39954 46226
rect 40010 46170 40078 46226
rect 40134 46170 40202 46226
rect 40258 46170 40326 46226
rect 40382 46170 40478 46226
rect 39858 46102 40478 46170
rect 39858 46046 39954 46102
rect 40010 46046 40078 46102
rect 40134 46046 40202 46102
rect 40258 46046 40326 46102
rect 40382 46046 40478 46102
rect 39858 45978 40478 46046
rect 39858 45922 39954 45978
rect 40010 45922 40078 45978
rect 40134 45922 40202 45978
rect 40258 45922 40326 45978
rect 40382 45922 40478 45978
rect 39858 28350 40478 45922
rect 39858 28294 39954 28350
rect 40010 28294 40078 28350
rect 40134 28294 40202 28350
rect 40258 28294 40326 28350
rect 40382 28294 40478 28350
rect 39858 28226 40478 28294
rect 39858 28170 39954 28226
rect 40010 28170 40078 28226
rect 40134 28170 40202 28226
rect 40258 28170 40326 28226
rect 40382 28170 40478 28226
rect 39858 28102 40478 28170
rect 39858 28046 39954 28102
rect 40010 28046 40078 28102
rect 40134 28046 40202 28102
rect 40258 28046 40326 28102
rect 40382 28046 40478 28102
rect 39858 27978 40478 28046
rect 39858 27922 39954 27978
rect 40010 27922 40078 27978
rect 40134 27922 40202 27978
rect 40258 27922 40326 27978
rect 40382 27922 40478 27978
rect 39858 10350 40478 27922
rect 43596 82404 43652 82414
rect 39858 10294 39954 10350
rect 40010 10294 40078 10350
rect 40134 10294 40202 10350
rect 40258 10294 40326 10350
rect 40382 10294 40478 10350
rect 39858 10226 40478 10294
rect 39858 10170 39954 10226
rect 40010 10170 40078 10226
rect 40134 10170 40202 10226
rect 40258 10170 40326 10226
rect 40382 10170 40478 10226
rect 39858 10102 40478 10170
rect 39858 10046 39954 10102
rect 40010 10046 40078 10102
rect 40134 10046 40202 10102
rect 40258 10046 40326 10102
rect 40382 10046 40478 10102
rect 39858 9978 40478 10046
rect 39858 9922 39954 9978
rect 40010 9922 40078 9978
rect 40134 9922 40202 9978
rect 40258 9922 40326 9978
rect 40382 9922 40478 9978
rect 39858 -1120 40478 9922
rect 42476 16858 42532 16868
rect 40908 5518 40964 5528
rect 40908 3780 40964 5462
rect 40908 3714 40964 3724
rect 42476 3332 42532 16802
rect 43148 8578 43204 8588
rect 43148 3780 43204 8522
rect 43148 3714 43204 3724
rect 42476 3266 42532 3276
rect 43596 1558 43652 82348
rect 46844 81060 46900 81070
rect 46732 34678 46788 34688
rect 46620 31258 46676 31268
rect 46508 25318 46564 25328
rect 44716 15238 44772 15248
rect 44268 5158 44324 5168
rect 44268 3780 44324 5102
rect 44268 3714 44324 3724
rect 44716 3780 44772 15182
rect 45612 11998 45668 12008
rect 44716 3714 44772 3724
rect 44940 7858 44996 7868
rect 44940 3780 44996 7802
rect 44940 3714 44996 3724
rect 45612 3780 45668 11942
rect 46508 8428 46564 25262
rect 45612 3714 45668 3724
rect 46396 8372 46564 8428
rect 46396 3556 46452 8372
rect 46620 3898 46676 31202
rect 46508 3842 46676 3898
rect 46508 3780 46564 3842
rect 46508 3714 46564 3724
rect 46620 3718 46676 3728
rect 46396 3490 46452 3500
rect 46284 3444 46340 3454
rect 45836 3358 45892 3370
rect 45836 3266 45892 3276
rect 43820 3108 43876 3118
rect 43820 2818 43876 3052
rect 43820 2752 43876 2762
rect 46284 2324 46340 3388
rect 46284 2258 46340 2268
rect 43596 1492 43652 1502
rect 46620 1428 46676 3662
rect 46732 3556 46788 34622
rect 46844 14518 46900 81004
rect 46844 14452 46900 14462
rect 46956 14338 47012 82684
rect 47628 82628 47684 82638
rect 47168 58350 47488 58384
rect 47168 58294 47238 58350
rect 47294 58294 47362 58350
rect 47418 58294 47488 58350
rect 47168 58226 47488 58294
rect 47168 58170 47238 58226
rect 47294 58170 47362 58226
rect 47418 58170 47488 58226
rect 47168 58102 47488 58170
rect 47168 58046 47238 58102
rect 47294 58046 47362 58102
rect 47418 58046 47488 58102
rect 47168 57978 47488 58046
rect 47168 57922 47238 57978
rect 47294 57922 47362 57978
rect 47418 57922 47488 57978
rect 47168 57888 47488 57922
rect 47168 40350 47488 40384
rect 47168 40294 47238 40350
rect 47294 40294 47362 40350
rect 47418 40294 47488 40350
rect 47168 40226 47488 40294
rect 47168 40170 47238 40226
rect 47294 40170 47362 40226
rect 47418 40170 47488 40226
rect 47168 40102 47488 40170
rect 47168 40046 47238 40102
rect 47294 40046 47362 40102
rect 47418 40046 47488 40102
rect 47168 39978 47488 40046
rect 47168 39922 47238 39978
rect 47294 39922 47362 39978
rect 47418 39922 47488 39978
rect 47168 39888 47488 39922
rect 47168 22350 47488 22384
rect 47168 22294 47238 22350
rect 47294 22294 47362 22350
rect 47418 22294 47488 22350
rect 47168 22226 47488 22294
rect 47168 22170 47238 22226
rect 47294 22170 47362 22226
rect 47418 22170 47488 22226
rect 47168 22102 47488 22170
rect 47168 22046 47238 22102
rect 47294 22046 47362 22102
rect 47418 22046 47488 22102
rect 47168 21978 47488 22046
rect 47168 21922 47238 21978
rect 47294 21922 47362 21978
rect 47418 21922 47488 21978
rect 47168 21888 47488 21922
rect 46844 14282 47012 14338
rect 46844 3780 46900 14282
rect 46844 3714 46900 3724
rect 46956 14158 47012 14168
rect 46732 3490 46788 3500
rect 46956 3444 47012 14102
rect 47628 3780 47684 82572
rect 47852 81508 47908 324268
rect 66858 310350 67478 327922
rect 66858 310294 66954 310350
rect 67010 310294 67078 310350
rect 67134 310294 67202 310350
rect 67258 310294 67326 310350
rect 67382 310294 67478 310350
rect 66858 310226 67478 310294
rect 66858 310170 66954 310226
rect 67010 310170 67078 310226
rect 67134 310170 67202 310226
rect 67258 310170 67326 310226
rect 67382 310170 67478 310226
rect 66858 310102 67478 310170
rect 66858 310046 66954 310102
rect 67010 310046 67078 310102
rect 67134 310046 67202 310102
rect 67258 310046 67326 310102
rect 67382 310046 67478 310102
rect 66858 309978 67478 310046
rect 66858 309922 66954 309978
rect 67010 309922 67078 309978
rect 67134 309922 67202 309978
rect 67258 309922 67326 309978
rect 67382 309922 67478 309978
rect 66858 292350 67478 309922
rect 66858 292294 66954 292350
rect 67010 292294 67078 292350
rect 67134 292294 67202 292350
rect 67258 292294 67326 292350
rect 67382 292294 67478 292350
rect 66858 292226 67478 292294
rect 66858 292170 66954 292226
rect 67010 292170 67078 292226
rect 67134 292170 67202 292226
rect 67258 292170 67326 292226
rect 67382 292170 67478 292226
rect 66858 292102 67478 292170
rect 66858 292046 66954 292102
rect 67010 292046 67078 292102
rect 67134 292046 67202 292102
rect 67258 292046 67326 292102
rect 67382 292046 67478 292102
rect 66858 291978 67478 292046
rect 66858 291922 66954 291978
rect 67010 291922 67078 291978
rect 67134 291922 67202 291978
rect 67258 291922 67326 291978
rect 67382 291922 67478 291978
rect 66858 274350 67478 291922
rect 66858 274294 66954 274350
rect 67010 274294 67078 274350
rect 67134 274294 67202 274350
rect 67258 274294 67326 274350
rect 67382 274294 67478 274350
rect 66858 274226 67478 274294
rect 66858 274170 66954 274226
rect 67010 274170 67078 274226
rect 67134 274170 67202 274226
rect 67258 274170 67326 274226
rect 67382 274170 67478 274226
rect 66858 274102 67478 274170
rect 66858 274046 66954 274102
rect 67010 274046 67078 274102
rect 67134 274046 67202 274102
rect 67258 274046 67326 274102
rect 67382 274046 67478 274102
rect 66858 273978 67478 274046
rect 66858 273922 66954 273978
rect 67010 273922 67078 273978
rect 67134 273922 67202 273978
rect 67258 273922 67326 273978
rect 67382 273922 67478 273978
rect 66858 256350 67478 273922
rect 66858 256294 66954 256350
rect 67010 256294 67078 256350
rect 67134 256294 67202 256350
rect 67258 256294 67326 256350
rect 67382 256294 67478 256350
rect 66858 256226 67478 256294
rect 66858 256170 66954 256226
rect 67010 256170 67078 256226
rect 67134 256170 67202 256226
rect 67258 256170 67326 256226
rect 67382 256170 67478 256226
rect 66858 256102 67478 256170
rect 66858 256046 66954 256102
rect 67010 256046 67078 256102
rect 67134 256046 67202 256102
rect 67258 256046 67326 256102
rect 67382 256046 67478 256102
rect 66858 255978 67478 256046
rect 66858 255922 66954 255978
rect 67010 255922 67078 255978
rect 67134 255922 67202 255978
rect 67258 255922 67326 255978
rect 67382 255922 67478 255978
rect 66858 238350 67478 255922
rect 66858 238294 66954 238350
rect 67010 238294 67078 238350
rect 67134 238294 67202 238350
rect 67258 238294 67326 238350
rect 67382 238294 67478 238350
rect 66858 238226 67478 238294
rect 66858 238170 66954 238226
rect 67010 238170 67078 238226
rect 67134 238170 67202 238226
rect 67258 238170 67326 238226
rect 67382 238170 67478 238226
rect 66858 238102 67478 238170
rect 66858 238046 66954 238102
rect 67010 238046 67078 238102
rect 67134 238046 67202 238102
rect 67258 238046 67326 238102
rect 67382 238046 67478 238102
rect 66858 237978 67478 238046
rect 66858 237922 66954 237978
rect 67010 237922 67078 237978
rect 67134 237922 67202 237978
rect 67258 237922 67326 237978
rect 67382 237922 67478 237978
rect 66858 220350 67478 237922
rect 66858 220294 66954 220350
rect 67010 220294 67078 220350
rect 67134 220294 67202 220350
rect 67258 220294 67326 220350
rect 67382 220294 67478 220350
rect 66858 220226 67478 220294
rect 66858 220170 66954 220226
rect 67010 220170 67078 220226
rect 67134 220170 67202 220226
rect 67258 220170 67326 220226
rect 67382 220170 67478 220226
rect 66858 220102 67478 220170
rect 66858 220046 66954 220102
rect 67010 220046 67078 220102
rect 67134 220046 67202 220102
rect 67258 220046 67326 220102
rect 67382 220046 67478 220102
rect 66858 219978 67478 220046
rect 66858 219922 66954 219978
rect 67010 219922 67078 219978
rect 67134 219922 67202 219978
rect 67258 219922 67326 219978
rect 67382 219922 67478 219978
rect 66858 202350 67478 219922
rect 66858 202294 66954 202350
rect 67010 202294 67078 202350
rect 67134 202294 67202 202350
rect 67258 202294 67326 202350
rect 67382 202294 67478 202350
rect 66858 202226 67478 202294
rect 66858 202170 66954 202226
rect 67010 202170 67078 202226
rect 67134 202170 67202 202226
rect 67258 202170 67326 202226
rect 67382 202170 67478 202226
rect 66858 202102 67478 202170
rect 66858 202046 66954 202102
rect 67010 202046 67078 202102
rect 67134 202046 67202 202102
rect 67258 202046 67326 202102
rect 67382 202046 67478 202102
rect 66858 201978 67478 202046
rect 66858 201922 66954 201978
rect 67010 201922 67078 201978
rect 67134 201922 67202 201978
rect 67258 201922 67326 201978
rect 67382 201922 67478 201978
rect 66858 184350 67478 201922
rect 66858 184294 66954 184350
rect 67010 184294 67078 184350
rect 67134 184294 67202 184350
rect 67258 184294 67326 184350
rect 67382 184294 67478 184350
rect 66858 184226 67478 184294
rect 66858 184170 66954 184226
rect 67010 184170 67078 184226
rect 67134 184170 67202 184226
rect 67258 184170 67326 184226
rect 67382 184170 67478 184226
rect 66858 184102 67478 184170
rect 66858 184046 66954 184102
rect 67010 184046 67078 184102
rect 67134 184046 67202 184102
rect 67258 184046 67326 184102
rect 67382 184046 67478 184102
rect 66858 183978 67478 184046
rect 66858 183922 66954 183978
rect 67010 183922 67078 183978
rect 67134 183922 67202 183978
rect 67258 183922 67326 183978
rect 67382 183922 67478 183978
rect 66858 166350 67478 183922
rect 66858 166294 66954 166350
rect 67010 166294 67078 166350
rect 67134 166294 67202 166350
rect 67258 166294 67326 166350
rect 67382 166294 67478 166350
rect 66858 166226 67478 166294
rect 66858 166170 66954 166226
rect 67010 166170 67078 166226
rect 67134 166170 67202 166226
rect 67258 166170 67326 166226
rect 67382 166170 67478 166226
rect 66858 166102 67478 166170
rect 66858 166046 66954 166102
rect 67010 166046 67078 166102
rect 67134 166046 67202 166102
rect 67258 166046 67326 166102
rect 67382 166046 67478 166102
rect 66858 165978 67478 166046
rect 66858 165922 66954 165978
rect 67010 165922 67078 165978
rect 67134 165922 67202 165978
rect 67258 165922 67326 165978
rect 67382 165922 67478 165978
rect 66858 148350 67478 165922
rect 66858 148294 66954 148350
rect 67010 148294 67078 148350
rect 67134 148294 67202 148350
rect 67258 148294 67326 148350
rect 67382 148294 67478 148350
rect 66858 148226 67478 148294
rect 66858 148170 66954 148226
rect 67010 148170 67078 148226
rect 67134 148170 67202 148226
rect 67258 148170 67326 148226
rect 67382 148170 67478 148226
rect 66858 148102 67478 148170
rect 66858 148046 66954 148102
rect 67010 148046 67078 148102
rect 67134 148046 67202 148102
rect 67258 148046 67326 148102
rect 67382 148046 67478 148102
rect 66858 147978 67478 148046
rect 66858 147922 66954 147978
rect 67010 147922 67078 147978
rect 67134 147922 67202 147978
rect 67258 147922 67326 147978
rect 67382 147922 67478 147978
rect 66858 130350 67478 147922
rect 66858 130294 66954 130350
rect 67010 130294 67078 130350
rect 67134 130294 67202 130350
rect 67258 130294 67326 130350
rect 67382 130294 67478 130350
rect 66858 130226 67478 130294
rect 66858 130170 66954 130226
rect 67010 130170 67078 130226
rect 67134 130170 67202 130226
rect 67258 130170 67326 130226
rect 67382 130170 67478 130226
rect 66858 130102 67478 130170
rect 66858 130046 66954 130102
rect 67010 130046 67078 130102
rect 67134 130046 67202 130102
rect 67258 130046 67326 130102
rect 67382 130046 67478 130102
rect 66858 129978 67478 130046
rect 66858 129922 66954 129978
rect 67010 129922 67078 129978
rect 67134 129922 67202 129978
rect 67258 129922 67326 129978
rect 67382 129922 67478 129978
rect 66858 112350 67478 129922
rect 66858 112294 66954 112350
rect 67010 112294 67078 112350
rect 67134 112294 67202 112350
rect 67258 112294 67326 112350
rect 67382 112294 67478 112350
rect 66858 112226 67478 112294
rect 66858 112170 66954 112226
rect 67010 112170 67078 112226
rect 67134 112170 67202 112226
rect 67258 112170 67326 112226
rect 67382 112170 67478 112226
rect 66858 112102 67478 112170
rect 66858 112046 66954 112102
rect 67010 112046 67078 112102
rect 67134 112046 67202 112102
rect 67258 112046 67326 112102
rect 67382 112046 67478 112102
rect 66858 111978 67478 112046
rect 66858 111922 66954 111978
rect 67010 111922 67078 111978
rect 67134 111922 67202 111978
rect 67258 111922 67326 111978
rect 67382 111922 67478 111978
rect 66858 94350 67478 111922
rect 66858 94294 66954 94350
rect 67010 94294 67078 94350
rect 67134 94294 67202 94350
rect 67258 94294 67326 94350
rect 67382 94294 67478 94350
rect 66858 94226 67478 94294
rect 66858 94170 66954 94226
rect 67010 94170 67078 94226
rect 67134 94170 67202 94226
rect 67258 94170 67326 94226
rect 67382 94170 67478 94226
rect 66858 94102 67478 94170
rect 66858 94046 66954 94102
rect 67010 94046 67078 94102
rect 67134 94046 67202 94102
rect 67258 94046 67326 94102
rect 67382 94046 67478 94102
rect 66858 93978 67478 94046
rect 66858 93922 66954 93978
rect 67010 93922 67078 93978
rect 67134 93922 67202 93978
rect 67258 93922 67326 93978
rect 67382 93922 67478 93978
rect 47852 81442 47908 81452
rect 48524 82516 48580 82526
rect 48300 80948 48356 80958
rect 47628 3714 47684 3724
rect 48188 36298 48244 36308
rect 48188 3780 48244 36242
rect 48188 3714 48244 3724
rect 46956 3378 47012 3388
rect 48300 3444 48356 80892
rect 48412 80836 48468 80846
rect 48412 3556 48468 80780
rect 48524 3780 48580 82460
rect 65436 79828 65492 79838
rect 60284 76468 60340 76478
rect 52780 76244 52836 76254
rect 49196 47818 49252 47828
rect 48524 3714 48580 3724
rect 48972 44578 49028 44588
rect 48972 3780 49028 44522
rect 48972 3714 49028 3724
rect 49196 3780 49252 47762
rect 51212 37738 51268 37748
rect 50316 24418 50372 24428
rect 50204 19198 50260 19208
rect 50092 14338 50148 14348
rect 49196 3714 49252 3724
rect 49868 12538 49924 12548
rect 49868 3780 49924 12482
rect 49868 3714 49924 3724
rect 48412 3490 48468 3500
rect 48300 3378 48356 3388
rect 50092 3444 50148 14282
rect 50204 3556 50260 19142
rect 50316 3780 50372 24362
rect 50988 17578 51044 17588
rect 50316 3714 50372 3724
rect 50540 15958 50596 15968
rect 50540 3780 50596 15902
rect 50540 3714 50596 3724
rect 50988 3780 51044 17522
rect 50988 3714 51044 3724
rect 51212 3780 51268 37682
rect 51996 30898 52052 30908
rect 51884 24238 51940 24248
rect 51212 3714 51268 3724
rect 51772 19018 51828 19028
rect 51772 3780 51828 18962
rect 51772 3714 51828 3724
rect 50204 3490 50260 3500
rect 50092 3378 50148 3388
rect 51884 3444 51940 24182
rect 51996 3556 52052 30842
rect 52556 29278 52612 29288
rect 52332 14158 52388 14168
rect 52332 3780 52388 14102
rect 52332 3714 52388 3724
rect 51996 3490 52052 3500
rect 51884 3378 51940 3388
rect 52556 3332 52612 29222
rect 52556 3266 52612 3276
rect 49868 2212 49924 2222
rect 48076 1652 48132 1662
rect 48076 1558 48132 1596
rect 48076 1492 48132 1502
rect 48636 1558 48692 1568
rect 46620 1362 46676 1372
rect 48636 1428 48692 1502
rect 49868 1540 49924 2156
rect 49868 1474 49924 1484
rect 48636 1362 48692 1372
rect 52780 1378 52836 76188
rect 57484 73444 57540 73454
rect 56364 72884 56420 72894
rect 56140 69418 56196 69428
rect 54572 59878 54628 59888
rect 53676 56278 53732 56288
rect 53452 29098 53508 29108
rect 53340 24598 53396 24608
rect 53228 8938 53284 8948
rect 53116 4116 53172 4126
rect 53116 2324 53172 4060
rect 53228 3780 53284 8882
rect 53340 3898 53396 24542
rect 53452 20188 53508 29042
rect 53452 20132 53620 20188
rect 53340 3842 53508 3898
rect 53228 3714 53284 3724
rect 53452 3780 53508 3842
rect 53452 3714 53508 3724
rect 53564 3556 53620 20132
rect 53676 7678 53732 56222
rect 54124 41158 54180 41168
rect 53676 7612 53732 7622
rect 53900 20638 53956 20648
rect 53564 3490 53620 3500
rect 53788 5338 53844 5348
rect 53116 2258 53172 2268
rect 52780 1312 52836 1322
rect 53452 1652 53508 1662
rect 53452 1018 53508 1596
rect 53452 952 53508 962
rect 53788 420 53844 5282
rect 53900 3780 53956 20582
rect 54124 8428 54180 41102
rect 53900 3714 53956 3724
rect 54012 8372 54180 8428
rect 54348 32518 54404 32528
rect 54012 1428 54068 8372
rect 54124 4116 54180 4126
rect 54124 3780 54180 4060
rect 54124 3714 54180 3724
rect 54348 3780 54404 32462
rect 54348 3714 54404 3724
rect 54572 3444 54628 59822
rect 55692 42778 55748 42788
rect 55468 20458 55524 20468
rect 55468 20188 55524 20402
rect 55468 20132 55636 20188
rect 55244 17398 55300 17408
rect 55244 3780 55300 17342
rect 55244 3714 55300 3724
rect 55356 13978 55412 13988
rect 55356 3556 55412 13922
rect 55356 3490 55412 3500
rect 55580 3556 55636 20132
rect 55692 3780 55748 42722
rect 56140 20188 56196 69362
rect 56140 20132 56308 20188
rect 55692 3714 55748 3724
rect 55580 3490 55636 3500
rect 56140 3538 56196 3548
rect 54572 3378 54628 3388
rect 56140 3332 56196 3482
rect 56140 3266 56196 3276
rect 56252 1558 56308 20132
rect 56364 13438 56420 72828
rect 57036 51418 57092 51428
rect 56364 13372 56420 13382
rect 56700 18838 56756 18848
rect 56700 3780 56756 18782
rect 56700 3714 56756 3724
rect 56924 15778 56980 15788
rect 56924 3780 56980 15722
rect 57036 6778 57092 51362
rect 57036 6712 57092 6722
rect 57260 10918 57316 10928
rect 56924 3714 56980 3724
rect 57148 4228 57204 4238
rect 56588 3108 56644 3118
rect 56588 2998 56644 3052
rect 56588 2932 56644 2942
rect 57148 2324 57204 4172
rect 57260 3780 57316 10862
rect 57260 3714 57316 3724
rect 57484 3556 57540 73388
rect 58492 73332 58548 73342
rect 58044 73108 58100 73118
rect 57708 54658 57764 54668
rect 57484 3490 57540 3500
rect 57596 4452 57652 4462
rect 57596 3332 57652 4396
rect 57708 3780 57764 54602
rect 57708 3714 57764 3724
rect 57932 7318 57988 7328
rect 57932 3780 57988 7262
rect 57932 3714 57988 3724
rect 57596 3266 57652 3276
rect 57148 2258 57204 2268
rect 56252 1492 56308 1502
rect 54012 1362 54068 1372
rect 58044 1198 58100 73052
rect 58380 37558 58436 37568
rect 58380 3780 58436 37502
rect 58380 3714 58436 3724
rect 58492 3332 58548 73276
rect 58716 61138 58772 61148
rect 58716 25138 58772 61082
rect 59500 47638 59556 47648
rect 59276 40978 59332 40988
rect 58716 25082 58884 25138
rect 58828 20188 58884 25082
rect 58828 20132 59108 20188
rect 59052 3780 59108 20132
rect 58492 3266 58548 3276
rect 58940 3718 58996 3728
rect 59052 3714 59108 3724
rect 59276 3780 59332 40922
rect 59276 3714 59332 3724
rect 59500 3780 59556 47582
rect 60172 36118 60228 36128
rect 59500 3714 59556 3724
rect 59724 7678 59780 7688
rect 59724 3780 59780 7622
rect 59724 3714 59780 3724
rect 60172 3780 60228 36062
rect 60172 3714 60228 3724
rect 58940 2324 58996 3662
rect 60284 3556 60340 76412
rect 60396 76356 60452 76366
rect 60396 3780 60452 76300
rect 62076 74788 62132 74798
rect 61964 74564 62020 74574
rect 61068 52858 61124 52868
rect 60396 3714 60452 3724
rect 60844 32338 60900 32348
rect 60844 3780 60900 32282
rect 60844 3714 60900 3724
rect 61068 3780 61124 52802
rect 61852 37378 61908 37388
rect 61740 35938 61796 35948
rect 61068 3714 61124 3724
rect 61292 25858 61348 25868
rect 61292 3780 61348 25802
rect 61628 4228 61684 4238
rect 61628 3892 61684 4172
rect 61628 3826 61684 3836
rect 61292 3714 61348 3724
rect 61740 3780 61796 35882
rect 61740 3714 61796 3724
rect 60284 3490 60340 3500
rect 61852 3332 61908 37322
rect 61852 3266 61908 3276
rect 58940 2258 58996 2268
rect 60508 3220 60564 3230
rect 60508 2324 60564 3164
rect 60508 2258 60564 2268
rect 58044 1132 58100 1142
rect 58156 1652 58212 1662
rect 53788 354 53844 364
rect 58156 118 58212 1596
rect 61516 1652 61572 1662
rect 61516 1558 61572 1596
rect 61964 1652 62020 74508
rect 62076 3556 62132 74732
rect 65324 74676 65380 74686
rect 65212 70678 65268 70688
rect 62528 64350 62848 64384
rect 62528 64294 62598 64350
rect 62654 64294 62722 64350
rect 62778 64294 62848 64350
rect 62528 64226 62848 64294
rect 62528 64170 62598 64226
rect 62654 64170 62722 64226
rect 62778 64170 62848 64226
rect 62528 64102 62848 64170
rect 62528 64046 62598 64102
rect 62654 64046 62722 64102
rect 62778 64046 62848 64102
rect 62528 63978 62848 64046
rect 62528 63922 62598 63978
rect 62654 63922 62722 63978
rect 62778 63922 62848 63978
rect 62528 63888 62848 63922
rect 63196 62938 63252 62948
rect 62528 46350 62848 46384
rect 62528 46294 62598 46350
rect 62654 46294 62722 46350
rect 62778 46294 62848 46350
rect 62528 46226 62848 46294
rect 62528 46170 62598 46226
rect 62654 46170 62722 46226
rect 62778 46170 62848 46226
rect 62528 46102 62848 46170
rect 62528 46046 62598 46102
rect 62654 46046 62722 46102
rect 62778 46046 62848 46102
rect 62528 45978 62848 46046
rect 62528 45922 62598 45978
rect 62654 45922 62722 45978
rect 62778 45922 62848 45978
rect 62528 45888 62848 45922
rect 62528 28350 62848 28384
rect 62528 28294 62598 28350
rect 62654 28294 62722 28350
rect 62778 28294 62848 28350
rect 62528 28226 62848 28294
rect 62528 28170 62598 28226
rect 62654 28170 62722 28226
rect 62778 28170 62848 28226
rect 62528 28102 62848 28170
rect 62528 28046 62598 28102
rect 62654 28046 62722 28102
rect 62778 28046 62848 28102
rect 62528 27978 62848 28046
rect 62528 27922 62598 27978
rect 62654 27922 62722 27978
rect 62778 27922 62848 27978
rect 62528 27888 62848 27922
rect 62528 10350 62848 10384
rect 62528 10294 62598 10350
rect 62654 10294 62722 10350
rect 62778 10294 62848 10350
rect 62528 10226 62848 10294
rect 62528 10170 62598 10226
rect 62654 10170 62722 10226
rect 62778 10170 62848 10226
rect 62528 10102 62848 10170
rect 62528 10046 62598 10102
rect 62654 10046 62722 10102
rect 62778 10046 62848 10102
rect 62528 9978 62848 10046
rect 62528 9922 62598 9978
rect 62654 9922 62722 9978
rect 62778 9922 62848 9978
rect 62528 9888 62848 9922
rect 62972 6778 63028 6788
rect 62860 4340 62916 4350
rect 62076 3490 62132 3500
rect 62188 4228 62244 4238
rect 61964 1586 62020 1596
rect 61516 1492 61572 1502
rect 62188 868 62244 4172
rect 62860 3780 62916 4284
rect 62860 3714 62916 3724
rect 62972 2660 63028 6722
rect 63196 3332 63252 62882
rect 63644 60058 63700 60068
rect 63532 44758 63588 44768
rect 63420 18658 63476 18668
rect 63308 13798 63364 13808
rect 63308 3668 63364 13742
rect 63308 3602 63364 3612
rect 63196 3266 63252 3276
rect 63420 3108 63476 18602
rect 63532 3220 63588 44702
rect 63644 3780 63700 60002
rect 64428 49618 64484 49628
rect 63980 34498 64036 34508
rect 63644 3714 63700 3724
rect 63756 7138 63812 7148
rect 63756 3668 63812 7082
rect 63980 3780 64036 34442
rect 63980 3714 64036 3724
rect 64204 15598 64260 15608
rect 64204 3780 64260 15542
rect 64204 3714 64260 3724
rect 64428 3780 64484 49562
rect 65100 39538 65156 39548
rect 64876 5698 64932 5708
rect 64428 3714 64484 3724
rect 64764 5518 64820 5528
rect 63756 3602 63812 3612
rect 63532 3154 63588 3164
rect 63980 3332 64036 3342
rect 63420 3042 63476 3052
rect 62972 2594 63028 2604
rect 63196 2660 63252 2670
rect 63196 2436 63252 2604
rect 63196 2370 63252 2380
rect 63980 2324 64036 3276
rect 64764 2660 64820 5462
rect 64876 3668 64932 5642
rect 65100 3780 65156 39482
rect 65212 6598 65268 70622
rect 65212 6532 65268 6542
rect 65100 3714 65156 3724
rect 64876 3602 64932 3612
rect 65324 3668 65380 74620
rect 65436 3780 65492 79772
rect 66858 76350 67478 93922
rect 70578 598172 71198 598268
rect 70578 598116 70674 598172
rect 70730 598116 70798 598172
rect 70854 598116 70922 598172
rect 70978 598116 71046 598172
rect 71102 598116 71198 598172
rect 70578 598048 71198 598116
rect 70578 597992 70674 598048
rect 70730 597992 70798 598048
rect 70854 597992 70922 598048
rect 70978 597992 71046 598048
rect 71102 597992 71198 598048
rect 70578 597924 71198 597992
rect 70578 597868 70674 597924
rect 70730 597868 70798 597924
rect 70854 597868 70922 597924
rect 70978 597868 71046 597924
rect 71102 597868 71198 597924
rect 70578 597800 71198 597868
rect 70578 597744 70674 597800
rect 70730 597744 70798 597800
rect 70854 597744 70922 597800
rect 70978 597744 71046 597800
rect 71102 597744 71198 597800
rect 70578 586350 71198 597744
rect 70578 586294 70674 586350
rect 70730 586294 70798 586350
rect 70854 586294 70922 586350
rect 70978 586294 71046 586350
rect 71102 586294 71198 586350
rect 70578 586226 71198 586294
rect 70578 586170 70674 586226
rect 70730 586170 70798 586226
rect 70854 586170 70922 586226
rect 70978 586170 71046 586226
rect 71102 586170 71198 586226
rect 70578 586102 71198 586170
rect 70578 586046 70674 586102
rect 70730 586046 70798 586102
rect 70854 586046 70922 586102
rect 70978 586046 71046 586102
rect 71102 586046 71198 586102
rect 70578 585978 71198 586046
rect 70578 585922 70674 585978
rect 70730 585922 70798 585978
rect 70854 585922 70922 585978
rect 70978 585922 71046 585978
rect 71102 585922 71198 585978
rect 70578 568350 71198 585922
rect 70578 568294 70674 568350
rect 70730 568294 70798 568350
rect 70854 568294 70922 568350
rect 70978 568294 71046 568350
rect 71102 568294 71198 568350
rect 70578 568226 71198 568294
rect 70578 568170 70674 568226
rect 70730 568170 70798 568226
rect 70854 568170 70922 568226
rect 70978 568170 71046 568226
rect 71102 568170 71198 568226
rect 70578 568102 71198 568170
rect 70578 568046 70674 568102
rect 70730 568046 70798 568102
rect 70854 568046 70922 568102
rect 70978 568046 71046 568102
rect 71102 568046 71198 568102
rect 70578 567978 71198 568046
rect 70578 567922 70674 567978
rect 70730 567922 70798 567978
rect 70854 567922 70922 567978
rect 70978 567922 71046 567978
rect 71102 567922 71198 567978
rect 70578 550350 71198 567922
rect 70578 550294 70674 550350
rect 70730 550294 70798 550350
rect 70854 550294 70922 550350
rect 70978 550294 71046 550350
rect 71102 550294 71198 550350
rect 70578 550226 71198 550294
rect 70578 550170 70674 550226
rect 70730 550170 70798 550226
rect 70854 550170 70922 550226
rect 70978 550170 71046 550226
rect 71102 550170 71198 550226
rect 70578 550102 71198 550170
rect 70578 550046 70674 550102
rect 70730 550046 70798 550102
rect 70854 550046 70922 550102
rect 70978 550046 71046 550102
rect 71102 550046 71198 550102
rect 70578 549978 71198 550046
rect 70578 549922 70674 549978
rect 70730 549922 70798 549978
rect 70854 549922 70922 549978
rect 70978 549922 71046 549978
rect 71102 549922 71198 549978
rect 70578 532350 71198 549922
rect 70578 532294 70674 532350
rect 70730 532294 70798 532350
rect 70854 532294 70922 532350
rect 70978 532294 71046 532350
rect 71102 532294 71198 532350
rect 70578 532226 71198 532294
rect 70578 532170 70674 532226
rect 70730 532170 70798 532226
rect 70854 532170 70922 532226
rect 70978 532170 71046 532226
rect 71102 532170 71198 532226
rect 70578 532102 71198 532170
rect 70578 532046 70674 532102
rect 70730 532046 70798 532102
rect 70854 532046 70922 532102
rect 70978 532046 71046 532102
rect 71102 532046 71198 532102
rect 70578 531978 71198 532046
rect 70578 531922 70674 531978
rect 70730 531922 70798 531978
rect 70854 531922 70922 531978
rect 70978 531922 71046 531978
rect 71102 531922 71198 531978
rect 70578 514350 71198 531922
rect 70578 514294 70674 514350
rect 70730 514294 70798 514350
rect 70854 514294 70922 514350
rect 70978 514294 71046 514350
rect 71102 514294 71198 514350
rect 70578 514226 71198 514294
rect 70578 514170 70674 514226
rect 70730 514170 70798 514226
rect 70854 514170 70922 514226
rect 70978 514170 71046 514226
rect 71102 514170 71198 514226
rect 70578 514102 71198 514170
rect 70578 514046 70674 514102
rect 70730 514046 70798 514102
rect 70854 514046 70922 514102
rect 70978 514046 71046 514102
rect 71102 514046 71198 514102
rect 70578 513978 71198 514046
rect 70578 513922 70674 513978
rect 70730 513922 70798 513978
rect 70854 513922 70922 513978
rect 70978 513922 71046 513978
rect 71102 513922 71198 513978
rect 70578 496350 71198 513922
rect 70578 496294 70674 496350
rect 70730 496294 70798 496350
rect 70854 496294 70922 496350
rect 70978 496294 71046 496350
rect 71102 496294 71198 496350
rect 70578 496226 71198 496294
rect 70578 496170 70674 496226
rect 70730 496170 70798 496226
rect 70854 496170 70922 496226
rect 70978 496170 71046 496226
rect 71102 496170 71198 496226
rect 70578 496102 71198 496170
rect 70578 496046 70674 496102
rect 70730 496046 70798 496102
rect 70854 496046 70922 496102
rect 70978 496046 71046 496102
rect 71102 496046 71198 496102
rect 70578 495978 71198 496046
rect 70578 495922 70674 495978
rect 70730 495922 70798 495978
rect 70854 495922 70922 495978
rect 70978 495922 71046 495978
rect 71102 495922 71198 495978
rect 70578 478350 71198 495922
rect 70578 478294 70674 478350
rect 70730 478294 70798 478350
rect 70854 478294 70922 478350
rect 70978 478294 71046 478350
rect 71102 478294 71198 478350
rect 70578 478226 71198 478294
rect 70578 478170 70674 478226
rect 70730 478170 70798 478226
rect 70854 478170 70922 478226
rect 70978 478170 71046 478226
rect 71102 478170 71198 478226
rect 70578 478102 71198 478170
rect 70578 478046 70674 478102
rect 70730 478046 70798 478102
rect 70854 478046 70922 478102
rect 70978 478046 71046 478102
rect 71102 478046 71198 478102
rect 70578 477978 71198 478046
rect 70578 477922 70674 477978
rect 70730 477922 70798 477978
rect 70854 477922 70922 477978
rect 70978 477922 71046 477978
rect 71102 477922 71198 477978
rect 70578 460350 71198 477922
rect 70578 460294 70674 460350
rect 70730 460294 70798 460350
rect 70854 460294 70922 460350
rect 70978 460294 71046 460350
rect 71102 460294 71198 460350
rect 70578 460226 71198 460294
rect 70578 460170 70674 460226
rect 70730 460170 70798 460226
rect 70854 460170 70922 460226
rect 70978 460170 71046 460226
rect 71102 460170 71198 460226
rect 70578 460102 71198 460170
rect 70578 460046 70674 460102
rect 70730 460046 70798 460102
rect 70854 460046 70922 460102
rect 70978 460046 71046 460102
rect 71102 460046 71198 460102
rect 70578 459978 71198 460046
rect 70578 459922 70674 459978
rect 70730 459922 70798 459978
rect 70854 459922 70922 459978
rect 70978 459922 71046 459978
rect 71102 459922 71198 459978
rect 70578 442350 71198 459922
rect 97578 597212 98198 598268
rect 97578 597156 97674 597212
rect 97730 597156 97798 597212
rect 97854 597156 97922 597212
rect 97978 597156 98046 597212
rect 98102 597156 98198 597212
rect 97578 597088 98198 597156
rect 97578 597032 97674 597088
rect 97730 597032 97798 597088
rect 97854 597032 97922 597088
rect 97978 597032 98046 597088
rect 98102 597032 98198 597088
rect 97578 596964 98198 597032
rect 97578 596908 97674 596964
rect 97730 596908 97798 596964
rect 97854 596908 97922 596964
rect 97978 596908 98046 596964
rect 98102 596908 98198 596964
rect 97578 596840 98198 596908
rect 97578 596784 97674 596840
rect 97730 596784 97798 596840
rect 97854 596784 97922 596840
rect 97978 596784 98046 596840
rect 98102 596784 98198 596840
rect 97578 580350 98198 596784
rect 101298 598172 101918 598268
rect 101298 598116 101394 598172
rect 101450 598116 101518 598172
rect 101574 598116 101642 598172
rect 101698 598116 101766 598172
rect 101822 598116 101918 598172
rect 101298 598048 101918 598116
rect 101298 597992 101394 598048
rect 101450 597992 101518 598048
rect 101574 597992 101642 598048
rect 101698 597992 101766 598048
rect 101822 597992 101918 598048
rect 101298 597924 101918 597992
rect 101298 597868 101394 597924
rect 101450 597868 101518 597924
rect 101574 597868 101642 597924
rect 101698 597868 101766 597924
rect 101822 597868 101918 597924
rect 101298 597800 101918 597868
rect 101298 597744 101394 597800
rect 101450 597744 101518 597800
rect 101574 597744 101642 597800
rect 101698 597744 101766 597800
rect 101822 597744 101918 597800
rect 97578 580294 97674 580350
rect 97730 580294 97798 580350
rect 97854 580294 97922 580350
rect 97978 580294 98046 580350
rect 98102 580294 98198 580350
rect 97578 580226 98198 580294
rect 97578 580170 97674 580226
rect 97730 580170 97798 580226
rect 97854 580170 97922 580226
rect 97978 580170 98046 580226
rect 98102 580170 98198 580226
rect 97578 580102 98198 580170
rect 97578 580046 97674 580102
rect 97730 580046 97798 580102
rect 97854 580046 97922 580102
rect 97978 580046 98046 580102
rect 98102 580046 98198 580102
rect 97578 579978 98198 580046
rect 97578 579922 97674 579978
rect 97730 579922 97798 579978
rect 97854 579922 97922 579978
rect 97978 579922 98046 579978
rect 98102 579922 98198 579978
rect 97578 562350 98198 579922
rect 99260 590212 99316 590222
rect 99260 572908 99316 590156
rect 97578 562294 97674 562350
rect 97730 562294 97798 562350
rect 97854 562294 97922 562350
rect 97978 562294 98046 562350
rect 98102 562294 98198 562350
rect 97578 562226 98198 562294
rect 97578 562170 97674 562226
rect 97730 562170 97798 562226
rect 97854 562170 97922 562226
rect 97978 562170 98046 562226
rect 98102 562170 98198 562226
rect 97578 562102 98198 562170
rect 97578 562046 97674 562102
rect 97730 562046 97798 562102
rect 97854 562046 97922 562102
rect 97978 562046 98046 562102
rect 98102 562046 98198 562102
rect 97578 561978 98198 562046
rect 97578 561922 97674 561978
rect 97730 561922 97798 561978
rect 97854 561922 97922 561978
rect 97978 561922 98046 561978
rect 98102 561922 98198 561978
rect 97578 544350 98198 561922
rect 97578 544294 97674 544350
rect 97730 544294 97798 544350
rect 97854 544294 97922 544350
rect 97978 544294 98046 544350
rect 98102 544294 98198 544350
rect 97578 544226 98198 544294
rect 97578 544170 97674 544226
rect 97730 544170 97798 544226
rect 97854 544170 97922 544226
rect 97978 544170 98046 544226
rect 98102 544170 98198 544226
rect 97578 544102 98198 544170
rect 97578 544046 97674 544102
rect 97730 544046 97798 544102
rect 97854 544046 97922 544102
rect 97978 544046 98046 544102
rect 98102 544046 98198 544102
rect 97578 543978 98198 544046
rect 97578 543922 97674 543978
rect 97730 543922 97798 543978
rect 97854 543922 97922 543978
rect 97978 543922 98046 543978
rect 98102 543922 98198 543978
rect 97578 526350 98198 543922
rect 97578 526294 97674 526350
rect 97730 526294 97798 526350
rect 97854 526294 97922 526350
rect 97978 526294 98046 526350
rect 98102 526294 98198 526350
rect 97578 526226 98198 526294
rect 97578 526170 97674 526226
rect 97730 526170 97798 526226
rect 97854 526170 97922 526226
rect 97978 526170 98046 526226
rect 98102 526170 98198 526226
rect 97578 526102 98198 526170
rect 97578 526046 97674 526102
rect 97730 526046 97798 526102
rect 97854 526046 97922 526102
rect 97978 526046 98046 526102
rect 98102 526046 98198 526102
rect 97578 525978 98198 526046
rect 97578 525922 97674 525978
rect 97730 525922 97798 525978
rect 97854 525922 97922 525978
rect 97978 525922 98046 525978
rect 98102 525922 98198 525978
rect 97578 508350 98198 525922
rect 97578 508294 97674 508350
rect 97730 508294 97798 508350
rect 97854 508294 97922 508350
rect 97978 508294 98046 508350
rect 98102 508294 98198 508350
rect 97578 508226 98198 508294
rect 97578 508170 97674 508226
rect 97730 508170 97798 508226
rect 97854 508170 97922 508226
rect 97978 508170 98046 508226
rect 98102 508170 98198 508226
rect 97578 508102 98198 508170
rect 97578 508046 97674 508102
rect 97730 508046 97798 508102
rect 97854 508046 97922 508102
rect 97978 508046 98046 508102
rect 98102 508046 98198 508102
rect 97578 507978 98198 508046
rect 97578 507922 97674 507978
rect 97730 507922 97798 507978
rect 97854 507922 97922 507978
rect 97978 507922 98046 507978
rect 98102 507922 98198 507978
rect 97578 490350 98198 507922
rect 97578 490294 97674 490350
rect 97730 490294 97798 490350
rect 97854 490294 97922 490350
rect 97978 490294 98046 490350
rect 98102 490294 98198 490350
rect 97578 490226 98198 490294
rect 97578 490170 97674 490226
rect 97730 490170 97798 490226
rect 97854 490170 97922 490226
rect 97978 490170 98046 490226
rect 98102 490170 98198 490226
rect 97578 490102 98198 490170
rect 97578 490046 97674 490102
rect 97730 490046 97798 490102
rect 97854 490046 97922 490102
rect 97978 490046 98046 490102
rect 98102 490046 98198 490102
rect 97578 489978 98198 490046
rect 97578 489922 97674 489978
rect 97730 489922 97798 489978
rect 97854 489922 97922 489978
rect 97978 489922 98046 489978
rect 98102 489922 98198 489978
rect 97578 472350 98198 489922
rect 97578 472294 97674 472350
rect 97730 472294 97798 472350
rect 97854 472294 97922 472350
rect 97978 472294 98046 472350
rect 98102 472294 98198 472350
rect 97578 472226 98198 472294
rect 97578 472170 97674 472226
rect 97730 472170 97798 472226
rect 97854 472170 97922 472226
rect 97978 472170 98046 472226
rect 98102 472170 98198 472226
rect 97578 472102 98198 472170
rect 97578 472046 97674 472102
rect 97730 472046 97798 472102
rect 97854 472046 97922 472102
rect 97978 472046 98046 472102
rect 98102 472046 98198 472102
rect 97578 471978 98198 472046
rect 97578 471922 97674 471978
rect 97730 471922 97798 471978
rect 97854 471922 97922 471978
rect 97978 471922 98046 471978
rect 98102 471922 98198 471978
rect 97578 454350 98198 471922
rect 97578 454294 97674 454350
rect 97730 454294 97798 454350
rect 97854 454294 97922 454350
rect 97978 454294 98046 454350
rect 98102 454294 98198 454350
rect 97578 454226 98198 454294
rect 97578 454170 97674 454226
rect 97730 454170 97798 454226
rect 97854 454170 97922 454226
rect 97978 454170 98046 454226
rect 98102 454170 98198 454226
rect 97578 454102 98198 454170
rect 97578 454046 97674 454102
rect 97730 454046 97798 454102
rect 97854 454046 97922 454102
rect 97978 454046 98046 454102
rect 98102 454046 98198 454102
rect 97578 453978 98198 454046
rect 97578 453922 97674 453978
rect 97730 453922 97798 453978
rect 97854 453922 97922 453978
rect 97978 453922 98046 453978
rect 98102 453922 98198 453978
rect 70578 442294 70674 442350
rect 70730 442294 70798 442350
rect 70854 442294 70922 442350
rect 70978 442294 71046 442350
rect 71102 442294 71198 442350
rect 70578 442226 71198 442294
rect 70578 442170 70674 442226
rect 70730 442170 70798 442226
rect 70854 442170 70922 442226
rect 70978 442170 71046 442226
rect 71102 442170 71198 442226
rect 70578 442102 71198 442170
rect 70578 442046 70674 442102
rect 70730 442046 70798 442102
rect 70854 442046 70922 442102
rect 70978 442046 71046 442102
rect 71102 442046 71198 442102
rect 70578 441978 71198 442046
rect 70578 441922 70674 441978
rect 70730 441922 70798 441978
rect 70854 441922 70922 441978
rect 70978 441922 71046 441978
rect 71102 441922 71198 441978
rect 70578 424350 71198 441922
rect 70578 424294 70674 424350
rect 70730 424294 70798 424350
rect 70854 424294 70922 424350
rect 70978 424294 71046 424350
rect 71102 424294 71198 424350
rect 70578 424226 71198 424294
rect 70578 424170 70674 424226
rect 70730 424170 70798 424226
rect 70854 424170 70922 424226
rect 70978 424170 71046 424226
rect 71102 424170 71198 424226
rect 70578 424102 71198 424170
rect 70578 424046 70674 424102
rect 70730 424046 70798 424102
rect 70854 424046 70922 424102
rect 70978 424046 71046 424102
rect 71102 424046 71198 424102
rect 70578 423978 71198 424046
rect 70578 423922 70674 423978
rect 70730 423922 70798 423978
rect 70854 423922 70922 423978
rect 70978 423922 71046 423978
rect 71102 423922 71198 423978
rect 70578 406350 71198 423922
rect 86492 443268 86548 443278
rect 70578 406294 70674 406350
rect 70730 406294 70798 406350
rect 70854 406294 70922 406350
rect 70978 406294 71046 406350
rect 71102 406294 71198 406350
rect 70578 406226 71198 406294
rect 70578 406170 70674 406226
rect 70730 406170 70798 406226
rect 70854 406170 70922 406226
rect 70978 406170 71046 406226
rect 71102 406170 71198 406226
rect 70578 406102 71198 406170
rect 70578 406046 70674 406102
rect 70730 406046 70798 406102
rect 70854 406046 70922 406102
rect 70978 406046 71046 406102
rect 71102 406046 71198 406102
rect 70578 405978 71198 406046
rect 70578 405922 70674 405978
rect 70730 405922 70798 405978
rect 70854 405922 70922 405978
rect 70978 405922 71046 405978
rect 71102 405922 71198 405978
rect 70578 388350 71198 405922
rect 70578 388294 70674 388350
rect 70730 388294 70798 388350
rect 70854 388294 70922 388350
rect 70978 388294 71046 388350
rect 71102 388294 71198 388350
rect 70578 388226 71198 388294
rect 70578 388170 70674 388226
rect 70730 388170 70798 388226
rect 70854 388170 70922 388226
rect 70978 388170 71046 388226
rect 71102 388170 71198 388226
rect 70578 388102 71198 388170
rect 70578 388046 70674 388102
rect 70730 388046 70798 388102
rect 70854 388046 70922 388102
rect 70978 388046 71046 388102
rect 71102 388046 71198 388102
rect 70578 387978 71198 388046
rect 70578 387922 70674 387978
rect 70730 387922 70798 387978
rect 70854 387922 70922 387978
rect 70978 387922 71046 387978
rect 71102 387922 71198 387978
rect 70578 370350 71198 387922
rect 70578 370294 70674 370350
rect 70730 370294 70798 370350
rect 70854 370294 70922 370350
rect 70978 370294 71046 370350
rect 71102 370294 71198 370350
rect 70578 370226 71198 370294
rect 70578 370170 70674 370226
rect 70730 370170 70798 370226
rect 70854 370170 70922 370226
rect 70978 370170 71046 370226
rect 71102 370170 71198 370226
rect 70578 370102 71198 370170
rect 70578 370046 70674 370102
rect 70730 370046 70798 370102
rect 70854 370046 70922 370102
rect 70978 370046 71046 370102
rect 71102 370046 71198 370102
rect 70578 369978 71198 370046
rect 70578 369922 70674 369978
rect 70730 369922 70798 369978
rect 70854 369922 70922 369978
rect 70978 369922 71046 369978
rect 71102 369922 71198 369978
rect 70578 352350 71198 369922
rect 70578 352294 70674 352350
rect 70730 352294 70798 352350
rect 70854 352294 70922 352350
rect 70978 352294 71046 352350
rect 71102 352294 71198 352350
rect 70578 352226 71198 352294
rect 70578 352170 70674 352226
rect 70730 352170 70798 352226
rect 70854 352170 70922 352226
rect 70978 352170 71046 352226
rect 71102 352170 71198 352226
rect 70578 352102 71198 352170
rect 70578 352046 70674 352102
rect 70730 352046 70798 352102
rect 70854 352046 70922 352102
rect 70978 352046 71046 352102
rect 71102 352046 71198 352102
rect 70578 351978 71198 352046
rect 70578 351922 70674 351978
rect 70730 351922 70798 351978
rect 70854 351922 70922 351978
rect 70978 351922 71046 351978
rect 71102 351922 71198 351978
rect 70578 334350 71198 351922
rect 70578 334294 70674 334350
rect 70730 334294 70798 334350
rect 70854 334294 70922 334350
rect 70978 334294 71046 334350
rect 71102 334294 71198 334350
rect 70578 334226 71198 334294
rect 70578 334170 70674 334226
rect 70730 334170 70798 334226
rect 70854 334170 70922 334226
rect 70978 334170 71046 334226
rect 71102 334170 71198 334226
rect 70578 334102 71198 334170
rect 70578 334046 70674 334102
rect 70730 334046 70798 334102
rect 70854 334046 70922 334102
rect 70978 334046 71046 334102
rect 71102 334046 71198 334102
rect 70578 333978 71198 334046
rect 70578 333922 70674 333978
rect 70730 333922 70798 333978
rect 70854 333922 70922 333978
rect 70978 333922 71046 333978
rect 71102 333922 71198 333978
rect 70578 316350 71198 333922
rect 70578 316294 70674 316350
rect 70730 316294 70798 316350
rect 70854 316294 70922 316350
rect 70978 316294 71046 316350
rect 71102 316294 71198 316350
rect 70578 316226 71198 316294
rect 70578 316170 70674 316226
rect 70730 316170 70798 316226
rect 70854 316170 70922 316226
rect 70978 316170 71046 316226
rect 71102 316170 71198 316226
rect 70578 316102 71198 316170
rect 70578 316046 70674 316102
rect 70730 316046 70798 316102
rect 70854 316046 70922 316102
rect 70978 316046 71046 316102
rect 71102 316046 71198 316102
rect 70578 315978 71198 316046
rect 70578 315922 70674 315978
rect 70730 315922 70798 315978
rect 70854 315922 70922 315978
rect 70978 315922 71046 315978
rect 71102 315922 71198 315978
rect 70578 298350 71198 315922
rect 70578 298294 70674 298350
rect 70730 298294 70798 298350
rect 70854 298294 70922 298350
rect 70978 298294 71046 298350
rect 71102 298294 71198 298350
rect 70578 298226 71198 298294
rect 70578 298170 70674 298226
rect 70730 298170 70798 298226
rect 70854 298170 70922 298226
rect 70978 298170 71046 298226
rect 71102 298170 71198 298226
rect 70578 298102 71198 298170
rect 70578 298046 70674 298102
rect 70730 298046 70798 298102
rect 70854 298046 70922 298102
rect 70978 298046 71046 298102
rect 71102 298046 71198 298102
rect 70578 297978 71198 298046
rect 70578 297922 70674 297978
rect 70730 297922 70798 297978
rect 70854 297922 70922 297978
rect 70978 297922 71046 297978
rect 71102 297922 71198 297978
rect 70578 280350 71198 297922
rect 70578 280294 70674 280350
rect 70730 280294 70798 280350
rect 70854 280294 70922 280350
rect 70978 280294 71046 280350
rect 71102 280294 71198 280350
rect 70578 280226 71198 280294
rect 70578 280170 70674 280226
rect 70730 280170 70798 280226
rect 70854 280170 70922 280226
rect 70978 280170 71046 280226
rect 71102 280170 71198 280226
rect 70578 280102 71198 280170
rect 70578 280046 70674 280102
rect 70730 280046 70798 280102
rect 70854 280046 70922 280102
rect 70978 280046 71046 280102
rect 71102 280046 71198 280102
rect 70578 279978 71198 280046
rect 70578 279922 70674 279978
rect 70730 279922 70798 279978
rect 70854 279922 70922 279978
rect 70978 279922 71046 279978
rect 71102 279922 71198 279978
rect 70578 262350 71198 279922
rect 70578 262294 70674 262350
rect 70730 262294 70798 262350
rect 70854 262294 70922 262350
rect 70978 262294 71046 262350
rect 71102 262294 71198 262350
rect 70578 262226 71198 262294
rect 70578 262170 70674 262226
rect 70730 262170 70798 262226
rect 70854 262170 70922 262226
rect 70978 262170 71046 262226
rect 71102 262170 71198 262226
rect 70578 262102 71198 262170
rect 70578 262046 70674 262102
rect 70730 262046 70798 262102
rect 70854 262046 70922 262102
rect 70978 262046 71046 262102
rect 71102 262046 71198 262102
rect 70578 261978 71198 262046
rect 70578 261922 70674 261978
rect 70730 261922 70798 261978
rect 70854 261922 70922 261978
rect 70978 261922 71046 261978
rect 71102 261922 71198 261978
rect 70578 244350 71198 261922
rect 70578 244294 70674 244350
rect 70730 244294 70798 244350
rect 70854 244294 70922 244350
rect 70978 244294 71046 244350
rect 71102 244294 71198 244350
rect 70578 244226 71198 244294
rect 70578 244170 70674 244226
rect 70730 244170 70798 244226
rect 70854 244170 70922 244226
rect 70978 244170 71046 244226
rect 71102 244170 71198 244226
rect 70578 244102 71198 244170
rect 70578 244046 70674 244102
rect 70730 244046 70798 244102
rect 70854 244046 70922 244102
rect 70978 244046 71046 244102
rect 71102 244046 71198 244102
rect 70578 243978 71198 244046
rect 70578 243922 70674 243978
rect 70730 243922 70798 243978
rect 70854 243922 70922 243978
rect 70978 243922 71046 243978
rect 71102 243922 71198 243978
rect 70578 226350 71198 243922
rect 70578 226294 70674 226350
rect 70730 226294 70798 226350
rect 70854 226294 70922 226350
rect 70978 226294 71046 226350
rect 71102 226294 71198 226350
rect 70578 226226 71198 226294
rect 70578 226170 70674 226226
rect 70730 226170 70798 226226
rect 70854 226170 70922 226226
rect 70978 226170 71046 226226
rect 71102 226170 71198 226226
rect 70578 226102 71198 226170
rect 70578 226046 70674 226102
rect 70730 226046 70798 226102
rect 70854 226046 70922 226102
rect 70978 226046 71046 226102
rect 71102 226046 71198 226102
rect 70578 225978 71198 226046
rect 70578 225922 70674 225978
rect 70730 225922 70798 225978
rect 70854 225922 70922 225978
rect 70978 225922 71046 225978
rect 71102 225922 71198 225978
rect 70578 208350 71198 225922
rect 70578 208294 70674 208350
rect 70730 208294 70798 208350
rect 70854 208294 70922 208350
rect 70978 208294 71046 208350
rect 71102 208294 71198 208350
rect 70578 208226 71198 208294
rect 70578 208170 70674 208226
rect 70730 208170 70798 208226
rect 70854 208170 70922 208226
rect 70978 208170 71046 208226
rect 71102 208170 71198 208226
rect 70578 208102 71198 208170
rect 70578 208046 70674 208102
rect 70730 208046 70798 208102
rect 70854 208046 70922 208102
rect 70978 208046 71046 208102
rect 71102 208046 71198 208102
rect 70578 207978 71198 208046
rect 70578 207922 70674 207978
rect 70730 207922 70798 207978
rect 70854 207922 70922 207978
rect 70978 207922 71046 207978
rect 71102 207922 71198 207978
rect 70578 190350 71198 207922
rect 70578 190294 70674 190350
rect 70730 190294 70798 190350
rect 70854 190294 70922 190350
rect 70978 190294 71046 190350
rect 71102 190294 71198 190350
rect 70578 190226 71198 190294
rect 70578 190170 70674 190226
rect 70730 190170 70798 190226
rect 70854 190170 70922 190226
rect 70978 190170 71046 190226
rect 71102 190170 71198 190226
rect 70578 190102 71198 190170
rect 70578 190046 70674 190102
rect 70730 190046 70798 190102
rect 70854 190046 70922 190102
rect 70978 190046 71046 190102
rect 71102 190046 71198 190102
rect 70578 189978 71198 190046
rect 70578 189922 70674 189978
rect 70730 189922 70798 189978
rect 70854 189922 70922 189978
rect 70978 189922 71046 189978
rect 71102 189922 71198 189978
rect 70578 172350 71198 189922
rect 70578 172294 70674 172350
rect 70730 172294 70798 172350
rect 70854 172294 70922 172350
rect 70978 172294 71046 172350
rect 71102 172294 71198 172350
rect 70578 172226 71198 172294
rect 70578 172170 70674 172226
rect 70730 172170 70798 172226
rect 70854 172170 70922 172226
rect 70978 172170 71046 172226
rect 71102 172170 71198 172226
rect 70578 172102 71198 172170
rect 70578 172046 70674 172102
rect 70730 172046 70798 172102
rect 70854 172046 70922 172102
rect 70978 172046 71046 172102
rect 71102 172046 71198 172102
rect 70578 171978 71198 172046
rect 70578 171922 70674 171978
rect 70730 171922 70798 171978
rect 70854 171922 70922 171978
rect 70978 171922 71046 171978
rect 71102 171922 71198 171978
rect 70578 154350 71198 171922
rect 70578 154294 70674 154350
rect 70730 154294 70798 154350
rect 70854 154294 70922 154350
rect 70978 154294 71046 154350
rect 71102 154294 71198 154350
rect 70578 154226 71198 154294
rect 70578 154170 70674 154226
rect 70730 154170 70798 154226
rect 70854 154170 70922 154226
rect 70978 154170 71046 154226
rect 71102 154170 71198 154226
rect 70578 154102 71198 154170
rect 70578 154046 70674 154102
rect 70730 154046 70798 154102
rect 70854 154046 70922 154102
rect 70978 154046 71046 154102
rect 71102 154046 71198 154102
rect 70578 153978 71198 154046
rect 70578 153922 70674 153978
rect 70730 153922 70798 153978
rect 70854 153922 70922 153978
rect 70978 153922 71046 153978
rect 71102 153922 71198 153978
rect 70578 136350 71198 153922
rect 70578 136294 70674 136350
rect 70730 136294 70798 136350
rect 70854 136294 70922 136350
rect 70978 136294 71046 136350
rect 71102 136294 71198 136350
rect 70578 136226 71198 136294
rect 70578 136170 70674 136226
rect 70730 136170 70798 136226
rect 70854 136170 70922 136226
rect 70978 136170 71046 136226
rect 71102 136170 71198 136226
rect 70578 136102 71198 136170
rect 70578 136046 70674 136102
rect 70730 136046 70798 136102
rect 70854 136046 70922 136102
rect 70978 136046 71046 136102
rect 71102 136046 71198 136102
rect 70578 135978 71198 136046
rect 70578 135922 70674 135978
rect 70730 135922 70798 135978
rect 70854 135922 70922 135978
rect 70978 135922 71046 135978
rect 71102 135922 71198 135978
rect 70578 118350 71198 135922
rect 70578 118294 70674 118350
rect 70730 118294 70798 118350
rect 70854 118294 70922 118350
rect 70978 118294 71046 118350
rect 71102 118294 71198 118350
rect 70578 118226 71198 118294
rect 70578 118170 70674 118226
rect 70730 118170 70798 118226
rect 70854 118170 70922 118226
rect 70978 118170 71046 118226
rect 71102 118170 71198 118226
rect 70578 118102 71198 118170
rect 70578 118046 70674 118102
rect 70730 118046 70798 118102
rect 70854 118046 70922 118102
rect 70978 118046 71046 118102
rect 71102 118046 71198 118102
rect 70578 117978 71198 118046
rect 70578 117922 70674 117978
rect 70730 117922 70798 117978
rect 70854 117922 70922 117978
rect 70978 117922 71046 117978
rect 71102 117922 71198 117978
rect 70578 100350 71198 117922
rect 70578 100294 70674 100350
rect 70730 100294 70798 100350
rect 70854 100294 70922 100350
rect 70978 100294 71046 100350
rect 71102 100294 71198 100350
rect 70578 100226 71198 100294
rect 70578 100170 70674 100226
rect 70730 100170 70798 100226
rect 70854 100170 70922 100226
rect 70978 100170 71046 100226
rect 71102 100170 71198 100226
rect 70578 100102 71198 100170
rect 70578 100046 70674 100102
rect 70730 100046 70798 100102
rect 70854 100046 70922 100102
rect 70978 100046 71046 100102
rect 71102 100046 71198 100102
rect 70578 99978 71198 100046
rect 70578 99922 70674 99978
rect 70730 99922 70798 99978
rect 70854 99922 70922 99978
rect 70978 99922 71046 99978
rect 71102 99922 71198 99978
rect 70578 82350 71198 99922
rect 70578 82294 70674 82350
rect 70730 82294 70798 82350
rect 70854 82294 70922 82350
rect 70978 82294 71046 82350
rect 71102 82294 71198 82350
rect 70578 82226 71198 82294
rect 70578 82170 70674 82226
rect 70730 82170 70798 82226
rect 70854 82170 70922 82226
rect 70978 82170 71046 82226
rect 71102 82170 71198 82226
rect 70578 82102 71198 82170
rect 70578 82046 70674 82102
rect 70730 82046 70798 82102
rect 70854 82046 70922 82102
rect 70978 82046 71046 82102
rect 71102 82046 71198 82102
rect 70578 81978 71198 82046
rect 70578 81922 70674 81978
rect 70730 81922 70798 81978
rect 70854 81922 70922 81978
rect 70978 81922 71046 81978
rect 71102 81922 71198 81978
rect 70364 80724 70420 80734
rect 66858 76294 66954 76350
rect 67010 76294 67078 76350
rect 67134 76294 67202 76350
rect 67258 76294 67326 76350
rect 67382 76294 67478 76350
rect 66858 76226 67478 76294
rect 66858 76170 66954 76226
rect 67010 76170 67078 76226
rect 67134 76170 67202 76226
rect 67258 76170 67326 76226
rect 67382 76170 67478 76226
rect 66858 76102 67478 76170
rect 66858 76046 66954 76102
rect 67010 76046 67078 76102
rect 67134 76046 67202 76102
rect 67258 76046 67326 76102
rect 67382 76046 67478 76102
rect 66858 75978 67478 76046
rect 66858 75922 66954 75978
rect 67010 75922 67078 75978
rect 67134 75922 67202 75978
rect 67258 75922 67326 75978
rect 67382 75922 67478 75978
rect 66668 72996 66724 73006
rect 66556 67618 66612 67628
rect 66444 56458 66500 56468
rect 66332 32698 66388 32708
rect 66220 26218 66276 26228
rect 65436 3714 65492 3724
rect 65996 13438 66052 13448
rect 65996 3780 66052 13382
rect 65996 3714 66052 3724
rect 65324 3602 65380 3612
rect 66220 3668 66276 26162
rect 66332 3780 66388 32642
rect 66332 3714 66388 3724
rect 66220 3602 66276 3612
rect 66444 3668 66500 56402
rect 66444 3602 66500 3612
rect 66556 3388 66612 67562
rect 66668 3780 66724 72940
rect 66668 3714 66724 3724
rect 66858 58350 67478 75922
rect 70252 78260 70308 78270
rect 66858 58294 66954 58350
rect 67010 58294 67078 58350
rect 67134 58294 67202 58350
rect 67258 58294 67326 58350
rect 67382 58294 67478 58350
rect 66858 58226 67478 58294
rect 66858 58170 66954 58226
rect 67010 58170 67078 58226
rect 67134 58170 67202 58226
rect 67258 58170 67326 58226
rect 67382 58170 67478 58226
rect 66858 58102 67478 58170
rect 66858 58046 66954 58102
rect 67010 58046 67078 58102
rect 67134 58046 67202 58102
rect 67258 58046 67326 58102
rect 67382 58046 67478 58102
rect 66858 57978 67478 58046
rect 66858 57922 66954 57978
rect 67010 57922 67078 57978
rect 67134 57922 67202 57978
rect 67258 57922 67326 57978
rect 67382 57922 67478 57978
rect 66858 40350 67478 57922
rect 66858 40294 66954 40350
rect 67010 40294 67078 40350
rect 67134 40294 67202 40350
rect 67258 40294 67326 40350
rect 67382 40294 67478 40350
rect 66858 40226 67478 40294
rect 66858 40170 66954 40226
rect 67010 40170 67078 40226
rect 67134 40170 67202 40226
rect 67258 40170 67326 40226
rect 67382 40170 67478 40226
rect 66858 40102 67478 40170
rect 66858 40046 66954 40102
rect 67010 40046 67078 40102
rect 67134 40046 67202 40102
rect 67258 40046 67326 40102
rect 67382 40046 67478 40102
rect 66858 39978 67478 40046
rect 66858 39922 66954 39978
rect 67010 39922 67078 39978
rect 67134 39922 67202 39978
rect 67258 39922 67326 39978
rect 67382 39922 67478 39978
rect 66858 22350 67478 39922
rect 66858 22294 66954 22350
rect 67010 22294 67078 22350
rect 67134 22294 67202 22350
rect 67258 22294 67326 22350
rect 67382 22294 67478 22350
rect 66858 22226 67478 22294
rect 66858 22170 66954 22226
rect 67010 22170 67078 22226
rect 67134 22170 67202 22226
rect 67258 22170 67326 22226
rect 67382 22170 67478 22226
rect 66858 22102 67478 22170
rect 66858 22046 66954 22102
rect 67010 22046 67078 22102
rect 67134 22046 67202 22102
rect 67258 22046 67326 22102
rect 67382 22046 67478 22102
rect 66858 21978 67478 22046
rect 66858 21922 66954 21978
rect 67010 21922 67078 21978
rect 67134 21922 67202 21978
rect 67258 21922 67326 21978
rect 67382 21922 67478 21978
rect 66858 4350 67478 21922
rect 66858 4294 66954 4350
rect 67010 4294 67078 4350
rect 67134 4294 67202 4350
rect 67258 4294 67326 4350
rect 67382 4294 67478 4350
rect 66858 4226 67478 4294
rect 66858 4170 66954 4226
rect 67010 4170 67078 4226
rect 67134 4170 67202 4226
rect 67258 4170 67326 4226
rect 67382 4170 67478 4226
rect 66858 4102 67478 4170
rect 66858 4046 66954 4102
rect 67010 4046 67078 4102
rect 67134 4046 67202 4102
rect 67258 4046 67326 4102
rect 67382 4046 67478 4102
rect 66858 3978 67478 4046
rect 66858 3922 66954 3978
rect 67010 3922 67078 3978
rect 67134 3922 67202 3978
rect 67258 3922 67326 3978
rect 67382 3922 67478 3978
rect 66556 3332 66724 3388
rect 66668 3108 66724 3332
rect 66668 3042 66724 3052
rect 64764 2594 64820 2604
rect 63980 2258 64036 2268
rect 62412 1540 62468 1550
rect 62412 1378 62468 1484
rect 62412 1312 62468 1322
rect 65772 1540 65828 1550
rect 65772 1198 65828 1484
rect 65772 1132 65828 1142
rect 62188 802 62244 812
rect 58156 52 58212 62
rect 39858 -1176 39954 -1120
rect 40010 -1176 40078 -1120
rect 40134 -1176 40202 -1120
rect 40258 -1176 40326 -1120
rect 40382 -1176 40478 -1120
rect 39858 -1244 40478 -1176
rect 39858 -1300 39954 -1244
rect 40010 -1300 40078 -1244
rect 40134 -1300 40202 -1244
rect 40258 -1300 40326 -1244
rect 40382 -1300 40478 -1244
rect 39858 -1368 40478 -1300
rect 39858 -1424 39954 -1368
rect 40010 -1424 40078 -1368
rect 40134 -1424 40202 -1368
rect 40258 -1424 40326 -1368
rect 40382 -1424 40478 -1368
rect 39858 -1492 40478 -1424
rect 39858 -1548 39954 -1492
rect 40010 -1548 40078 -1492
rect 40134 -1548 40202 -1492
rect 40258 -1548 40326 -1492
rect 40382 -1548 40478 -1492
rect 39858 -1644 40478 -1548
rect 66858 -160 67478 3922
rect 67788 74452 67844 74462
rect 67788 3780 67844 74396
rect 69132 74340 69188 74350
rect 68796 72772 68852 72782
rect 68684 70858 68740 70868
rect 68572 52678 68628 52688
rect 68460 32158 68516 32168
rect 68348 6598 68404 6608
rect 67788 3714 67844 3724
rect 68124 4116 68180 4126
rect 68124 2772 68180 4060
rect 68348 3108 68404 6542
rect 68460 3780 68516 32102
rect 68460 3714 68516 3724
rect 68572 3556 68628 52622
rect 68572 3490 68628 3500
rect 68684 3220 68740 70802
rect 68796 3668 68852 72716
rect 68908 4116 68964 4126
rect 68908 3780 68964 4060
rect 68908 3714 68964 3724
rect 69132 3780 69188 74284
rect 70140 69058 70196 69068
rect 69132 3714 69188 3724
rect 69468 54838 69524 54848
rect 69468 3780 69524 54782
rect 70028 30358 70084 30368
rect 69468 3714 69524 3724
rect 69916 22798 69972 22808
rect 68796 3602 68852 3612
rect 69916 3668 69972 22742
rect 69916 3602 69972 3612
rect 70028 3388 70084 30302
rect 70140 4116 70196 69002
rect 70140 4050 70196 4060
rect 70252 3898 70308 78204
rect 70140 3842 70308 3898
rect 70140 3780 70196 3842
rect 70140 3714 70196 3724
rect 70364 3780 70420 80668
rect 70364 3714 70420 3724
rect 70578 64350 71198 81922
rect 76412 416836 76468 416846
rect 75852 79604 75908 79614
rect 70578 64294 70674 64350
rect 70730 64294 70798 64350
rect 70854 64294 70922 64350
rect 70978 64294 71046 64350
rect 71102 64294 71198 64350
rect 70578 64226 71198 64294
rect 70578 64170 70674 64226
rect 70730 64170 70798 64226
rect 70854 64170 70922 64226
rect 70978 64170 71046 64226
rect 71102 64170 71198 64226
rect 70578 64102 71198 64170
rect 70578 64046 70674 64102
rect 70730 64046 70798 64102
rect 70854 64046 70922 64102
rect 70978 64046 71046 64102
rect 71102 64046 71198 64102
rect 70578 63978 71198 64046
rect 70578 63922 70674 63978
rect 70730 63922 70798 63978
rect 70854 63922 70922 63978
rect 70978 63922 71046 63978
rect 71102 63922 71198 63978
rect 70578 46350 71198 63922
rect 70578 46294 70674 46350
rect 70730 46294 70798 46350
rect 70854 46294 70922 46350
rect 70978 46294 71046 46350
rect 71102 46294 71198 46350
rect 70578 46226 71198 46294
rect 70578 46170 70674 46226
rect 70730 46170 70798 46226
rect 70854 46170 70922 46226
rect 70978 46170 71046 46226
rect 71102 46170 71198 46226
rect 70578 46102 71198 46170
rect 70578 46046 70674 46102
rect 70730 46046 70798 46102
rect 70854 46046 70922 46102
rect 70978 46046 71046 46102
rect 71102 46046 71198 46102
rect 70578 45978 71198 46046
rect 70578 45922 70674 45978
rect 70730 45922 70798 45978
rect 70854 45922 70922 45978
rect 70978 45922 71046 45978
rect 71102 45922 71198 45978
rect 70578 28350 71198 45922
rect 70578 28294 70674 28350
rect 70730 28294 70798 28350
rect 70854 28294 70922 28350
rect 70978 28294 71046 28350
rect 71102 28294 71198 28350
rect 70578 28226 71198 28294
rect 70578 28170 70674 28226
rect 70730 28170 70798 28226
rect 70854 28170 70922 28226
rect 70978 28170 71046 28226
rect 71102 28170 71198 28226
rect 70578 28102 71198 28170
rect 70578 28046 70674 28102
rect 70730 28046 70798 28102
rect 70854 28046 70922 28102
rect 70978 28046 71046 28102
rect 71102 28046 71198 28102
rect 70578 27978 71198 28046
rect 70578 27922 70674 27978
rect 70730 27922 70798 27978
rect 70854 27922 70922 27978
rect 70978 27922 71046 27978
rect 71102 27922 71198 27978
rect 70578 10350 71198 27922
rect 71708 78148 71764 78158
rect 70578 10294 70674 10350
rect 70730 10294 70798 10350
rect 70854 10294 70922 10350
rect 70978 10294 71046 10350
rect 71102 10294 71198 10350
rect 70578 10226 71198 10294
rect 70578 10170 70674 10226
rect 70730 10170 70798 10226
rect 70854 10170 70922 10226
rect 70978 10170 71046 10226
rect 71102 10170 71198 10226
rect 70578 10102 71198 10170
rect 70578 10046 70674 10102
rect 70730 10046 70798 10102
rect 70854 10046 70922 10102
rect 70978 10046 71046 10102
rect 71102 10046 71198 10102
rect 70578 9978 71198 10046
rect 70578 9922 70674 9978
rect 70730 9922 70798 9978
rect 70854 9922 70922 9978
rect 70978 9922 71046 9978
rect 71102 9922 71198 9978
rect 68684 3154 68740 3164
rect 69804 3332 70084 3388
rect 69804 3220 69860 3332
rect 69804 3154 69860 3164
rect 68348 3042 68404 3052
rect 68124 2706 68180 2716
rect 66858 -216 66954 -160
rect 67010 -216 67078 -160
rect 67134 -216 67202 -160
rect 67258 -216 67326 -160
rect 67382 -216 67478 -160
rect 66858 -284 67478 -216
rect 66858 -340 66954 -284
rect 67010 -340 67078 -284
rect 67134 -340 67202 -284
rect 67258 -340 67326 -284
rect 67382 -340 67478 -284
rect 66858 -408 67478 -340
rect 66858 -464 66954 -408
rect 67010 -464 67078 -408
rect 67134 -464 67202 -408
rect 67258 -464 67326 -408
rect 67382 -464 67478 -408
rect 66858 -532 67478 -464
rect 66858 -588 66954 -532
rect 67010 -588 67078 -532
rect 67134 -588 67202 -532
rect 67258 -588 67326 -532
rect 67382 -588 67478 -532
rect 66858 -1644 67478 -588
rect 70578 -1120 71198 9922
rect 71596 13438 71652 13448
rect 71596 3780 71652 13382
rect 71596 3714 71652 3724
rect 71708 3668 71764 78092
rect 73052 77924 73108 77934
rect 72492 76132 72548 76142
rect 72044 51598 72100 51608
rect 71932 25138 71988 25148
rect 71932 3780 71988 25082
rect 71932 3714 71988 3724
rect 71708 3602 71764 3612
rect 72044 3444 72100 51542
rect 72268 4116 72324 4126
rect 72268 3780 72324 4060
rect 72268 3714 72324 3724
rect 72492 3780 72548 76076
rect 72492 3714 72548 3724
rect 72716 74228 72772 74238
rect 72716 3780 72772 74172
rect 72940 42418 72996 42428
rect 72940 34498 72996 42362
rect 72940 34432 72996 34442
rect 73052 30358 73108 77868
rect 74508 77812 74564 77822
rect 73836 76020 73892 76030
rect 73052 30292 73108 30302
rect 73164 59698 73220 59708
rect 73052 26938 73108 26948
rect 73052 24598 73108 26882
rect 73164 26218 73220 59642
rect 73724 40798 73780 40808
rect 73164 26152 73220 26162
rect 73612 30538 73668 30548
rect 73052 24532 73108 24542
rect 73500 26038 73556 26048
rect 72716 3714 72772 3724
rect 73164 17218 73220 17228
rect 73164 3780 73220 17162
rect 73164 3714 73220 3724
rect 73500 3780 73556 25982
rect 73500 3714 73556 3724
rect 73612 3668 73668 30482
rect 73724 4116 73780 40742
rect 73724 4050 73780 4060
rect 73836 3780 73892 75964
rect 73948 51238 74004 51248
rect 73948 47818 74004 51182
rect 73948 47752 74004 47762
rect 73836 3714 73892 3724
rect 74172 4004 74228 4014
rect 73612 3602 73668 3612
rect 72044 3378 72100 3388
rect 74172 2884 74228 3948
rect 74508 3780 74564 77756
rect 75404 75908 75460 75918
rect 74508 3714 74564 3724
rect 74732 73556 74788 73566
rect 74732 3220 74788 73500
rect 74732 3154 74788 3164
rect 74844 59518 74900 59528
rect 74172 2818 74228 2828
rect 74844 2772 74900 59462
rect 75292 43858 75348 43868
rect 74844 2706 74900 2716
rect 74956 35758 75012 35768
rect 74956 1652 75012 35702
rect 75180 33958 75236 33968
rect 75068 4564 75124 4574
rect 75068 3220 75124 4508
rect 75180 3780 75236 33902
rect 75180 3714 75236 3724
rect 75292 3668 75348 43802
rect 75404 3780 75460 75852
rect 75516 45658 75572 45668
rect 75516 36298 75572 45602
rect 75516 36232 75572 36242
rect 75404 3714 75460 3724
rect 75852 3780 75908 79548
rect 76412 65458 76468 416780
rect 84812 79940 84868 79950
rect 76412 65392 76468 65402
rect 76524 79716 76580 79726
rect 76412 62578 76468 62588
rect 75852 3714 75908 3724
rect 76076 42238 76132 42248
rect 76076 3780 76132 42182
rect 76412 13438 76468 62522
rect 76412 13372 76468 13382
rect 76524 4564 76580 79660
rect 81564 79492 81620 79502
rect 78316 79380 78372 79390
rect 76636 78036 76692 78046
rect 76636 25138 76692 77980
rect 76636 25072 76692 25082
rect 77084 74116 77140 74126
rect 76860 24058 76916 24068
rect 76524 4498 76580 4508
rect 76748 19378 76804 19388
rect 76076 3714 76132 3724
rect 75292 3602 75348 3612
rect 76748 3668 76804 19322
rect 76748 3602 76804 3612
rect 75068 3154 75124 3164
rect 76860 3108 76916 24002
rect 76972 21718 77028 21728
rect 76972 3780 77028 21662
rect 76972 3714 77028 3724
rect 77084 3556 77140 74060
rect 77888 58350 78208 58384
rect 77888 58294 77958 58350
rect 78014 58294 78082 58350
rect 78138 58294 78208 58350
rect 77888 58226 78208 58294
rect 77888 58170 77958 58226
rect 78014 58170 78082 58226
rect 78138 58170 78208 58226
rect 77888 58102 78208 58170
rect 77888 58046 77958 58102
rect 78014 58046 78082 58102
rect 78138 58046 78208 58102
rect 77888 57978 78208 58046
rect 77888 57922 77958 57978
rect 78014 57922 78082 57978
rect 78138 57922 78208 57978
rect 77888 57888 78208 57922
rect 77888 40350 78208 40384
rect 77888 40294 77958 40350
rect 78014 40294 78082 40350
rect 78138 40294 78208 40350
rect 77888 40226 78208 40294
rect 77888 40170 77958 40226
rect 78014 40170 78082 40226
rect 78138 40170 78208 40226
rect 77888 40102 78208 40170
rect 77888 40046 77958 40102
rect 78014 40046 78082 40102
rect 78138 40046 78208 40102
rect 77888 39978 78208 40046
rect 77888 39922 77958 39978
rect 78014 39922 78082 39978
rect 78138 39922 78208 39978
rect 77888 39888 78208 39922
rect 77644 25138 77700 25148
rect 77084 3490 77140 3500
rect 77308 9118 77364 9128
rect 76860 3042 76916 3052
rect 74956 1586 75012 1596
rect 76300 1652 76356 1662
rect 76300 1558 76356 1596
rect 76300 1492 76356 1502
rect 77308 1428 77364 9062
rect 77644 3780 77700 25082
rect 77888 22350 78208 22384
rect 77888 22294 77958 22350
rect 78014 22294 78082 22350
rect 78138 22294 78208 22350
rect 77888 22226 78208 22294
rect 77888 22170 77958 22226
rect 78014 22170 78082 22226
rect 78138 22170 78208 22226
rect 77888 22102 78208 22170
rect 77888 22046 77958 22102
rect 78014 22046 78082 22102
rect 78138 22046 78208 22102
rect 77888 21978 78208 22046
rect 77888 21922 77958 21978
rect 78014 21922 78082 21978
rect 78138 21922 78208 21978
rect 77888 21888 78208 21922
rect 78316 21718 78372 79324
rect 78876 79268 78932 79278
rect 78428 64738 78484 64748
rect 78428 51418 78484 64682
rect 78428 51352 78484 51362
rect 78540 55018 78596 55028
rect 78316 21652 78372 21662
rect 78428 48718 78484 48728
rect 77644 3714 77700 3724
rect 77980 5338 78036 5348
rect 77980 2660 78036 5282
rect 78428 3220 78484 48662
rect 78428 3154 78484 3164
rect 77980 2594 78036 2604
rect 77308 1362 77364 1372
rect 78540 532 78596 54962
rect 78652 20278 78708 20288
rect 78652 2548 78708 20222
rect 78876 3780 78932 79212
rect 78876 3714 78932 3724
rect 79436 77700 79492 77710
rect 79436 3780 79492 77644
rect 81452 75796 81508 75806
rect 80108 72658 80164 72668
rect 79884 60418 79940 60428
rect 79772 53038 79828 53048
rect 79772 15148 79828 52982
rect 79884 44758 79940 60362
rect 79884 44692 79940 44702
rect 79996 55918 80052 55928
rect 79660 15092 79828 15148
rect 79884 37198 79940 37208
rect 79548 4564 79604 4574
rect 79548 4004 79604 4508
rect 79548 3938 79604 3948
rect 79436 3714 79492 3724
rect 78652 2482 78708 2492
rect 79660 1316 79716 15092
rect 79772 4228 79828 4238
rect 79772 2884 79828 4172
rect 79884 3556 79940 37142
rect 79996 25138 80052 55862
rect 79996 25072 80052 25082
rect 79996 12178 80052 12188
rect 79996 3892 80052 12122
rect 79996 3826 80052 3836
rect 80108 3668 80164 72602
rect 81228 65818 81284 65828
rect 80556 61318 80612 61328
rect 80556 59878 80612 61262
rect 80556 59812 80612 59822
rect 80556 34318 80612 34328
rect 80556 32698 80612 34262
rect 80556 32632 80612 32642
rect 80780 33778 80836 33788
rect 80556 26218 80612 26228
rect 80108 3602 80164 3612
rect 80444 23878 80500 23888
rect 79884 3490 79940 3500
rect 79772 2818 79828 2828
rect 80444 2772 80500 23822
rect 80556 3780 80612 26162
rect 80668 4564 80724 4574
rect 80668 3892 80724 4508
rect 80668 3826 80724 3836
rect 80556 3714 80612 3724
rect 80780 3780 80836 33722
rect 80780 3714 80836 3724
rect 81228 3780 81284 65762
rect 81228 3714 81284 3724
rect 81452 3556 81508 75740
rect 81564 48718 81620 79436
rect 81564 48652 81620 48662
rect 81788 79156 81844 79166
rect 81676 44038 81732 44048
rect 81452 3490 81508 3500
rect 81564 41338 81620 41348
rect 80444 2706 80500 2716
rect 79660 1250 79716 1260
rect 80556 1764 80612 1774
rect 80108 1204 80164 1214
rect 80108 868 80164 1148
rect 80556 1092 80612 1708
rect 81564 1558 81620 41282
rect 81676 33958 81732 43982
rect 81676 33892 81732 33902
rect 81676 23698 81732 23708
rect 81676 3332 81732 23642
rect 81788 20188 81844 79100
rect 83020 77588 83076 77598
rect 82572 74900 82628 74910
rect 81788 20132 82068 20188
rect 81900 6778 81956 6788
rect 81900 3668 81956 6722
rect 82012 3780 82068 20132
rect 82012 3714 82068 3724
rect 82124 4228 82180 4238
rect 81900 3602 81956 3612
rect 82124 3668 82180 4172
rect 82572 3780 82628 74844
rect 82572 3714 82628 3724
rect 82796 32698 82852 32708
rect 82796 3780 82852 32642
rect 82796 3714 82852 3724
rect 82908 5518 82964 5528
rect 82124 3602 82180 3612
rect 82908 3668 82964 5462
rect 83020 3780 83076 77532
rect 84588 72478 84644 72488
rect 83132 69238 83188 69248
rect 83132 55018 83188 69182
rect 83356 67798 83412 67808
rect 83132 54952 83188 54962
rect 83244 60958 83300 60968
rect 83020 3714 83076 3724
rect 83132 44398 83188 44408
rect 82908 3602 82964 3612
rect 83132 3388 83188 44342
rect 83244 26218 83300 60902
rect 83356 54838 83412 67742
rect 83356 54772 83412 54782
rect 84140 67438 84196 67448
rect 83804 35578 83860 35588
rect 83244 26152 83300 26162
rect 83692 28918 83748 28928
rect 81676 3266 81732 3276
rect 83020 3332 83188 3388
rect 83244 12358 83300 12368
rect 81564 1492 81620 1502
rect 81788 1558 81844 1568
rect 81788 1316 81844 1502
rect 81788 1250 81844 1260
rect 80556 1026 80612 1036
rect 80108 802 80164 812
rect 83020 868 83076 3332
rect 83244 1652 83300 12302
rect 83580 8578 83636 8588
rect 83580 2884 83636 8522
rect 83692 3780 83748 28862
rect 83692 3714 83748 3724
rect 83804 3668 83860 35522
rect 84140 3780 84196 67382
rect 84140 3714 84196 3724
rect 84588 3780 84644 72422
rect 84700 64918 84756 64928
rect 84700 60058 84756 64862
rect 84700 59992 84756 60002
rect 84588 3714 84644 3724
rect 84700 4340 84756 4350
rect 83804 3602 83860 3612
rect 83580 2818 83636 2828
rect 83244 1586 83300 1596
rect 83020 802 83076 812
rect 84700 756 84756 4284
rect 84812 3556 84868 79884
rect 85932 79318 85988 79328
rect 85596 77476 85652 77486
rect 84924 65998 84980 66008
rect 84924 51598 84980 65942
rect 84924 51532 84980 51542
rect 85484 51058 85540 51068
rect 84812 3490 84868 3500
rect 84924 37018 84980 37028
rect 84700 690 84756 700
rect 78540 466 78596 476
rect 84924 308 84980 36962
rect 85036 25498 85092 25508
rect 85036 2996 85092 25442
rect 85484 15148 85540 51002
rect 85372 15092 85540 15148
rect 85372 3668 85428 15092
rect 85596 3898 85652 77420
rect 85484 3842 85652 3898
rect 85708 4564 85764 4574
rect 85484 3780 85540 3842
rect 85484 3714 85540 3724
rect 85372 3602 85428 3612
rect 85036 2930 85092 2940
rect 85708 1018 85764 4508
rect 85932 3780 85988 79262
rect 86492 63658 86548 443212
rect 97578 436350 98198 453922
rect 97578 436294 97674 436350
rect 97730 436294 97798 436350
rect 97854 436294 97922 436350
rect 97978 436294 98046 436350
rect 98102 436294 98198 436350
rect 97578 436226 98198 436294
rect 97578 436170 97674 436226
rect 97730 436170 97798 436226
rect 97854 436170 97922 436226
rect 97978 436170 98046 436226
rect 98102 436170 98198 436226
rect 97578 436102 98198 436170
rect 97578 436046 97674 436102
rect 97730 436046 97798 436102
rect 97854 436046 97922 436102
rect 97978 436046 98046 436102
rect 98102 436046 98198 436102
rect 97578 435978 98198 436046
rect 97578 435922 97674 435978
rect 97730 435922 97798 435978
rect 97854 435922 97922 435978
rect 97978 435922 98046 435978
rect 98102 435922 98198 435978
rect 97578 418350 98198 435922
rect 97578 418294 97674 418350
rect 97730 418294 97798 418350
rect 97854 418294 97922 418350
rect 97978 418294 98046 418350
rect 98102 418294 98198 418350
rect 97578 418226 98198 418294
rect 97578 418170 97674 418226
rect 97730 418170 97798 418226
rect 97854 418170 97922 418226
rect 97978 418170 98046 418226
rect 98102 418170 98198 418226
rect 97578 418102 98198 418170
rect 97578 418046 97674 418102
rect 97730 418046 97798 418102
rect 97854 418046 97922 418102
rect 97978 418046 98046 418102
rect 98102 418046 98198 418102
rect 97578 417978 98198 418046
rect 97578 417922 97674 417978
rect 97730 417922 97798 417978
rect 97854 417922 97922 417978
rect 97978 417922 98046 417978
rect 98102 417922 98198 417978
rect 97578 400350 98198 417922
rect 97578 400294 97674 400350
rect 97730 400294 97798 400350
rect 97854 400294 97922 400350
rect 97978 400294 98046 400350
rect 98102 400294 98198 400350
rect 97578 400226 98198 400294
rect 97578 400170 97674 400226
rect 97730 400170 97798 400226
rect 97854 400170 97922 400226
rect 97978 400170 98046 400226
rect 98102 400170 98198 400226
rect 97578 400102 98198 400170
rect 97578 400046 97674 400102
rect 97730 400046 97798 400102
rect 97854 400046 97922 400102
rect 97978 400046 98046 400102
rect 98102 400046 98198 400102
rect 97578 399978 98198 400046
rect 97578 399922 97674 399978
rect 97730 399922 97798 399978
rect 97854 399922 97922 399978
rect 97978 399922 98046 399978
rect 98102 399922 98198 399978
rect 97578 382350 98198 399922
rect 97578 382294 97674 382350
rect 97730 382294 97798 382350
rect 97854 382294 97922 382350
rect 97978 382294 98046 382350
rect 98102 382294 98198 382350
rect 97578 382226 98198 382294
rect 97578 382170 97674 382226
rect 97730 382170 97798 382226
rect 97854 382170 97922 382226
rect 97978 382170 98046 382226
rect 98102 382170 98198 382226
rect 97578 382102 98198 382170
rect 97578 382046 97674 382102
rect 97730 382046 97798 382102
rect 97854 382046 97922 382102
rect 97978 382046 98046 382102
rect 98102 382046 98198 382102
rect 97578 381978 98198 382046
rect 97578 381922 97674 381978
rect 97730 381922 97798 381978
rect 97854 381922 97922 381978
rect 97978 381922 98046 381978
rect 98102 381922 98198 381978
rect 97578 364350 98198 381922
rect 97578 364294 97674 364350
rect 97730 364294 97798 364350
rect 97854 364294 97922 364350
rect 97978 364294 98046 364350
rect 98102 364294 98198 364350
rect 97578 364226 98198 364294
rect 97578 364170 97674 364226
rect 97730 364170 97798 364226
rect 97854 364170 97922 364226
rect 97978 364170 98046 364226
rect 98102 364170 98198 364226
rect 97578 364102 98198 364170
rect 97578 364046 97674 364102
rect 97730 364046 97798 364102
rect 97854 364046 97922 364102
rect 97978 364046 98046 364102
rect 98102 364046 98198 364102
rect 97578 363978 98198 364046
rect 97578 363922 97674 363978
rect 97730 363922 97798 363978
rect 97854 363922 97922 363978
rect 97978 363922 98046 363978
rect 98102 363922 98198 363978
rect 97578 346350 98198 363922
rect 97578 346294 97674 346350
rect 97730 346294 97798 346350
rect 97854 346294 97922 346350
rect 97978 346294 98046 346350
rect 98102 346294 98198 346350
rect 97578 346226 98198 346294
rect 97578 346170 97674 346226
rect 97730 346170 97798 346226
rect 97854 346170 97922 346226
rect 97978 346170 98046 346226
rect 98102 346170 98198 346226
rect 97578 346102 98198 346170
rect 97578 346046 97674 346102
rect 97730 346046 97798 346102
rect 97854 346046 97922 346102
rect 97978 346046 98046 346102
rect 98102 346046 98198 346102
rect 97578 345978 98198 346046
rect 97578 345922 97674 345978
rect 97730 345922 97798 345978
rect 97854 345922 97922 345978
rect 97978 345922 98046 345978
rect 98102 345922 98198 345978
rect 97578 328350 98198 345922
rect 97578 328294 97674 328350
rect 97730 328294 97798 328350
rect 97854 328294 97922 328350
rect 97978 328294 98046 328350
rect 98102 328294 98198 328350
rect 97578 328226 98198 328294
rect 97578 328170 97674 328226
rect 97730 328170 97798 328226
rect 97854 328170 97922 328226
rect 97978 328170 98046 328226
rect 98102 328170 98198 328226
rect 97578 328102 98198 328170
rect 97578 328046 97674 328102
rect 97730 328046 97798 328102
rect 97854 328046 97922 328102
rect 97978 328046 98046 328102
rect 98102 328046 98198 328102
rect 97578 327978 98198 328046
rect 97578 327922 97674 327978
rect 97730 327922 97798 327978
rect 97854 327922 97922 327978
rect 97978 327922 98046 327978
rect 98102 327922 98198 327978
rect 97578 310350 98198 327922
rect 97578 310294 97674 310350
rect 97730 310294 97798 310350
rect 97854 310294 97922 310350
rect 97978 310294 98046 310350
rect 98102 310294 98198 310350
rect 97578 310226 98198 310294
rect 97578 310170 97674 310226
rect 97730 310170 97798 310226
rect 97854 310170 97922 310226
rect 97978 310170 98046 310226
rect 98102 310170 98198 310226
rect 97578 310102 98198 310170
rect 97578 310046 97674 310102
rect 97730 310046 97798 310102
rect 97854 310046 97922 310102
rect 97978 310046 98046 310102
rect 98102 310046 98198 310102
rect 97578 309978 98198 310046
rect 97578 309922 97674 309978
rect 97730 309922 97798 309978
rect 97854 309922 97922 309978
rect 97978 309922 98046 309978
rect 98102 309922 98198 309978
rect 97578 292350 98198 309922
rect 97578 292294 97674 292350
rect 97730 292294 97798 292350
rect 97854 292294 97922 292350
rect 97978 292294 98046 292350
rect 98102 292294 98198 292350
rect 97578 292226 98198 292294
rect 97578 292170 97674 292226
rect 97730 292170 97798 292226
rect 97854 292170 97922 292226
rect 97978 292170 98046 292226
rect 98102 292170 98198 292226
rect 97578 292102 98198 292170
rect 97578 292046 97674 292102
rect 97730 292046 97798 292102
rect 97854 292046 97922 292102
rect 97978 292046 98046 292102
rect 98102 292046 98198 292102
rect 97578 291978 98198 292046
rect 97578 291922 97674 291978
rect 97730 291922 97798 291978
rect 97854 291922 97922 291978
rect 97978 291922 98046 291978
rect 98102 291922 98198 291978
rect 97578 274350 98198 291922
rect 97578 274294 97674 274350
rect 97730 274294 97798 274350
rect 97854 274294 97922 274350
rect 97978 274294 98046 274350
rect 98102 274294 98198 274350
rect 97578 274226 98198 274294
rect 97578 274170 97674 274226
rect 97730 274170 97798 274226
rect 97854 274170 97922 274226
rect 97978 274170 98046 274226
rect 98102 274170 98198 274226
rect 97578 274102 98198 274170
rect 97578 274046 97674 274102
rect 97730 274046 97798 274102
rect 97854 274046 97922 274102
rect 97978 274046 98046 274102
rect 98102 274046 98198 274102
rect 97578 273978 98198 274046
rect 97578 273922 97674 273978
rect 97730 273922 97798 273978
rect 97854 273922 97922 273978
rect 97978 273922 98046 273978
rect 98102 273922 98198 273978
rect 97578 256350 98198 273922
rect 97578 256294 97674 256350
rect 97730 256294 97798 256350
rect 97854 256294 97922 256350
rect 97978 256294 98046 256350
rect 98102 256294 98198 256350
rect 97578 256226 98198 256294
rect 97578 256170 97674 256226
rect 97730 256170 97798 256226
rect 97854 256170 97922 256226
rect 97978 256170 98046 256226
rect 98102 256170 98198 256226
rect 97578 256102 98198 256170
rect 97578 256046 97674 256102
rect 97730 256046 97798 256102
rect 97854 256046 97922 256102
rect 97978 256046 98046 256102
rect 98102 256046 98198 256102
rect 97578 255978 98198 256046
rect 97578 255922 97674 255978
rect 97730 255922 97798 255978
rect 97854 255922 97922 255978
rect 97978 255922 98046 255978
rect 98102 255922 98198 255978
rect 97578 238350 98198 255922
rect 97578 238294 97674 238350
rect 97730 238294 97798 238350
rect 97854 238294 97922 238350
rect 97978 238294 98046 238350
rect 98102 238294 98198 238350
rect 97578 238226 98198 238294
rect 97578 238170 97674 238226
rect 97730 238170 97798 238226
rect 97854 238170 97922 238226
rect 97978 238170 98046 238226
rect 98102 238170 98198 238226
rect 97578 238102 98198 238170
rect 97578 238046 97674 238102
rect 97730 238046 97798 238102
rect 97854 238046 97922 238102
rect 97978 238046 98046 238102
rect 98102 238046 98198 238102
rect 97578 237978 98198 238046
rect 97578 237922 97674 237978
rect 97730 237922 97798 237978
rect 97854 237922 97922 237978
rect 97978 237922 98046 237978
rect 98102 237922 98198 237978
rect 97578 220350 98198 237922
rect 97578 220294 97674 220350
rect 97730 220294 97798 220350
rect 97854 220294 97922 220350
rect 97978 220294 98046 220350
rect 98102 220294 98198 220350
rect 97578 220226 98198 220294
rect 97578 220170 97674 220226
rect 97730 220170 97798 220226
rect 97854 220170 97922 220226
rect 97978 220170 98046 220226
rect 98102 220170 98198 220226
rect 97578 220102 98198 220170
rect 97578 220046 97674 220102
rect 97730 220046 97798 220102
rect 97854 220046 97922 220102
rect 97978 220046 98046 220102
rect 98102 220046 98198 220102
rect 97578 219978 98198 220046
rect 97578 219922 97674 219978
rect 97730 219922 97798 219978
rect 97854 219922 97922 219978
rect 97978 219922 98046 219978
rect 98102 219922 98198 219978
rect 97578 202350 98198 219922
rect 97578 202294 97674 202350
rect 97730 202294 97798 202350
rect 97854 202294 97922 202350
rect 97978 202294 98046 202350
rect 98102 202294 98198 202350
rect 97578 202226 98198 202294
rect 97578 202170 97674 202226
rect 97730 202170 97798 202226
rect 97854 202170 97922 202226
rect 97978 202170 98046 202226
rect 98102 202170 98198 202226
rect 97578 202102 98198 202170
rect 97578 202046 97674 202102
rect 97730 202046 97798 202102
rect 97854 202046 97922 202102
rect 97978 202046 98046 202102
rect 98102 202046 98198 202102
rect 97578 201978 98198 202046
rect 97578 201922 97674 201978
rect 97730 201922 97798 201978
rect 97854 201922 97922 201978
rect 97978 201922 98046 201978
rect 98102 201922 98198 201978
rect 97578 184350 98198 201922
rect 97578 184294 97674 184350
rect 97730 184294 97798 184350
rect 97854 184294 97922 184350
rect 97978 184294 98046 184350
rect 98102 184294 98198 184350
rect 97578 184226 98198 184294
rect 97578 184170 97674 184226
rect 97730 184170 97798 184226
rect 97854 184170 97922 184226
rect 97978 184170 98046 184226
rect 98102 184170 98198 184226
rect 97578 184102 98198 184170
rect 97578 184046 97674 184102
rect 97730 184046 97798 184102
rect 97854 184046 97922 184102
rect 97978 184046 98046 184102
rect 98102 184046 98198 184102
rect 97578 183978 98198 184046
rect 97578 183922 97674 183978
rect 97730 183922 97798 183978
rect 97854 183922 97922 183978
rect 97978 183922 98046 183978
rect 98102 183922 98198 183978
rect 97578 166350 98198 183922
rect 97578 166294 97674 166350
rect 97730 166294 97798 166350
rect 97854 166294 97922 166350
rect 97978 166294 98046 166350
rect 98102 166294 98198 166350
rect 97578 166226 98198 166294
rect 97578 166170 97674 166226
rect 97730 166170 97798 166226
rect 97854 166170 97922 166226
rect 97978 166170 98046 166226
rect 98102 166170 98198 166226
rect 97578 166102 98198 166170
rect 97578 166046 97674 166102
rect 97730 166046 97798 166102
rect 97854 166046 97922 166102
rect 97978 166046 98046 166102
rect 98102 166046 98198 166102
rect 97578 165978 98198 166046
rect 97578 165922 97674 165978
rect 97730 165922 97798 165978
rect 97854 165922 97922 165978
rect 97978 165922 98046 165978
rect 98102 165922 98198 165978
rect 97578 148350 98198 165922
rect 97578 148294 97674 148350
rect 97730 148294 97798 148350
rect 97854 148294 97922 148350
rect 97978 148294 98046 148350
rect 98102 148294 98198 148350
rect 97578 148226 98198 148294
rect 97578 148170 97674 148226
rect 97730 148170 97798 148226
rect 97854 148170 97922 148226
rect 97978 148170 98046 148226
rect 98102 148170 98198 148226
rect 97578 148102 98198 148170
rect 97578 148046 97674 148102
rect 97730 148046 97798 148102
rect 97854 148046 97922 148102
rect 97978 148046 98046 148102
rect 98102 148046 98198 148102
rect 97578 147978 98198 148046
rect 97578 147922 97674 147978
rect 97730 147922 97798 147978
rect 97854 147922 97922 147978
rect 97978 147922 98046 147978
rect 98102 147922 98198 147978
rect 97578 130350 98198 147922
rect 97578 130294 97674 130350
rect 97730 130294 97798 130350
rect 97854 130294 97922 130350
rect 97978 130294 98046 130350
rect 98102 130294 98198 130350
rect 97578 130226 98198 130294
rect 97578 130170 97674 130226
rect 97730 130170 97798 130226
rect 97854 130170 97922 130226
rect 97978 130170 98046 130226
rect 98102 130170 98198 130226
rect 97578 130102 98198 130170
rect 97578 130046 97674 130102
rect 97730 130046 97798 130102
rect 97854 130046 97922 130102
rect 97978 130046 98046 130102
rect 98102 130046 98198 130102
rect 97578 129978 98198 130046
rect 97578 129922 97674 129978
rect 97730 129922 97798 129978
rect 97854 129922 97922 129978
rect 97978 129922 98046 129978
rect 98102 129922 98198 129978
rect 97578 112350 98198 129922
rect 97578 112294 97674 112350
rect 97730 112294 97798 112350
rect 97854 112294 97922 112350
rect 97978 112294 98046 112350
rect 98102 112294 98198 112350
rect 97578 112226 98198 112294
rect 97578 112170 97674 112226
rect 97730 112170 97798 112226
rect 97854 112170 97922 112226
rect 97978 112170 98046 112226
rect 98102 112170 98198 112226
rect 97578 112102 98198 112170
rect 97578 112046 97674 112102
rect 97730 112046 97798 112102
rect 97854 112046 97922 112102
rect 97978 112046 98046 112102
rect 98102 112046 98198 112102
rect 97578 111978 98198 112046
rect 97578 111922 97674 111978
rect 97730 111922 97798 111978
rect 97854 111922 97922 111978
rect 97978 111922 98046 111978
rect 98102 111922 98198 111978
rect 97578 94350 98198 111922
rect 97578 94294 97674 94350
rect 97730 94294 97798 94350
rect 97854 94294 97922 94350
rect 97978 94294 98046 94350
rect 98102 94294 98198 94350
rect 97578 94226 98198 94294
rect 97578 94170 97674 94226
rect 97730 94170 97798 94226
rect 97854 94170 97922 94226
rect 97978 94170 98046 94226
rect 98102 94170 98198 94226
rect 97578 94102 98198 94170
rect 97578 94046 97674 94102
rect 97730 94046 97798 94102
rect 97854 94046 97922 94102
rect 97978 94046 98046 94102
rect 98102 94046 98198 94102
rect 97578 93978 98198 94046
rect 97578 93922 97674 93978
rect 97730 93922 97798 93978
rect 97854 93922 97922 93978
rect 97978 93922 98046 93978
rect 98102 93922 98198 93978
rect 89740 79138 89796 79148
rect 86492 63592 86548 63602
rect 86604 78372 86660 78382
rect 85932 3714 85988 3724
rect 86156 47458 86212 47468
rect 86156 3780 86212 47402
rect 86156 3714 86212 3724
rect 86604 3332 86660 78316
rect 87948 76580 88004 76590
rect 87276 74098 87332 74108
rect 87164 59338 87220 59348
rect 87052 54478 87108 54488
rect 86940 22618 86996 22628
rect 86940 15148 86996 22562
rect 86716 15092 86996 15148
rect 86716 3444 86772 15092
rect 87052 5158 87108 54422
rect 86828 5102 87108 5158
rect 86828 3780 86884 5102
rect 86828 3714 86884 3724
rect 87164 3780 87220 59282
rect 87276 3892 87332 74042
rect 87388 66178 87444 66188
rect 87388 62938 87444 66122
rect 87388 62872 87444 62882
rect 87836 28738 87892 28748
rect 87836 25498 87892 28682
rect 87836 25432 87892 25442
rect 87500 16858 87556 16868
rect 87276 3826 87332 3836
rect 87388 6058 87444 6068
rect 87164 3714 87220 3724
rect 86716 3378 86772 3388
rect 86604 3266 86660 3276
rect 85932 1764 85988 1774
rect 85932 1540 85988 1708
rect 85932 1474 85988 1484
rect 87388 1378 87444 6002
rect 87500 2884 87556 16802
rect 87836 11818 87892 11828
rect 87724 11762 87836 11818
rect 87724 3780 87780 11762
rect 87836 11752 87892 11762
rect 87724 3714 87780 3724
rect 87948 3780 88004 76524
rect 88956 72298 89012 72308
rect 88284 71038 88340 71048
rect 88284 49618 88340 70982
rect 88844 62398 88900 62408
rect 88284 49552 88340 49562
rect 88732 52498 88788 52508
rect 87948 3714 88004 3724
rect 88172 49078 88228 49088
rect 87500 2818 87556 2828
rect 88172 1652 88228 49022
rect 88732 3444 88788 52442
rect 88844 3780 88900 62342
rect 88956 3892 89012 72242
rect 89516 59158 89572 59168
rect 89292 50878 89348 50888
rect 88956 3826 89012 3836
rect 89068 13618 89124 13628
rect 88844 3714 88900 3724
rect 89068 3780 89124 13562
rect 89068 3714 89124 3724
rect 89292 3780 89348 50822
rect 89292 3714 89348 3724
rect 89516 3780 89572 59102
rect 89516 3714 89572 3724
rect 89740 3780 89796 79082
rect 92316 77338 92372 77348
rect 91532 74004 91588 74014
rect 89852 71218 89908 71228
rect 89852 60418 89908 71162
rect 89852 60352 89908 60362
rect 90636 60778 90692 60788
rect 90412 54298 90468 54308
rect 89852 25678 89908 25688
rect 89852 19378 89908 25622
rect 89852 19312 89908 19322
rect 89740 3714 89796 3724
rect 89852 17038 89908 17048
rect 88732 3378 88788 3388
rect 89404 2818 89460 2828
rect 89404 1764 89460 2762
rect 89404 1698 89460 1708
rect 88172 1586 88228 1596
rect 89852 1558 89908 16982
rect 90412 3780 90468 54242
rect 90412 3714 90468 3724
rect 90636 3444 90692 60722
rect 90860 47278 90916 47288
rect 90748 45478 90804 45488
rect 90748 42778 90804 45422
rect 90748 42712 90804 42722
rect 90748 34138 90804 34148
rect 90748 28738 90804 34082
rect 90748 28672 90804 28682
rect 90636 3378 90692 3388
rect 90748 8578 90804 8588
rect 90748 1652 90804 8522
rect 90860 3780 90916 47222
rect 91308 38818 91364 38828
rect 90860 3714 90916 3724
rect 90972 11098 91028 11108
rect 90748 1586 90804 1596
rect 89852 1492 89908 1502
rect 87276 1322 87444 1378
rect 87276 1316 87332 1322
rect 87276 1250 87332 1260
rect 90972 1092 91028 11042
rect 91308 3780 91364 38762
rect 91420 4340 91476 4350
rect 91420 4004 91476 4284
rect 91420 3938 91476 3948
rect 91308 3714 91364 3724
rect 91532 2660 91588 73948
rect 91644 67978 91700 67988
rect 91644 56278 91700 67922
rect 91644 56212 91700 56222
rect 91756 66358 91812 66368
rect 91644 56098 91700 56108
rect 91644 39538 91700 56042
rect 91756 52858 91812 66302
rect 91756 52792 91812 52802
rect 91644 39472 91700 39482
rect 92204 30358 92260 30368
rect 92092 28738 92148 28748
rect 92092 3780 92148 28682
rect 92092 3714 92148 3724
rect 92204 3332 92260 30302
rect 92316 3444 92372 77282
rect 97578 76350 98198 93922
rect 99148 572852 99316 572908
rect 101298 586350 101918 597744
rect 128298 597212 128918 598268
rect 128298 597156 128394 597212
rect 128450 597156 128518 597212
rect 128574 597156 128642 597212
rect 128698 597156 128766 597212
rect 128822 597156 128918 597212
rect 128298 597088 128918 597156
rect 128298 597032 128394 597088
rect 128450 597032 128518 597088
rect 128574 597032 128642 597088
rect 128698 597032 128766 597088
rect 128822 597032 128918 597088
rect 128298 596964 128918 597032
rect 128298 596908 128394 596964
rect 128450 596908 128518 596964
rect 128574 596908 128642 596964
rect 128698 596908 128766 596964
rect 128822 596908 128918 596964
rect 128298 596840 128918 596908
rect 128298 596784 128394 596840
rect 128450 596784 128518 596840
rect 128574 596784 128642 596840
rect 128698 596784 128766 596840
rect 128822 596784 128918 596840
rect 101298 586294 101394 586350
rect 101450 586294 101518 586350
rect 101574 586294 101642 586350
rect 101698 586294 101766 586350
rect 101822 586294 101918 586350
rect 101298 586226 101918 586294
rect 101298 586170 101394 586226
rect 101450 586170 101518 586226
rect 101574 586170 101642 586226
rect 101698 586170 101766 586226
rect 101822 586170 101918 586226
rect 101298 586102 101918 586170
rect 101298 586046 101394 586102
rect 101450 586046 101518 586102
rect 101574 586046 101642 586102
rect 101698 586046 101766 586102
rect 101822 586046 101918 586102
rect 101298 585978 101918 586046
rect 101298 585922 101394 585978
rect 101450 585922 101518 585978
rect 101574 585922 101642 585978
rect 101698 585922 101766 585978
rect 101822 585922 101918 585978
rect 99148 80038 99204 572852
rect 99148 79972 99204 79982
rect 101298 568350 101918 585922
rect 101298 568294 101394 568350
rect 101450 568294 101518 568350
rect 101574 568294 101642 568350
rect 101698 568294 101766 568350
rect 101822 568294 101918 568350
rect 101298 568226 101918 568294
rect 101298 568170 101394 568226
rect 101450 568170 101518 568226
rect 101574 568170 101642 568226
rect 101698 568170 101766 568226
rect 101822 568170 101918 568226
rect 101298 568102 101918 568170
rect 101298 568046 101394 568102
rect 101450 568046 101518 568102
rect 101574 568046 101642 568102
rect 101698 568046 101766 568102
rect 101822 568046 101918 568102
rect 101298 567978 101918 568046
rect 101298 567922 101394 567978
rect 101450 567922 101518 567978
rect 101574 567922 101642 567978
rect 101698 567922 101766 567978
rect 101822 567922 101918 567978
rect 101298 550350 101918 567922
rect 101298 550294 101394 550350
rect 101450 550294 101518 550350
rect 101574 550294 101642 550350
rect 101698 550294 101766 550350
rect 101822 550294 101918 550350
rect 101298 550226 101918 550294
rect 101298 550170 101394 550226
rect 101450 550170 101518 550226
rect 101574 550170 101642 550226
rect 101698 550170 101766 550226
rect 101822 550170 101918 550226
rect 101298 550102 101918 550170
rect 101298 550046 101394 550102
rect 101450 550046 101518 550102
rect 101574 550046 101642 550102
rect 101698 550046 101766 550102
rect 101822 550046 101918 550102
rect 101298 549978 101918 550046
rect 101298 549922 101394 549978
rect 101450 549922 101518 549978
rect 101574 549922 101642 549978
rect 101698 549922 101766 549978
rect 101822 549922 101918 549978
rect 101298 532350 101918 549922
rect 101298 532294 101394 532350
rect 101450 532294 101518 532350
rect 101574 532294 101642 532350
rect 101698 532294 101766 532350
rect 101822 532294 101918 532350
rect 101298 532226 101918 532294
rect 101298 532170 101394 532226
rect 101450 532170 101518 532226
rect 101574 532170 101642 532226
rect 101698 532170 101766 532226
rect 101822 532170 101918 532226
rect 101298 532102 101918 532170
rect 101298 532046 101394 532102
rect 101450 532046 101518 532102
rect 101574 532046 101642 532102
rect 101698 532046 101766 532102
rect 101822 532046 101918 532102
rect 101298 531978 101918 532046
rect 101298 531922 101394 531978
rect 101450 531922 101518 531978
rect 101574 531922 101642 531978
rect 101698 531922 101766 531978
rect 101822 531922 101918 531978
rect 101298 514350 101918 531922
rect 101298 514294 101394 514350
rect 101450 514294 101518 514350
rect 101574 514294 101642 514350
rect 101698 514294 101766 514350
rect 101822 514294 101918 514350
rect 101298 514226 101918 514294
rect 101298 514170 101394 514226
rect 101450 514170 101518 514226
rect 101574 514170 101642 514226
rect 101698 514170 101766 514226
rect 101822 514170 101918 514226
rect 101298 514102 101918 514170
rect 101298 514046 101394 514102
rect 101450 514046 101518 514102
rect 101574 514046 101642 514102
rect 101698 514046 101766 514102
rect 101822 514046 101918 514102
rect 101298 513978 101918 514046
rect 101298 513922 101394 513978
rect 101450 513922 101518 513978
rect 101574 513922 101642 513978
rect 101698 513922 101766 513978
rect 101822 513922 101918 513978
rect 101298 496350 101918 513922
rect 101298 496294 101394 496350
rect 101450 496294 101518 496350
rect 101574 496294 101642 496350
rect 101698 496294 101766 496350
rect 101822 496294 101918 496350
rect 101298 496226 101918 496294
rect 101298 496170 101394 496226
rect 101450 496170 101518 496226
rect 101574 496170 101642 496226
rect 101698 496170 101766 496226
rect 101822 496170 101918 496226
rect 101298 496102 101918 496170
rect 101298 496046 101394 496102
rect 101450 496046 101518 496102
rect 101574 496046 101642 496102
rect 101698 496046 101766 496102
rect 101822 496046 101918 496102
rect 101298 495978 101918 496046
rect 101298 495922 101394 495978
rect 101450 495922 101518 495978
rect 101574 495922 101642 495978
rect 101698 495922 101766 495978
rect 101822 495922 101918 495978
rect 101298 478350 101918 495922
rect 101298 478294 101394 478350
rect 101450 478294 101518 478350
rect 101574 478294 101642 478350
rect 101698 478294 101766 478350
rect 101822 478294 101918 478350
rect 101298 478226 101918 478294
rect 101298 478170 101394 478226
rect 101450 478170 101518 478226
rect 101574 478170 101642 478226
rect 101698 478170 101766 478226
rect 101822 478170 101918 478226
rect 101298 478102 101918 478170
rect 101298 478046 101394 478102
rect 101450 478046 101518 478102
rect 101574 478046 101642 478102
rect 101698 478046 101766 478102
rect 101822 478046 101918 478102
rect 101298 477978 101918 478046
rect 101298 477922 101394 477978
rect 101450 477922 101518 477978
rect 101574 477922 101642 477978
rect 101698 477922 101766 477978
rect 101822 477922 101918 477978
rect 101298 460350 101918 477922
rect 101298 460294 101394 460350
rect 101450 460294 101518 460350
rect 101574 460294 101642 460350
rect 101698 460294 101766 460350
rect 101822 460294 101918 460350
rect 101298 460226 101918 460294
rect 101298 460170 101394 460226
rect 101450 460170 101518 460226
rect 101574 460170 101642 460226
rect 101698 460170 101766 460226
rect 101822 460170 101918 460226
rect 101298 460102 101918 460170
rect 101298 460046 101394 460102
rect 101450 460046 101518 460102
rect 101574 460046 101642 460102
rect 101698 460046 101766 460102
rect 101822 460046 101918 460102
rect 101298 459978 101918 460046
rect 101298 459922 101394 459978
rect 101450 459922 101518 459978
rect 101574 459922 101642 459978
rect 101698 459922 101766 459978
rect 101822 459922 101918 459978
rect 101298 442350 101918 459922
rect 101298 442294 101394 442350
rect 101450 442294 101518 442350
rect 101574 442294 101642 442350
rect 101698 442294 101766 442350
rect 101822 442294 101918 442350
rect 101298 442226 101918 442294
rect 101298 442170 101394 442226
rect 101450 442170 101518 442226
rect 101574 442170 101642 442226
rect 101698 442170 101766 442226
rect 101822 442170 101918 442226
rect 101298 442102 101918 442170
rect 101298 442046 101394 442102
rect 101450 442046 101518 442102
rect 101574 442046 101642 442102
rect 101698 442046 101766 442102
rect 101822 442046 101918 442102
rect 101298 441978 101918 442046
rect 101298 441922 101394 441978
rect 101450 441922 101518 441978
rect 101574 441922 101642 441978
rect 101698 441922 101766 441978
rect 101822 441922 101918 441978
rect 101298 424350 101918 441922
rect 101298 424294 101394 424350
rect 101450 424294 101518 424350
rect 101574 424294 101642 424350
rect 101698 424294 101766 424350
rect 101822 424294 101918 424350
rect 101298 424226 101918 424294
rect 101298 424170 101394 424226
rect 101450 424170 101518 424226
rect 101574 424170 101642 424226
rect 101698 424170 101766 424226
rect 101822 424170 101918 424226
rect 101298 424102 101918 424170
rect 101298 424046 101394 424102
rect 101450 424046 101518 424102
rect 101574 424046 101642 424102
rect 101698 424046 101766 424102
rect 101822 424046 101918 424102
rect 101298 423978 101918 424046
rect 101298 423922 101394 423978
rect 101450 423922 101518 423978
rect 101574 423922 101642 423978
rect 101698 423922 101766 423978
rect 101822 423922 101918 423978
rect 101298 406350 101918 423922
rect 101298 406294 101394 406350
rect 101450 406294 101518 406350
rect 101574 406294 101642 406350
rect 101698 406294 101766 406350
rect 101822 406294 101918 406350
rect 101298 406226 101918 406294
rect 101298 406170 101394 406226
rect 101450 406170 101518 406226
rect 101574 406170 101642 406226
rect 101698 406170 101766 406226
rect 101822 406170 101918 406226
rect 101298 406102 101918 406170
rect 101298 406046 101394 406102
rect 101450 406046 101518 406102
rect 101574 406046 101642 406102
rect 101698 406046 101766 406102
rect 101822 406046 101918 406102
rect 101298 405978 101918 406046
rect 101298 405922 101394 405978
rect 101450 405922 101518 405978
rect 101574 405922 101642 405978
rect 101698 405922 101766 405978
rect 101822 405922 101918 405978
rect 101298 388350 101918 405922
rect 101298 388294 101394 388350
rect 101450 388294 101518 388350
rect 101574 388294 101642 388350
rect 101698 388294 101766 388350
rect 101822 388294 101918 388350
rect 101298 388226 101918 388294
rect 101298 388170 101394 388226
rect 101450 388170 101518 388226
rect 101574 388170 101642 388226
rect 101698 388170 101766 388226
rect 101822 388170 101918 388226
rect 101298 388102 101918 388170
rect 101298 388046 101394 388102
rect 101450 388046 101518 388102
rect 101574 388046 101642 388102
rect 101698 388046 101766 388102
rect 101822 388046 101918 388102
rect 101298 387978 101918 388046
rect 101298 387922 101394 387978
rect 101450 387922 101518 387978
rect 101574 387922 101642 387978
rect 101698 387922 101766 387978
rect 101822 387922 101918 387978
rect 101298 370350 101918 387922
rect 101298 370294 101394 370350
rect 101450 370294 101518 370350
rect 101574 370294 101642 370350
rect 101698 370294 101766 370350
rect 101822 370294 101918 370350
rect 101298 370226 101918 370294
rect 101298 370170 101394 370226
rect 101450 370170 101518 370226
rect 101574 370170 101642 370226
rect 101698 370170 101766 370226
rect 101822 370170 101918 370226
rect 101298 370102 101918 370170
rect 101298 370046 101394 370102
rect 101450 370046 101518 370102
rect 101574 370046 101642 370102
rect 101698 370046 101766 370102
rect 101822 370046 101918 370102
rect 101298 369978 101918 370046
rect 101298 369922 101394 369978
rect 101450 369922 101518 369978
rect 101574 369922 101642 369978
rect 101698 369922 101766 369978
rect 101822 369922 101918 369978
rect 101298 352350 101918 369922
rect 101298 352294 101394 352350
rect 101450 352294 101518 352350
rect 101574 352294 101642 352350
rect 101698 352294 101766 352350
rect 101822 352294 101918 352350
rect 101298 352226 101918 352294
rect 101298 352170 101394 352226
rect 101450 352170 101518 352226
rect 101574 352170 101642 352226
rect 101698 352170 101766 352226
rect 101822 352170 101918 352226
rect 101298 352102 101918 352170
rect 101298 352046 101394 352102
rect 101450 352046 101518 352102
rect 101574 352046 101642 352102
rect 101698 352046 101766 352102
rect 101822 352046 101918 352102
rect 101298 351978 101918 352046
rect 101298 351922 101394 351978
rect 101450 351922 101518 351978
rect 101574 351922 101642 351978
rect 101698 351922 101766 351978
rect 101822 351922 101918 351978
rect 101298 334350 101918 351922
rect 101298 334294 101394 334350
rect 101450 334294 101518 334350
rect 101574 334294 101642 334350
rect 101698 334294 101766 334350
rect 101822 334294 101918 334350
rect 101298 334226 101918 334294
rect 101298 334170 101394 334226
rect 101450 334170 101518 334226
rect 101574 334170 101642 334226
rect 101698 334170 101766 334226
rect 101822 334170 101918 334226
rect 101298 334102 101918 334170
rect 101298 334046 101394 334102
rect 101450 334046 101518 334102
rect 101574 334046 101642 334102
rect 101698 334046 101766 334102
rect 101822 334046 101918 334102
rect 101298 333978 101918 334046
rect 101298 333922 101394 333978
rect 101450 333922 101518 333978
rect 101574 333922 101642 333978
rect 101698 333922 101766 333978
rect 101822 333922 101918 333978
rect 101298 316350 101918 333922
rect 101298 316294 101394 316350
rect 101450 316294 101518 316350
rect 101574 316294 101642 316350
rect 101698 316294 101766 316350
rect 101822 316294 101918 316350
rect 101298 316226 101918 316294
rect 101298 316170 101394 316226
rect 101450 316170 101518 316226
rect 101574 316170 101642 316226
rect 101698 316170 101766 316226
rect 101822 316170 101918 316226
rect 101298 316102 101918 316170
rect 101298 316046 101394 316102
rect 101450 316046 101518 316102
rect 101574 316046 101642 316102
rect 101698 316046 101766 316102
rect 101822 316046 101918 316102
rect 101298 315978 101918 316046
rect 101298 315922 101394 315978
rect 101450 315922 101518 315978
rect 101574 315922 101642 315978
rect 101698 315922 101766 315978
rect 101822 315922 101918 315978
rect 101298 298350 101918 315922
rect 101298 298294 101394 298350
rect 101450 298294 101518 298350
rect 101574 298294 101642 298350
rect 101698 298294 101766 298350
rect 101822 298294 101918 298350
rect 101298 298226 101918 298294
rect 101298 298170 101394 298226
rect 101450 298170 101518 298226
rect 101574 298170 101642 298226
rect 101698 298170 101766 298226
rect 101822 298170 101918 298226
rect 101298 298102 101918 298170
rect 101298 298046 101394 298102
rect 101450 298046 101518 298102
rect 101574 298046 101642 298102
rect 101698 298046 101766 298102
rect 101822 298046 101918 298102
rect 101298 297978 101918 298046
rect 101298 297922 101394 297978
rect 101450 297922 101518 297978
rect 101574 297922 101642 297978
rect 101698 297922 101766 297978
rect 101822 297922 101918 297978
rect 101298 280350 101918 297922
rect 101298 280294 101394 280350
rect 101450 280294 101518 280350
rect 101574 280294 101642 280350
rect 101698 280294 101766 280350
rect 101822 280294 101918 280350
rect 101298 280226 101918 280294
rect 101298 280170 101394 280226
rect 101450 280170 101518 280226
rect 101574 280170 101642 280226
rect 101698 280170 101766 280226
rect 101822 280170 101918 280226
rect 101298 280102 101918 280170
rect 101298 280046 101394 280102
rect 101450 280046 101518 280102
rect 101574 280046 101642 280102
rect 101698 280046 101766 280102
rect 101822 280046 101918 280102
rect 101298 279978 101918 280046
rect 101298 279922 101394 279978
rect 101450 279922 101518 279978
rect 101574 279922 101642 279978
rect 101698 279922 101766 279978
rect 101822 279922 101918 279978
rect 101298 262350 101918 279922
rect 101298 262294 101394 262350
rect 101450 262294 101518 262350
rect 101574 262294 101642 262350
rect 101698 262294 101766 262350
rect 101822 262294 101918 262350
rect 101298 262226 101918 262294
rect 101298 262170 101394 262226
rect 101450 262170 101518 262226
rect 101574 262170 101642 262226
rect 101698 262170 101766 262226
rect 101822 262170 101918 262226
rect 101298 262102 101918 262170
rect 101298 262046 101394 262102
rect 101450 262046 101518 262102
rect 101574 262046 101642 262102
rect 101698 262046 101766 262102
rect 101822 262046 101918 262102
rect 101298 261978 101918 262046
rect 101298 261922 101394 261978
rect 101450 261922 101518 261978
rect 101574 261922 101642 261978
rect 101698 261922 101766 261978
rect 101822 261922 101918 261978
rect 101298 244350 101918 261922
rect 101298 244294 101394 244350
rect 101450 244294 101518 244350
rect 101574 244294 101642 244350
rect 101698 244294 101766 244350
rect 101822 244294 101918 244350
rect 101298 244226 101918 244294
rect 101298 244170 101394 244226
rect 101450 244170 101518 244226
rect 101574 244170 101642 244226
rect 101698 244170 101766 244226
rect 101822 244170 101918 244226
rect 101298 244102 101918 244170
rect 101298 244046 101394 244102
rect 101450 244046 101518 244102
rect 101574 244046 101642 244102
rect 101698 244046 101766 244102
rect 101822 244046 101918 244102
rect 101298 243978 101918 244046
rect 101298 243922 101394 243978
rect 101450 243922 101518 243978
rect 101574 243922 101642 243978
rect 101698 243922 101766 243978
rect 101822 243922 101918 243978
rect 101298 226350 101918 243922
rect 101298 226294 101394 226350
rect 101450 226294 101518 226350
rect 101574 226294 101642 226350
rect 101698 226294 101766 226350
rect 101822 226294 101918 226350
rect 101298 226226 101918 226294
rect 101298 226170 101394 226226
rect 101450 226170 101518 226226
rect 101574 226170 101642 226226
rect 101698 226170 101766 226226
rect 101822 226170 101918 226226
rect 101298 226102 101918 226170
rect 101298 226046 101394 226102
rect 101450 226046 101518 226102
rect 101574 226046 101642 226102
rect 101698 226046 101766 226102
rect 101822 226046 101918 226102
rect 101298 225978 101918 226046
rect 101298 225922 101394 225978
rect 101450 225922 101518 225978
rect 101574 225922 101642 225978
rect 101698 225922 101766 225978
rect 101822 225922 101918 225978
rect 101298 208350 101918 225922
rect 101298 208294 101394 208350
rect 101450 208294 101518 208350
rect 101574 208294 101642 208350
rect 101698 208294 101766 208350
rect 101822 208294 101918 208350
rect 101298 208226 101918 208294
rect 101298 208170 101394 208226
rect 101450 208170 101518 208226
rect 101574 208170 101642 208226
rect 101698 208170 101766 208226
rect 101822 208170 101918 208226
rect 101298 208102 101918 208170
rect 101298 208046 101394 208102
rect 101450 208046 101518 208102
rect 101574 208046 101642 208102
rect 101698 208046 101766 208102
rect 101822 208046 101918 208102
rect 101298 207978 101918 208046
rect 101298 207922 101394 207978
rect 101450 207922 101518 207978
rect 101574 207922 101642 207978
rect 101698 207922 101766 207978
rect 101822 207922 101918 207978
rect 101298 190350 101918 207922
rect 101298 190294 101394 190350
rect 101450 190294 101518 190350
rect 101574 190294 101642 190350
rect 101698 190294 101766 190350
rect 101822 190294 101918 190350
rect 101298 190226 101918 190294
rect 101298 190170 101394 190226
rect 101450 190170 101518 190226
rect 101574 190170 101642 190226
rect 101698 190170 101766 190226
rect 101822 190170 101918 190226
rect 101298 190102 101918 190170
rect 101298 190046 101394 190102
rect 101450 190046 101518 190102
rect 101574 190046 101642 190102
rect 101698 190046 101766 190102
rect 101822 190046 101918 190102
rect 101298 189978 101918 190046
rect 101298 189922 101394 189978
rect 101450 189922 101518 189978
rect 101574 189922 101642 189978
rect 101698 189922 101766 189978
rect 101822 189922 101918 189978
rect 101298 172350 101918 189922
rect 101298 172294 101394 172350
rect 101450 172294 101518 172350
rect 101574 172294 101642 172350
rect 101698 172294 101766 172350
rect 101822 172294 101918 172350
rect 101298 172226 101918 172294
rect 101298 172170 101394 172226
rect 101450 172170 101518 172226
rect 101574 172170 101642 172226
rect 101698 172170 101766 172226
rect 101822 172170 101918 172226
rect 101298 172102 101918 172170
rect 101298 172046 101394 172102
rect 101450 172046 101518 172102
rect 101574 172046 101642 172102
rect 101698 172046 101766 172102
rect 101822 172046 101918 172102
rect 101298 171978 101918 172046
rect 101298 171922 101394 171978
rect 101450 171922 101518 171978
rect 101574 171922 101642 171978
rect 101698 171922 101766 171978
rect 101822 171922 101918 171978
rect 101298 154350 101918 171922
rect 101298 154294 101394 154350
rect 101450 154294 101518 154350
rect 101574 154294 101642 154350
rect 101698 154294 101766 154350
rect 101822 154294 101918 154350
rect 101298 154226 101918 154294
rect 101298 154170 101394 154226
rect 101450 154170 101518 154226
rect 101574 154170 101642 154226
rect 101698 154170 101766 154226
rect 101822 154170 101918 154226
rect 101298 154102 101918 154170
rect 101298 154046 101394 154102
rect 101450 154046 101518 154102
rect 101574 154046 101642 154102
rect 101698 154046 101766 154102
rect 101822 154046 101918 154102
rect 101298 153978 101918 154046
rect 101298 153922 101394 153978
rect 101450 153922 101518 153978
rect 101574 153922 101642 153978
rect 101698 153922 101766 153978
rect 101822 153922 101918 153978
rect 101298 136350 101918 153922
rect 101298 136294 101394 136350
rect 101450 136294 101518 136350
rect 101574 136294 101642 136350
rect 101698 136294 101766 136350
rect 101822 136294 101918 136350
rect 101298 136226 101918 136294
rect 101298 136170 101394 136226
rect 101450 136170 101518 136226
rect 101574 136170 101642 136226
rect 101698 136170 101766 136226
rect 101822 136170 101918 136226
rect 101298 136102 101918 136170
rect 101298 136046 101394 136102
rect 101450 136046 101518 136102
rect 101574 136046 101642 136102
rect 101698 136046 101766 136102
rect 101822 136046 101918 136102
rect 101298 135978 101918 136046
rect 101298 135922 101394 135978
rect 101450 135922 101518 135978
rect 101574 135922 101642 135978
rect 101698 135922 101766 135978
rect 101822 135922 101918 135978
rect 101298 118350 101918 135922
rect 101298 118294 101394 118350
rect 101450 118294 101518 118350
rect 101574 118294 101642 118350
rect 101698 118294 101766 118350
rect 101822 118294 101918 118350
rect 101298 118226 101918 118294
rect 101298 118170 101394 118226
rect 101450 118170 101518 118226
rect 101574 118170 101642 118226
rect 101698 118170 101766 118226
rect 101822 118170 101918 118226
rect 101298 118102 101918 118170
rect 101298 118046 101394 118102
rect 101450 118046 101518 118102
rect 101574 118046 101642 118102
rect 101698 118046 101766 118102
rect 101822 118046 101918 118102
rect 101298 117978 101918 118046
rect 101298 117922 101394 117978
rect 101450 117922 101518 117978
rect 101574 117922 101642 117978
rect 101698 117922 101766 117978
rect 101822 117922 101918 117978
rect 101298 100350 101918 117922
rect 101298 100294 101394 100350
rect 101450 100294 101518 100350
rect 101574 100294 101642 100350
rect 101698 100294 101766 100350
rect 101822 100294 101918 100350
rect 101298 100226 101918 100294
rect 101298 100170 101394 100226
rect 101450 100170 101518 100226
rect 101574 100170 101642 100226
rect 101698 100170 101766 100226
rect 101822 100170 101918 100226
rect 101298 100102 101918 100170
rect 101298 100046 101394 100102
rect 101450 100046 101518 100102
rect 101574 100046 101642 100102
rect 101698 100046 101766 100102
rect 101822 100046 101918 100102
rect 101298 99978 101918 100046
rect 101298 99922 101394 99978
rect 101450 99922 101518 99978
rect 101574 99922 101642 99978
rect 101698 99922 101766 99978
rect 101822 99922 101918 99978
rect 101298 82350 101918 99922
rect 120988 590212 121044 590222
rect 101298 82294 101394 82350
rect 101450 82294 101518 82350
rect 101574 82294 101642 82350
rect 101698 82294 101766 82350
rect 101822 82294 101918 82350
rect 101298 82226 101918 82294
rect 101298 82170 101394 82226
rect 101450 82170 101518 82226
rect 101574 82170 101642 82226
rect 101698 82170 101766 82226
rect 101822 82170 101918 82226
rect 101298 82102 101918 82170
rect 101298 82046 101394 82102
rect 101450 82046 101518 82102
rect 101574 82046 101642 82102
rect 101698 82046 101766 82102
rect 101822 82046 101918 82102
rect 101298 81978 101918 82046
rect 101298 81922 101394 81978
rect 101450 81922 101518 81978
rect 101574 81922 101642 81978
rect 101698 81922 101766 81978
rect 101822 81922 101918 81978
rect 97578 76294 97674 76350
rect 97730 76294 97798 76350
rect 97854 76294 97922 76350
rect 97978 76294 98046 76350
rect 98102 76294 98198 76350
rect 97578 76226 98198 76294
rect 97578 76170 97674 76226
rect 97730 76170 97798 76226
rect 97854 76170 97922 76226
rect 97978 76170 98046 76226
rect 98102 76170 98198 76226
rect 97578 76102 98198 76170
rect 97578 76046 97674 76102
rect 97730 76046 97798 76102
rect 97854 76046 97922 76102
rect 97978 76046 98046 76102
rect 98102 76046 98198 76102
rect 97578 75978 98198 76046
rect 97578 75922 97674 75978
rect 97730 75922 97798 75978
rect 97854 75922 97922 75978
rect 97978 75922 98046 75978
rect 98102 75922 98198 75978
rect 94444 75684 94500 75694
rect 93248 64350 93568 64384
rect 93248 64294 93318 64350
rect 93374 64294 93442 64350
rect 93498 64294 93568 64350
rect 93248 64226 93568 64294
rect 93248 64170 93318 64226
rect 93374 64170 93442 64226
rect 93498 64170 93568 64226
rect 93248 64102 93568 64170
rect 93248 64046 93318 64102
rect 93374 64046 93442 64102
rect 93498 64046 93568 64102
rect 93248 63978 93568 64046
rect 93248 63922 93318 63978
rect 93374 63922 93442 63978
rect 93498 63922 93568 63978
rect 93248 63888 93568 63922
rect 92876 60598 92932 60608
rect 92764 57358 92820 57368
rect 92428 8758 92484 8768
rect 92428 5518 92484 8702
rect 92428 5452 92484 5462
rect 92764 4340 92820 57302
rect 92764 4274 92820 4284
rect 92316 3378 92372 3388
rect 92204 3266 92260 3276
rect 92876 3332 92932 60542
rect 94220 52318 94276 52328
rect 93248 46350 93568 46384
rect 93248 46294 93318 46350
rect 93374 46294 93442 46350
rect 93498 46294 93568 46350
rect 93248 46226 93568 46294
rect 93248 46170 93318 46226
rect 93374 46170 93442 46226
rect 93498 46170 93568 46226
rect 93248 46102 93568 46170
rect 93248 46046 93318 46102
rect 93374 46046 93442 46102
rect 93498 46046 93568 46102
rect 93248 45978 93568 46046
rect 93248 45922 93318 45978
rect 93374 45922 93442 45978
rect 93498 45922 93568 45978
rect 93248 45888 93568 45922
rect 93248 28350 93568 28384
rect 93248 28294 93318 28350
rect 93374 28294 93442 28350
rect 93498 28294 93568 28350
rect 93248 28226 93568 28294
rect 93248 28170 93318 28226
rect 93374 28170 93442 28226
rect 93498 28170 93568 28226
rect 93248 28102 93568 28170
rect 93248 28046 93318 28102
rect 93374 28046 93442 28102
rect 93498 28046 93568 28102
rect 93248 27978 93568 28046
rect 93248 27922 93318 27978
rect 93374 27922 93442 27978
rect 93498 27922 93568 27978
rect 93248 27888 93568 27922
rect 93884 25498 93940 25508
rect 93772 16858 93828 16868
rect 93660 15238 93716 15248
rect 93100 10738 93156 10748
rect 92988 10682 93100 10738
rect 92988 3892 93044 10682
rect 93100 10672 93156 10682
rect 93248 10350 93568 10384
rect 93248 10294 93318 10350
rect 93374 10294 93442 10350
rect 93498 10294 93568 10350
rect 93248 10226 93568 10294
rect 93248 10170 93318 10226
rect 93374 10170 93442 10226
rect 93498 10170 93568 10226
rect 93248 10102 93568 10170
rect 93248 10046 93318 10102
rect 93374 10046 93442 10102
rect 93498 10046 93568 10102
rect 93248 9978 93568 10046
rect 93248 9922 93318 9978
rect 93374 9922 93442 9978
rect 93498 9922 93568 9978
rect 93248 9888 93568 9922
rect 93212 5338 93268 5348
rect 92988 3826 93044 3836
rect 93100 4618 93156 4628
rect 93100 3444 93156 4562
rect 93100 3378 93156 3388
rect 92876 3266 92932 3276
rect 91532 2594 91588 2604
rect 93212 2660 93268 5282
rect 93324 4564 93380 4574
rect 93324 3892 93380 4508
rect 93324 3826 93380 3836
rect 93436 4340 93492 4350
rect 93436 3444 93492 4284
rect 93660 3780 93716 15182
rect 93660 3714 93716 3724
rect 93436 3378 93492 3388
rect 93772 3220 93828 16802
rect 93884 11818 93940 25442
rect 93884 11752 93940 11762
rect 93772 3154 93828 3164
rect 93884 5158 93940 5168
rect 93212 2594 93268 2604
rect 93884 1204 93940 5102
rect 94220 3780 94276 52262
rect 94220 3714 94276 3724
rect 94444 3220 94500 75628
rect 94892 71398 94948 71408
rect 94892 54658 94948 71342
rect 95676 62218 95732 62228
rect 95564 58978 95620 58988
rect 94892 54592 94948 54602
rect 95452 55738 95508 55748
rect 94892 54118 94948 54128
rect 94892 15238 94948 54062
rect 95340 44218 95396 44228
rect 95340 41338 95396 44162
rect 95340 41272 95396 41282
rect 94892 15172 94948 15182
rect 95340 15058 95396 15068
rect 95004 15002 95340 15058
rect 94444 3154 94500 3164
rect 94892 7498 94948 7508
rect 93996 1876 94052 1886
rect 93996 1428 94052 1820
rect 93996 1362 94052 1372
rect 93884 1138 93940 1148
rect 90972 1026 91028 1036
rect 85708 952 85764 962
rect 94892 532 94948 7442
rect 95004 1540 95060 15002
rect 95340 14992 95396 15002
rect 95340 6958 95396 6968
rect 95228 2996 95284 3006
rect 95228 2660 95284 2940
rect 95228 2594 95284 2604
rect 95340 1652 95396 6902
rect 95452 3780 95508 55682
rect 95452 3714 95508 3724
rect 95564 3332 95620 58922
rect 95676 3444 95732 62162
rect 97578 58350 98198 75922
rect 100156 77364 100212 77374
rect 97578 58294 97674 58350
rect 97730 58294 97798 58350
rect 97854 58294 97922 58350
rect 97978 58294 98046 58350
rect 98102 58294 98198 58350
rect 97578 58226 98198 58294
rect 97578 58170 97674 58226
rect 97730 58170 97798 58226
rect 97854 58170 97922 58226
rect 97978 58170 98046 58226
rect 98102 58170 98198 58226
rect 97578 58102 98198 58170
rect 97578 58046 97674 58102
rect 97730 58046 97798 58102
rect 97854 58046 97922 58102
rect 97978 58046 98046 58102
rect 98102 58046 98198 58102
rect 97578 57978 98198 58046
rect 97578 57922 97674 57978
rect 97730 57922 97798 57978
rect 97854 57922 97922 57978
rect 97978 57922 98046 57978
rect 98102 57922 98198 57978
rect 96460 57178 96516 57188
rect 96236 50698 96292 50708
rect 96012 47098 96068 47108
rect 95676 3378 95732 3388
rect 95900 15238 95956 15248
rect 95564 3266 95620 3276
rect 95900 2772 95956 15182
rect 96012 3780 96068 47042
rect 96012 3714 96068 3724
rect 96236 3780 96292 50642
rect 96236 3714 96292 3724
rect 96348 5518 96404 5528
rect 95900 2706 95956 2716
rect 96348 2548 96404 5462
rect 96460 3780 96516 57122
rect 96572 54658 96628 54668
rect 96572 53038 96628 54602
rect 96572 52972 96628 52982
rect 97356 50518 97412 50528
rect 97244 40618 97300 40628
rect 96460 3714 96516 3724
rect 97132 15238 97188 15248
rect 97132 3332 97188 15182
rect 97244 3780 97300 40562
rect 97244 3714 97300 3724
rect 97356 3444 97412 50462
rect 97356 3378 97412 3388
rect 97578 40350 98198 57922
rect 99932 74278 99988 74288
rect 99372 55558 99428 55568
rect 97578 40294 97674 40350
rect 97730 40294 97798 40350
rect 97854 40294 97922 40350
rect 97978 40294 98046 40350
rect 98102 40294 98198 40350
rect 97578 40226 98198 40294
rect 97578 40170 97674 40226
rect 97730 40170 97798 40226
rect 97854 40170 97922 40226
rect 97978 40170 98046 40226
rect 98102 40170 98198 40226
rect 97578 40102 98198 40170
rect 97578 40046 97674 40102
rect 97730 40046 97798 40102
rect 97854 40046 97922 40102
rect 97978 40046 98046 40102
rect 98102 40046 98198 40102
rect 97578 39978 98198 40046
rect 97578 39922 97674 39978
rect 97730 39922 97798 39978
rect 97854 39922 97922 39978
rect 97978 39922 98046 39978
rect 98102 39922 98198 39978
rect 97578 22350 98198 39922
rect 97578 22294 97674 22350
rect 97730 22294 97798 22350
rect 97854 22294 97922 22350
rect 97978 22294 98046 22350
rect 98102 22294 98198 22350
rect 97578 22226 98198 22294
rect 97578 22170 97674 22226
rect 97730 22170 97798 22226
rect 97854 22170 97922 22226
rect 97978 22170 98046 22226
rect 98102 22170 98198 22226
rect 97578 22102 98198 22170
rect 97578 22046 97674 22102
rect 97730 22046 97798 22102
rect 97854 22046 97922 22102
rect 97978 22046 98046 22102
rect 98102 22046 98198 22102
rect 97578 21978 98198 22046
rect 97578 21922 97674 21978
rect 97730 21922 97798 21978
rect 97854 21922 97922 21978
rect 97978 21922 98046 21978
rect 98102 21922 98198 21978
rect 97578 4350 98198 21922
rect 97578 4294 97674 4350
rect 97730 4294 97798 4350
rect 97854 4294 97922 4350
rect 97978 4294 98046 4350
rect 98102 4294 98198 4350
rect 97578 4226 98198 4294
rect 97578 4170 97674 4226
rect 97730 4170 97798 4226
rect 97854 4170 97922 4226
rect 97978 4170 98046 4226
rect 98102 4170 98198 4226
rect 97578 4102 98198 4170
rect 97578 4046 97674 4102
rect 97730 4046 97798 4102
rect 97854 4046 97922 4102
rect 97978 4046 98046 4102
rect 98102 4046 98198 4102
rect 97578 3978 98198 4046
rect 97578 3922 97674 3978
rect 97730 3922 97798 3978
rect 97854 3922 97922 3978
rect 97978 3922 98046 3978
rect 98102 3922 98198 3978
rect 97132 3266 97188 3276
rect 96348 2482 96404 2492
rect 95340 1586 95396 1596
rect 95004 1474 95060 1484
rect 94892 466 94948 476
rect 84924 242 84980 252
rect 70578 -1176 70674 -1120
rect 70730 -1176 70798 -1120
rect 70854 -1176 70922 -1120
rect 70978 -1176 71046 -1120
rect 71102 -1176 71198 -1120
rect 70578 -1244 71198 -1176
rect 70578 -1300 70674 -1244
rect 70730 -1300 70798 -1244
rect 70854 -1300 70922 -1244
rect 70978 -1300 71046 -1244
rect 71102 -1300 71198 -1244
rect 70578 -1368 71198 -1300
rect 70578 -1424 70674 -1368
rect 70730 -1424 70798 -1368
rect 70854 -1424 70922 -1368
rect 70978 -1424 71046 -1368
rect 71102 -1424 71198 -1368
rect 70578 -1492 71198 -1424
rect 70578 -1548 70674 -1492
rect 70730 -1548 70798 -1492
rect 70854 -1548 70922 -1492
rect 70978 -1548 71046 -1492
rect 71102 -1548 71198 -1492
rect 70578 -1644 71198 -1548
rect 97578 -160 98198 3922
rect 98588 52138 98644 52148
rect 98588 3780 98644 52082
rect 98588 3714 98644 3724
rect 98700 48898 98756 48908
rect 98700 3444 98756 48842
rect 98700 3378 98756 3388
rect 98812 19378 98868 19388
rect 98812 3332 98868 19322
rect 98812 3266 98868 3276
rect 99036 7858 99092 7868
rect 98924 3220 98980 3230
rect 98924 3112 98980 3122
rect 99036 2772 99092 7802
rect 99372 3780 99428 55502
rect 99820 31978 99876 31988
rect 99372 3714 99428 3724
rect 99596 6778 99652 6788
rect 99596 3780 99652 6722
rect 99596 3714 99652 3724
rect 99820 3780 99876 31922
rect 99932 19378 99988 74222
rect 99932 19312 99988 19322
rect 100044 42058 100100 42068
rect 100044 6058 100100 42002
rect 100044 5992 100100 6002
rect 99820 3714 99876 3724
rect 100156 3780 100212 77308
rect 100604 67258 100660 67268
rect 100156 3714 100212 3724
rect 100492 53938 100548 53948
rect 100492 3444 100548 53882
rect 100604 3780 100660 67202
rect 100604 3714 100660 3724
rect 101298 64350 101918 81922
rect 114268 82740 114324 82750
rect 110908 81060 110964 81070
rect 101298 64294 101394 64350
rect 101450 64294 101518 64350
rect 101574 64294 101642 64350
rect 101698 64294 101766 64350
rect 101822 64294 101918 64350
rect 101298 64226 101918 64294
rect 101298 64170 101394 64226
rect 101450 64170 101518 64226
rect 101574 64170 101642 64226
rect 101698 64170 101766 64226
rect 101822 64170 101918 64226
rect 101298 64102 101918 64170
rect 101298 64046 101394 64102
rect 101450 64046 101518 64102
rect 101574 64046 101642 64102
rect 101698 64046 101766 64102
rect 101822 64046 101918 64102
rect 101298 63978 101918 64046
rect 101298 63922 101394 63978
rect 101450 63922 101518 63978
rect 101574 63922 101642 63978
rect 101698 63922 101766 63978
rect 101822 63922 101918 63978
rect 101298 46350 101918 63922
rect 101298 46294 101394 46350
rect 101450 46294 101518 46350
rect 101574 46294 101642 46350
rect 101698 46294 101766 46350
rect 101822 46294 101918 46350
rect 101298 46226 101918 46294
rect 101298 46170 101394 46226
rect 101450 46170 101518 46226
rect 101574 46170 101642 46226
rect 101698 46170 101766 46226
rect 101822 46170 101918 46226
rect 101298 46102 101918 46170
rect 101298 46046 101394 46102
rect 101450 46046 101518 46102
rect 101574 46046 101642 46102
rect 101698 46046 101766 46102
rect 101822 46046 101918 46102
rect 101298 45978 101918 46046
rect 101298 45922 101394 45978
rect 101450 45922 101518 45978
rect 101574 45922 101642 45978
rect 101698 45922 101766 45978
rect 101822 45922 101918 45978
rect 101298 28350 101918 45922
rect 101298 28294 101394 28350
rect 101450 28294 101518 28350
rect 101574 28294 101642 28350
rect 101698 28294 101766 28350
rect 101822 28294 101918 28350
rect 101298 28226 101918 28294
rect 101298 28170 101394 28226
rect 101450 28170 101518 28226
rect 101574 28170 101642 28226
rect 101698 28170 101766 28226
rect 101822 28170 101918 28226
rect 101298 28102 101918 28170
rect 101298 28046 101394 28102
rect 101450 28046 101518 28102
rect 101574 28046 101642 28102
rect 101698 28046 101766 28102
rect 101822 28046 101918 28102
rect 101298 27978 101918 28046
rect 101298 27922 101394 27978
rect 101450 27922 101518 27978
rect 101574 27922 101642 27978
rect 101698 27922 101766 27978
rect 101822 27922 101918 27978
rect 101298 10350 101918 27922
rect 101298 10294 101394 10350
rect 101450 10294 101518 10350
rect 101574 10294 101642 10350
rect 101698 10294 101766 10350
rect 101822 10294 101918 10350
rect 101298 10226 101918 10294
rect 101298 10170 101394 10226
rect 101450 10170 101518 10226
rect 101574 10170 101642 10226
rect 101698 10170 101766 10226
rect 101822 10170 101918 10226
rect 101298 10102 101918 10170
rect 101298 10046 101394 10102
rect 101450 10046 101518 10102
rect 101574 10046 101642 10102
rect 101698 10046 101766 10102
rect 101822 10046 101918 10102
rect 101298 9978 101918 10046
rect 101298 9922 101394 9978
rect 101450 9922 101518 9978
rect 101574 9922 101642 9978
rect 101698 9922 101766 9978
rect 101822 9922 101918 9978
rect 100492 3378 100548 3388
rect 99036 2706 99092 2716
rect 98476 1652 98532 1662
rect 98476 1198 98532 1596
rect 99148 1652 99204 1662
rect 99148 1378 99204 1596
rect 100492 1652 100548 1662
rect 100492 1558 100548 1596
rect 100492 1492 100548 1502
rect 99148 1312 99204 1322
rect 98476 1132 98532 1142
rect 97578 -216 97674 -160
rect 97730 -216 97798 -160
rect 97854 -216 97922 -160
rect 97978 -216 98046 -160
rect 98102 -216 98198 -160
rect 97578 -284 98198 -216
rect 97578 -340 97674 -284
rect 97730 -340 97798 -284
rect 97854 -340 97922 -284
rect 97978 -340 98046 -284
rect 98102 -340 98198 -284
rect 97578 -408 98198 -340
rect 97578 -464 97674 -408
rect 97730 -464 97798 -408
rect 97854 -464 97922 -408
rect 97978 -464 98046 -408
rect 98102 -464 98198 -408
rect 97578 -532 98198 -464
rect 97578 -588 97674 -532
rect 97730 -588 97798 -532
rect 97854 -588 97922 -532
rect 97978 -588 98046 -532
rect 98102 -588 98198 -532
rect 97578 -1644 98198 -588
rect 101298 -1120 101918 9922
rect 102060 65638 102116 65648
rect 102060 3444 102116 65582
rect 108608 58350 108928 58384
rect 108608 58294 108678 58350
rect 108734 58294 108802 58350
rect 108858 58294 108928 58350
rect 108608 58226 108928 58294
rect 108608 58170 108678 58226
rect 108734 58170 108802 58226
rect 108858 58170 108928 58226
rect 108608 58102 108928 58170
rect 108608 58046 108678 58102
rect 108734 58046 108802 58102
rect 108858 58046 108928 58102
rect 108608 57978 108928 58046
rect 108608 57922 108678 57978
rect 108734 57922 108802 57978
rect 108858 57922 108928 57978
rect 108608 57888 108928 57922
rect 110796 56458 110852 56468
rect 110796 49618 110852 56402
rect 110796 49552 110852 49562
rect 108608 40350 108928 40384
rect 108608 40294 108678 40350
rect 108734 40294 108802 40350
rect 108858 40294 108928 40350
rect 108608 40226 108928 40294
rect 108608 40170 108678 40226
rect 108734 40170 108802 40226
rect 108858 40170 108928 40226
rect 108608 40102 108928 40170
rect 108608 40046 108678 40102
rect 108734 40046 108802 40102
rect 108858 40046 108928 40102
rect 108608 39978 108928 40046
rect 108608 39922 108678 39978
rect 108734 39922 108802 39978
rect 108858 39922 108928 39978
rect 108608 39888 108928 39922
rect 103292 35398 103348 35408
rect 102396 20998 102452 21008
rect 102396 3780 102452 20942
rect 103292 4618 103348 35342
rect 109228 31258 109284 31268
rect 104076 30718 104132 30728
rect 104076 26038 104132 30662
rect 104076 25972 104132 25982
rect 107548 25318 107604 25328
rect 104188 11998 104244 12008
rect 103404 11818 103460 11828
rect 103404 6958 103460 11762
rect 103404 6892 103460 6902
rect 103292 4552 103348 4562
rect 102396 3714 102452 3724
rect 104188 3556 104244 11942
rect 104188 3490 104244 3500
rect 106540 3556 106596 3566
rect 102060 3378 102116 3388
rect 106540 3358 106596 3500
rect 107548 3556 107604 25262
rect 108332 25318 108388 25328
rect 108332 20998 108388 25262
rect 108608 22350 108928 22384
rect 108608 22294 108678 22350
rect 108734 22294 108802 22350
rect 108858 22294 108928 22350
rect 108608 22226 108928 22294
rect 108608 22170 108678 22226
rect 108734 22170 108802 22226
rect 108858 22170 108928 22226
rect 108608 22102 108928 22170
rect 108608 22046 108678 22102
rect 108734 22046 108802 22102
rect 108858 22046 108928 22102
rect 108608 21978 108928 22046
rect 108608 21922 108678 21978
rect 108734 21922 108802 21978
rect 108858 21922 108928 21978
rect 108608 21888 108928 21922
rect 108332 20932 108388 20942
rect 108332 7498 108388 7508
rect 108332 6958 108388 7442
rect 108332 6892 108388 6902
rect 107548 3490 107604 3500
rect 109228 3556 109284 31202
rect 109228 3490 109284 3500
rect 110908 3556 110964 81004
rect 111020 11998 111076 12008
rect 111020 11098 111076 11942
rect 111020 11032 111076 11042
rect 110908 3490 110964 3500
rect 114268 3444 114324 82684
rect 119308 80948 119364 80958
rect 115948 34678 116004 34688
rect 115836 33958 115892 33968
rect 115836 32698 115892 33902
rect 115836 32632 115892 32642
rect 115948 20188 116004 34622
rect 115948 20132 116116 20188
rect 116060 3556 116116 20132
rect 116060 3490 116116 3500
rect 119308 3556 119364 80892
rect 120988 78418 121044 590156
rect 128298 580350 128918 596784
rect 128298 580294 128394 580350
rect 128450 580294 128518 580350
rect 128574 580294 128642 580350
rect 128698 580294 128766 580350
rect 128822 580294 128918 580350
rect 128298 580226 128918 580294
rect 128298 580170 128394 580226
rect 128450 580170 128518 580226
rect 128574 580170 128642 580226
rect 128698 580170 128766 580226
rect 128822 580170 128918 580226
rect 128298 580102 128918 580170
rect 128298 580046 128394 580102
rect 128450 580046 128518 580102
rect 128574 580046 128642 580102
rect 128698 580046 128766 580102
rect 128822 580046 128918 580102
rect 128298 579978 128918 580046
rect 128298 579922 128394 579978
rect 128450 579922 128518 579978
rect 128574 579922 128642 579978
rect 128698 579922 128766 579978
rect 128822 579922 128918 579978
rect 128298 562350 128918 579922
rect 128298 562294 128394 562350
rect 128450 562294 128518 562350
rect 128574 562294 128642 562350
rect 128698 562294 128766 562350
rect 128822 562294 128918 562350
rect 128298 562226 128918 562294
rect 128298 562170 128394 562226
rect 128450 562170 128518 562226
rect 128574 562170 128642 562226
rect 128698 562170 128766 562226
rect 128822 562170 128918 562226
rect 128298 562102 128918 562170
rect 128298 562046 128394 562102
rect 128450 562046 128518 562102
rect 128574 562046 128642 562102
rect 128698 562046 128766 562102
rect 128822 562046 128918 562102
rect 128298 561978 128918 562046
rect 128298 561922 128394 561978
rect 128450 561922 128518 561978
rect 128574 561922 128642 561978
rect 128698 561922 128766 561978
rect 128822 561922 128918 561978
rect 128298 544350 128918 561922
rect 128298 544294 128394 544350
rect 128450 544294 128518 544350
rect 128574 544294 128642 544350
rect 128698 544294 128766 544350
rect 128822 544294 128918 544350
rect 128298 544226 128918 544294
rect 128298 544170 128394 544226
rect 128450 544170 128518 544226
rect 128574 544170 128642 544226
rect 128698 544170 128766 544226
rect 128822 544170 128918 544226
rect 128298 544102 128918 544170
rect 128298 544046 128394 544102
rect 128450 544046 128518 544102
rect 128574 544046 128642 544102
rect 128698 544046 128766 544102
rect 128822 544046 128918 544102
rect 128298 543978 128918 544046
rect 128298 543922 128394 543978
rect 128450 543922 128518 543978
rect 128574 543922 128642 543978
rect 128698 543922 128766 543978
rect 128822 543922 128918 543978
rect 128298 526350 128918 543922
rect 128298 526294 128394 526350
rect 128450 526294 128518 526350
rect 128574 526294 128642 526350
rect 128698 526294 128766 526350
rect 128822 526294 128918 526350
rect 128298 526226 128918 526294
rect 128298 526170 128394 526226
rect 128450 526170 128518 526226
rect 128574 526170 128642 526226
rect 128698 526170 128766 526226
rect 128822 526170 128918 526226
rect 128298 526102 128918 526170
rect 128298 526046 128394 526102
rect 128450 526046 128518 526102
rect 128574 526046 128642 526102
rect 128698 526046 128766 526102
rect 128822 526046 128918 526102
rect 128298 525978 128918 526046
rect 128298 525922 128394 525978
rect 128450 525922 128518 525978
rect 128574 525922 128642 525978
rect 128698 525922 128766 525978
rect 128822 525922 128918 525978
rect 128298 508350 128918 525922
rect 128298 508294 128394 508350
rect 128450 508294 128518 508350
rect 128574 508294 128642 508350
rect 128698 508294 128766 508350
rect 128822 508294 128918 508350
rect 128298 508226 128918 508294
rect 128298 508170 128394 508226
rect 128450 508170 128518 508226
rect 128574 508170 128642 508226
rect 128698 508170 128766 508226
rect 128822 508170 128918 508226
rect 128298 508102 128918 508170
rect 128298 508046 128394 508102
rect 128450 508046 128518 508102
rect 128574 508046 128642 508102
rect 128698 508046 128766 508102
rect 128822 508046 128918 508102
rect 128298 507978 128918 508046
rect 128298 507922 128394 507978
rect 128450 507922 128518 507978
rect 128574 507922 128642 507978
rect 128698 507922 128766 507978
rect 128822 507922 128918 507978
rect 128298 490350 128918 507922
rect 128298 490294 128394 490350
rect 128450 490294 128518 490350
rect 128574 490294 128642 490350
rect 128698 490294 128766 490350
rect 128822 490294 128918 490350
rect 128298 490226 128918 490294
rect 128298 490170 128394 490226
rect 128450 490170 128518 490226
rect 128574 490170 128642 490226
rect 128698 490170 128766 490226
rect 128822 490170 128918 490226
rect 128298 490102 128918 490170
rect 128298 490046 128394 490102
rect 128450 490046 128518 490102
rect 128574 490046 128642 490102
rect 128698 490046 128766 490102
rect 128822 490046 128918 490102
rect 128298 489978 128918 490046
rect 128298 489922 128394 489978
rect 128450 489922 128518 489978
rect 128574 489922 128642 489978
rect 128698 489922 128766 489978
rect 128822 489922 128918 489978
rect 128298 472350 128918 489922
rect 128298 472294 128394 472350
rect 128450 472294 128518 472350
rect 128574 472294 128642 472350
rect 128698 472294 128766 472350
rect 128822 472294 128918 472350
rect 128298 472226 128918 472294
rect 128298 472170 128394 472226
rect 128450 472170 128518 472226
rect 128574 472170 128642 472226
rect 128698 472170 128766 472226
rect 128822 472170 128918 472226
rect 128298 472102 128918 472170
rect 128298 472046 128394 472102
rect 128450 472046 128518 472102
rect 128574 472046 128642 472102
rect 128698 472046 128766 472102
rect 128822 472046 128918 472102
rect 128298 471978 128918 472046
rect 128298 471922 128394 471978
rect 128450 471922 128518 471978
rect 128574 471922 128642 471978
rect 128698 471922 128766 471978
rect 128822 471922 128918 471978
rect 128298 454350 128918 471922
rect 128298 454294 128394 454350
rect 128450 454294 128518 454350
rect 128574 454294 128642 454350
rect 128698 454294 128766 454350
rect 128822 454294 128918 454350
rect 128298 454226 128918 454294
rect 128298 454170 128394 454226
rect 128450 454170 128518 454226
rect 128574 454170 128642 454226
rect 128698 454170 128766 454226
rect 128822 454170 128918 454226
rect 128298 454102 128918 454170
rect 128298 454046 128394 454102
rect 128450 454046 128518 454102
rect 128574 454046 128642 454102
rect 128698 454046 128766 454102
rect 128822 454046 128918 454102
rect 128298 453978 128918 454046
rect 128298 453922 128394 453978
rect 128450 453922 128518 453978
rect 128574 453922 128642 453978
rect 128698 453922 128766 453978
rect 128822 453922 128918 453978
rect 128298 436350 128918 453922
rect 128298 436294 128394 436350
rect 128450 436294 128518 436350
rect 128574 436294 128642 436350
rect 128698 436294 128766 436350
rect 128822 436294 128918 436350
rect 128298 436226 128918 436294
rect 128298 436170 128394 436226
rect 128450 436170 128518 436226
rect 128574 436170 128642 436226
rect 128698 436170 128766 436226
rect 128822 436170 128918 436226
rect 128298 436102 128918 436170
rect 128298 436046 128394 436102
rect 128450 436046 128518 436102
rect 128574 436046 128642 436102
rect 128698 436046 128766 436102
rect 128822 436046 128918 436102
rect 128298 435978 128918 436046
rect 128298 435922 128394 435978
rect 128450 435922 128518 435978
rect 128574 435922 128642 435978
rect 128698 435922 128766 435978
rect 128822 435922 128918 435978
rect 128298 418350 128918 435922
rect 128298 418294 128394 418350
rect 128450 418294 128518 418350
rect 128574 418294 128642 418350
rect 128698 418294 128766 418350
rect 128822 418294 128918 418350
rect 128298 418226 128918 418294
rect 128298 418170 128394 418226
rect 128450 418170 128518 418226
rect 128574 418170 128642 418226
rect 128698 418170 128766 418226
rect 128822 418170 128918 418226
rect 128298 418102 128918 418170
rect 128298 418046 128394 418102
rect 128450 418046 128518 418102
rect 128574 418046 128642 418102
rect 128698 418046 128766 418102
rect 128822 418046 128918 418102
rect 128298 417978 128918 418046
rect 128298 417922 128394 417978
rect 128450 417922 128518 417978
rect 128574 417922 128642 417978
rect 128698 417922 128766 417978
rect 128822 417922 128918 417978
rect 128298 400350 128918 417922
rect 128298 400294 128394 400350
rect 128450 400294 128518 400350
rect 128574 400294 128642 400350
rect 128698 400294 128766 400350
rect 128822 400294 128918 400350
rect 128298 400226 128918 400294
rect 128298 400170 128394 400226
rect 128450 400170 128518 400226
rect 128574 400170 128642 400226
rect 128698 400170 128766 400226
rect 128822 400170 128918 400226
rect 128298 400102 128918 400170
rect 128298 400046 128394 400102
rect 128450 400046 128518 400102
rect 128574 400046 128642 400102
rect 128698 400046 128766 400102
rect 128822 400046 128918 400102
rect 128298 399978 128918 400046
rect 128298 399922 128394 399978
rect 128450 399922 128518 399978
rect 128574 399922 128642 399978
rect 128698 399922 128766 399978
rect 128822 399922 128918 399978
rect 128298 382350 128918 399922
rect 128298 382294 128394 382350
rect 128450 382294 128518 382350
rect 128574 382294 128642 382350
rect 128698 382294 128766 382350
rect 128822 382294 128918 382350
rect 128298 382226 128918 382294
rect 128298 382170 128394 382226
rect 128450 382170 128518 382226
rect 128574 382170 128642 382226
rect 128698 382170 128766 382226
rect 128822 382170 128918 382226
rect 128298 382102 128918 382170
rect 128298 382046 128394 382102
rect 128450 382046 128518 382102
rect 128574 382046 128642 382102
rect 128698 382046 128766 382102
rect 128822 382046 128918 382102
rect 128298 381978 128918 382046
rect 128298 381922 128394 381978
rect 128450 381922 128518 381978
rect 128574 381922 128642 381978
rect 128698 381922 128766 381978
rect 128822 381922 128918 381978
rect 128298 364350 128918 381922
rect 128298 364294 128394 364350
rect 128450 364294 128518 364350
rect 128574 364294 128642 364350
rect 128698 364294 128766 364350
rect 128822 364294 128918 364350
rect 128298 364226 128918 364294
rect 128298 364170 128394 364226
rect 128450 364170 128518 364226
rect 128574 364170 128642 364226
rect 128698 364170 128766 364226
rect 128822 364170 128918 364226
rect 128298 364102 128918 364170
rect 128298 364046 128394 364102
rect 128450 364046 128518 364102
rect 128574 364046 128642 364102
rect 128698 364046 128766 364102
rect 128822 364046 128918 364102
rect 128298 363978 128918 364046
rect 128298 363922 128394 363978
rect 128450 363922 128518 363978
rect 128574 363922 128642 363978
rect 128698 363922 128766 363978
rect 128822 363922 128918 363978
rect 128298 346350 128918 363922
rect 128298 346294 128394 346350
rect 128450 346294 128518 346350
rect 128574 346294 128642 346350
rect 128698 346294 128766 346350
rect 128822 346294 128918 346350
rect 128298 346226 128918 346294
rect 128298 346170 128394 346226
rect 128450 346170 128518 346226
rect 128574 346170 128642 346226
rect 128698 346170 128766 346226
rect 128822 346170 128918 346226
rect 128298 346102 128918 346170
rect 128298 346046 128394 346102
rect 128450 346046 128518 346102
rect 128574 346046 128642 346102
rect 128698 346046 128766 346102
rect 128822 346046 128918 346102
rect 128298 345978 128918 346046
rect 128298 345922 128394 345978
rect 128450 345922 128518 345978
rect 128574 345922 128642 345978
rect 128698 345922 128766 345978
rect 128822 345922 128918 345978
rect 128298 328350 128918 345922
rect 128298 328294 128394 328350
rect 128450 328294 128518 328350
rect 128574 328294 128642 328350
rect 128698 328294 128766 328350
rect 128822 328294 128918 328350
rect 128298 328226 128918 328294
rect 128298 328170 128394 328226
rect 128450 328170 128518 328226
rect 128574 328170 128642 328226
rect 128698 328170 128766 328226
rect 128822 328170 128918 328226
rect 128298 328102 128918 328170
rect 128298 328046 128394 328102
rect 128450 328046 128518 328102
rect 128574 328046 128642 328102
rect 128698 328046 128766 328102
rect 128822 328046 128918 328102
rect 128298 327978 128918 328046
rect 128298 327922 128394 327978
rect 128450 327922 128518 327978
rect 128574 327922 128642 327978
rect 128698 327922 128766 327978
rect 128822 327922 128918 327978
rect 126812 311108 126868 311118
rect 120988 78352 121044 78362
rect 121100 82628 121156 82638
rect 120092 54658 120148 54668
rect 120092 42778 120148 54602
rect 120092 42712 120148 42722
rect 120988 5338 121044 5348
rect 120988 4228 121044 5282
rect 120988 4162 121044 4172
rect 119308 3490 119364 3500
rect 121100 3556 121156 82572
rect 123788 74278 123844 74288
rect 121100 3490 121156 3500
rect 121772 74004 121828 74014
rect 114268 3378 114324 3388
rect 106540 3292 106596 3302
rect 121772 2548 121828 73948
rect 123788 20188 123844 74222
rect 126812 72548 126868 311052
rect 128298 310350 128918 327922
rect 128298 310294 128394 310350
rect 128450 310294 128518 310350
rect 128574 310294 128642 310350
rect 128698 310294 128766 310350
rect 128822 310294 128918 310350
rect 128298 310226 128918 310294
rect 128298 310170 128394 310226
rect 128450 310170 128518 310226
rect 128574 310170 128642 310226
rect 128698 310170 128766 310226
rect 128822 310170 128918 310226
rect 128298 310102 128918 310170
rect 128298 310046 128394 310102
rect 128450 310046 128518 310102
rect 128574 310046 128642 310102
rect 128698 310046 128766 310102
rect 128822 310046 128918 310102
rect 128298 309978 128918 310046
rect 128298 309922 128394 309978
rect 128450 309922 128518 309978
rect 128574 309922 128642 309978
rect 128698 309922 128766 309978
rect 128822 309922 128918 309978
rect 128298 292350 128918 309922
rect 128298 292294 128394 292350
rect 128450 292294 128518 292350
rect 128574 292294 128642 292350
rect 128698 292294 128766 292350
rect 128822 292294 128918 292350
rect 128298 292226 128918 292294
rect 128298 292170 128394 292226
rect 128450 292170 128518 292226
rect 128574 292170 128642 292226
rect 128698 292170 128766 292226
rect 128822 292170 128918 292226
rect 128298 292102 128918 292170
rect 128298 292046 128394 292102
rect 128450 292046 128518 292102
rect 128574 292046 128642 292102
rect 128698 292046 128766 292102
rect 128822 292046 128918 292102
rect 128298 291978 128918 292046
rect 128298 291922 128394 291978
rect 128450 291922 128518 291978
rect 128574 291922 128642 291978
rect 128698 291922 128766 291978
rect 128822 291922 128918 291978
rect 128298 274350 128918 291922
rect 128298 274294 128394 274350
rect 128450 274294 128518 274350
rect 128574 274294 128642 274350
rect 128698 274294 128766 274350
rect 128822 274294 128918 274350
rect 128298 274226 128918 274294
rect 128298 274170 128394 274226
rect 128450 274170 128518 274226
rect 128574 274170 128642 274226
rect 128698 274170 128766 274226
rect 128822 274170 128918 274226
rect 128298 274102 128918 274170
rect 128298 274046 128394 274102
rect 128450 274046 128518 274102
rect 128574 274046 128642 274102
rect 128698 274046 128766 274102
rect 128822 274046 128918 274102
rect 128298 273978 128918 274046
rect 128298 273922 128394 273978
rect 128450 273922 128518 273978
rect 128574 273922 128642 273978
rect 128698 273922 128766 273978
rect 128822 273922 128918 273978
rect 126812 72482 126868 72492
rect 126924 258244 126980 258254
rect 126924 60900 126980 258188
rect 128298 256350 128918 273922
rect 128298 256294 128394 256350
rect 128450 256294 128518 256350
rect 128574 256294 128642 256350
rect 128698 256294 128766 256350
rect 128822 256294 128918 256350
rect 128298 256226 128918 256294
rect 128298 256170 128394 256226
rect 128450 256170 128518 256226
rect 128574 256170 128642 256226
rect 128698 256170 128766 256226
rect 128822 256170 128918 256226
rect 128298 256102 128918 256170
rect 128298 256046 128394 256102
rect 128450 256046 128518 256102
rect 128574 256046 128642 256102
rect 128698 256046 128766 256102
rect 128822 256046 128918 256102
rect 128298 255978 128918 256046
rect 128298 255922 128394 255978
rect 128450 255922 128518 255978
rect 128574 255922 128642 255978
rect 128698 255922 128766 255978
rect 128822 255922 128918 255978
rect 128298 238350 128918 255922
rect 128298 238294 128394 238350
rect 128450 238294 128518 238350
rect 128574 238294 128642 238350
rect 128698 238294 128766 238350
rect 128822 238294 128918 238350
rect 128298 238226 128918 238294
rect 128298 238170 128394 238226
rect 128450 238170 128518 238226
rect 128574 238170 128642 238226
rect 128698 238170 128766 238226
rect 128822 238170 128918 238226
rect 128298 238102 128918 238170
rect 128298 238046 128394 238102
rect 128450 238046 128518 238102
rect 128574 238046 128642 238102
rect 128698 238046 128766 238102
rect 128822 238046 128918 238102
rect 128298 237978 128918 238046
rect 128298 237922 128394 237978
rect 128450 237922 128518 237978
rect 128574 237922 128642 237978
rect 128698 237922 128766 237978
rect 128822 237922 128918 237978
rect 128298 220350 128918 237922
rect 128298 220294 128394 220350
rect 128450 220294 128518 220350
rect 128574 220294 128642 220350
rect 128698 220294 128766 220350
rect 128822 220294 128918 220350
rect 128298 220226 128918 220294
rect 128298 220170 128394 220226
rect 128450 220170 128518 220226
rect 128574 220170 128642 220226
rect 128698 220170 128766 220226
rect 128822 220170 128918 220226
rect 128298 220102 128918 220170
rect 128298 220046 128394 220102
rect 128450 220046 128518 220102
rect 128574 220046 128642 220102
rect 128698 220046 128766 220102
rect 128822 220046 128918 220102
rect 128298 219978 128918 220046
rect 128298 219922 128394 219978
rect 128450 219922 128518 219978
rect 128574 219922 128642 219978
rect 128698 219922 128766 219978
rect 128822 219922 128918 219978
rect 126924 60834 126980 60844
rect 127036 218596 127092 218606
rect 126812 60004 126868 60014
rect 126028 45658 126084 45668
rect 123788 20132 124068 20188
rect 124012 10948 124068 20132
rect 124012 10882 124068 10892
rect 123452 6804 123508 6814
rect 123452 3332 123508 6748
rect 126028 4228 126084 45602
rect 126812 17220 126868 59948
rect 127036 52164 127092 218540
rect 128298 202350 128918 219922
rect 128298 202294 128394 202350
rect 128450 202294 128518 202350
rect 128574 202294 128642 202350
rect 128698 202294 128766 202350
rect 128822 202294 128918 202350
rect 128298 202226 128918 202294
rect 128298 202170 128394 202226
rect 128450 202170 128518 202226
rect 128574 202170 128642 202226
rect 128698 202170 128766 202226
rect 128822 202170 128918 202226
rect 128298 202102 128918 202170
rect 128298 202046 128394 202102
rect 128450 202046 128518 202102
rect 128574 202046 128642 202102
rect 128698 202046 128766 202102
rect 128822 202046 128918 202102
rect 128298 201978 128918 202046
rect 128298 201922 128394 201978
rect 128450 201922 128518 201978
rect 128574 201922 128642 201978
rect 128698 201922 128766 201978
rect 128822 201922 128918 201978
rect 128298 184350 128918 201922
rect 128298 184294 128394 184350
rect 128450 184294 128518 184350
rect 128574 184294 128642 184350
rect 128698 184294 128766 184350
rect 128822 184294 128918 184350
rect 128298 184226 128918 184294
rect 128298 184170 128394 184226
rect 128450 184170 128518 184226
rect 128574 184170 128642 184226
rect 128698 184170 128766 184226
rect 128822 184170 128918 184226
rect 128298 184102 128918 184170
rect 128298 184046 128394 184102
rect 128450 184046 128518 184102
rect 128574 184046 128642 184102
rect 128698 184046 128766 184102
rect 128822 184046 128918 184102
rect 128298 183978 128918 184046
rect 128298 183922 128394 183978
rect 128450 183922 128518 183978
rect 128574 183922 128642 183978
rect 128698 183922 128766 183978
rect 128822 183922 128918 183978
rect 127036 52098 127092 52108
rect 127148 178948 127204 178958
rect 127148 43428 127204 178892
rect 128298 166350 128918 183922
rect 128298 166294 128394 166350
rect 128450 166294 128518 166350
rect 128574 166294 128642 166350
rect 128698 166294 128766 166350
rect 128822 166294 128918 166350
rect 128298 166226 128918 166294
rect 128298 166170 128394 166226
rect 128450 166170 128518 166226
rect 128574 166170 128642 166226
rect 128698 166170 128766 166226
rect 128822 166170 128918 166226
rect 128298 166102 128918 166170
rect 128298 166046 128394 166102
rect 128450 166046 128518 166102
rect 128574 166046 128642 166102
rect 128698 166046 128766 166102
rect 128822 166046 128918 166102
rect 128298 165978 128918 166046
rect 128298 165922 128394 165978
rect 128450 165922 128518 165978
rect 128574 165922 128642 165978
rect 128698 165922 128766 165978
rect 128822 165922 128918 165978
rect 128298 148350 128918 165922
rect 128298 148294 128394 148350
rect 128450 148294 128518 148350
rect 128574 148294 128642 148350
rect 128698 148294 128766 148350
rect 128822 148294 128918 148350
rect 128298 148226 128918 148294
rect 128298 148170 128394 148226
rect 128450 148170 128518 148226
rect 128574 148170 128642 148226
rect 128698 148170 128766 148226
rect 128822 148170 128918 148226
rect 128298 148102 128918 148170
rect 128298 148046 128394 148102
rect 128450 148046 128518 148102
rect 128574 148046 128642 148102
rect 128698 148046 128766 148102
rect 128822 148046 128918 148102
rect 128298 147978 128918 148046
rect 128298 147922 128394 147978
rect 128450 147922 128518 147978
rect 128574 147922 128642 147978
rect 128698 147922 128766 147978
rect 128822 147922 128918 147978
rect 127148 43362 127204 43372
rect 127260 139300 127316 139310
rect 127260 34692 127316 139244
rect 128298 130350 128918 147922
rect 128298 130294 128394 130350
rect 128450 130294 128518 130350
rect 128574 130294 128642 130350
rect 128698 130294 128766 130350
rect 128822 130294 128918 130350
rect 128298 130226 128918 130294
rect 128298 130170 128394 130226
rect 128450 130170 128518 130226
rect 128574 130170 128642 130226
rect 128698 130170 128766 130226
rect 128822 130170 128918 130226
rect 128298 130102 128918 130170
rect 128298 130046 128394 130102
rect 128450 130046 128518 130102
rect 128574 130046 128642 130102
rect 128698 130046 128766 130102
rect 128822 130046 128918 130102
rect 128298 129978 128918 130046
rect 128298 129922 128394 129978
rect 128450 129922 128518 129978
rect 128574 129922 128642 129978
rect 128698 129922 128766 129978
rect 128822 129922 128918 129978
rect 128298 112350 128918 129922
rect 132018 598172 132638 598268
rect 132018 598116 132114 598172
rect 132170 598116 132238 598172
rect 132294 598116 132362 598172
rect 132418 598116 132486 598172
rect 132542 598116 132638 598172
rect 132018 598048 132638 598116
rect 132018 597992 132114 598048
rect 132170 597992 132238 598048
rect 132294 597992 132362 598048
rect 132418 597992 132486 598048
rect 132542 597992 132638 598048
rect 132018 597924 132638 597992
rect 132018 597868 132114 597924
rect 132170 597868 132238 597924
rect 132294 597868 132362 597924
rect 132418 597868 132486 597924
rect 132542 597868 132638 597924
rect 132018 597800 132638 597868
rect 132018 597744 132114 597800
rect 132170 597744 132238 597800
rect 132294 597744 132362 597800
rect 132418 597744 132486 597800
rect 132542 597744 132638 597800
rect 132018 586350 132638 597744
rect 132018 586294 132114 586350
rect 132170 586294 132238 586350
rect 132294 586294 132362 586350
rect 132418 586294 132486 586350
rect 132542 586294 132638 586350
rect 132018 586226 132638 586294
rect 132018 586170 132114 586226
rect 132170 586170 132238 586226
rect 132294 586170 132362 586226
rect 132418 586170 132486 586226
rect 132542 586170 132638 586226
rect 132018 586102 132638 586170
rect 132018 586046 132114 586102
rect 132170 586046 132238 586102
rect 132294 586046 132362 586102
rect 132418 586046 132486 586102
rect 132542 586046 132638 586102
rect 132018 585978 132638 586046
rect 132018 585922 132114 585978
rect 132170 585922 132238 585978
rect 132294 585922 132362 585978
rect 132418 585922 132486 585978
rect 132542 585922 132638 585978
rect 132018 568350 132638 585922
rect 132018 568294 132114 568350
rect 132170 568294 132238 568350
rect 132294 568294 132362 568350
rect 132418 568294 132486 568350
rect 132542 568294 132638 568350
rect 132018 568226 132638 568294
rect 132018 568170 132114 568226
rect 132170 568170 132238 568226
rect 132294 568170 132362 568226
rect 132418 568170 132486 568226
rect 132542 568170 132638 568226
rect 132018 568102 132638 568170
rect 132018 568046 132114 568102
rect 132170 568046 132238 568102
rect 132294 568046 132362 568102
rect 132418 568046 132486 568102
rect 132542 568046 132638 568102
rect 132018 567978 132638 568046
rect 132018 567922 132114 567978
rect 132170 567922 132238 567978
rect 132294 567922 132362 567978
rect 132418 567922 132486 567978
rect 132542 567922 132638 567978
rect 132018 550350 132638 567922
rect 132018 550294 132114 550350
rect 132170 550294 132238 550350
rect 132294 550294 132362 550350
rect 132418 550294 132486 550350
rect 132542 550294 132638 550350
rect 132018 550226 132638 550294
rect 132018 550170 132114 550226
rect 132170 550170 132238 550226
rect 132294 550170 132362 550226
rect 132418 550170 132486 550226
rect 132542 550170 132638 550226
rect 132018 550102 132638 550170
rect 132018 550046 132114 550102
rect 132170 550046 132238 550102
rect 132294 550046 132362 550102
rect 132418 550046 132486 550102
rect 132542 550046 132638 550102
rect 132018 549978 132638 550046
rect 132018 549922 132114 549978
rect 132170 549922 132238 549978
rect 132294 549922 132362 549978
rect 132418 549922 132486 549978
rect 132542 549922 132638 549978
rect 132018 532350 132638 549922
rect 132018 532294 132114 532350
rect 132170 532294 132238 532350
rect 132294 532294 132362 532350
rect 132418 532294 132486 532350
rect 132542 532294 132638 532350
rect 132018 532226 132638 532294
rect 132018 532170 132114 532226
rect 132170 532170 132238 532226
rect 132294 532170 132362 532226
rect 132418 532170 132486 532226
rect 132542 532170 132638 532226
rect 132018 532102 132638 532170
rect 132018 532046 132114 532102
rect 132170 532046 132238 532102
rect 132294 532046 132362 532102
rect 132418 532046 132486 532102
rect 132542 532046 132638 532102
rect 132018 531978 132638 532046
rect 132018 531922 132114 531978
rect 132170 531922 132238 531978
rect 132294 531922 132362 531978
rect 132418 531922 132486 531978
rect 132542 531922 132638 531978
rect 132018 514350 132638 531922
rect 132018 514294 132114 514350
rect 132170 514294 132238 514350
rect 132294 514294 132362 514350
rect 132418 514294 132486 514350
rect 132542 514294 132638 514350
rect 132018 514226 132638 514294
rect 132018 514170 132114 514226
rect 132170 514170 132238 514226
rect 132294 514170 132362 514226
rect 132418 514170 132486 514226
rect 132542 514170 132638 514226
rect 132018 514102 132638 514170
rect 132018 514046 132114 514102
rect 132170 514046 132238 514102
rect 132294 514046 132362 514102
rect 132418 514046 132486 514102
rect 132542 514046 132638 514102
rect 132018 513978 132638 514046
rect 132018 513922 132114 513978
rect 132170 513922 132238 513978
rect 132294 513922 132362 513978
rect 132418 513922 132486 513978
rect 132542 513922 132638 513978
rect 132018 496350 132638 513922
rect 132018 496294 132114 496350
rect 132170 496294 132238 496350
rect 132294 496294 132362 496350
rect 132418 496294 132486 496350
rect 132542 496294 132638 496350
rect 132018 496226 132638 496294
rect 132018 496170 132114 496226
rect 132170 496170 132238 496226
rect 132294 496170 132362 496226
rect 132418 496170 132486 496226
rect 132542 496170 132638 496226
rect 132018 496102 132638 496170
rect 132018 496046 132114 496102
rect 132170 496046 132238 496102
rect 132294 496046 132362 496102
rect 132418 496046 132486 496102
rect 132542 496046 132638 496102
rect 132018 495978 132638 496046
rect 132018 495922 132114 495978
rect 132170 495922 132238 495978
rect 132294 495922 132362 495978
rect 132418 495922 132486 495978
rect 132542 495922 132638 495978
rect 132018 478350 132638 495922
rect 132018 478294 132114 478350
rect 132170 478294 132238 478350
rect 132294 478294 132362 478350
rect 132418 478294 132486 478350
rect 132542 478294 132638 478350
rect 132018 478226 132638 478294
rect 132018 478170 132114 478226
rect 132170 478170 132238 478226
rect 132294 478170 132362 478226
rect 132418 478170 132486 478226
rect 132542 478170 132638 478226
rect 132018 478102 132638 478170
rect 132018 478046 132114 478102
rect 132170 478046 132238 478102
rect 132294 478046 132362 478102
rect 132418 478046 132486 478102
rect 132542 478046 132638 478102
rect 132018 477978 132638 478046
rect 132018 477922 132114 477978
rect 132170 477922 132238 477978
rect 132294 477922 132362 477978
rect 132418 477922 132486 477978
rect 132542 477922 132638 477978
rect 132018 460350 132638 477922
rect 132018 460294 132114 460350
rect 132170 460294 132238 460350
rect 132294 460294 132362 460350
rect 132418 460294 132486 460350
rect 132542 460294 132638 460350
rect 132018 460226 132638 460294
rect 132018 460170 132114 460226
rect 132170 460170 132238 460226
rect 132294 460170 132362 460226
rect 132418 460170 132486 460226
rect 132542 460170 132638 460226
rect 132018 460102 132638 460170
rect 132018 460046 132114 460102
rect 132170 460046 132238 460102
rect 132294 460046 132362 460102
rect 132418 460046 132486 460102
rect 132542 460046 132638 460102
rect 132018 459978 132638 460046
rect 132018 459922 132114 459978
rect 132170 459922 132238 459978
rect 132294 459922 132362 459978
rect 132418 459922 132486 459978
rect 132542 459922 132638 459978
rect 132018 442350 132638 459922
rect 132018 442294 132114 442350
rect 132170 442294 132238 442350
rect 132294 442294 132362 442350
rect 132418 442294 132486 442350
rect 132542 442294 132638 442350
rect 132018 442226 132638 442294
rect 132018 442170 132114 442226
rect 132170 442170 132238 442226
rect 132294 442170 132362 442226
rect 132418 442170 132486 442226
rect 132542 442170 132638 442226
rect 132018 442102 132638 442170
rect 132018 442046 132114 442102
rect 132170 442046 132238 442102
rect 132294 442046 132362 442102
rect 132418 442046 132486 442102
rect 132542 442046 132638 442102
rect 132018 441978 132638 442046
rect 132018 441922 132114 441978
rect 132170 441922 132238 441978
rect 132294 441922 132362 441978
rect 132418 441922 132486 441978
rect 132542 441922 132638 441978
rect 132018 424350 132638 441922
rect 132018 424294 132114 424350
rect 132170 424294 132238 424350
rect 132294 424294 132362 424350
rect 132418 424294 132486 424350
rect 132542 424294 132638 424350
rect 132018 424226 132638 424294
rect 132018 424170 132114 424226
rect 132170 424170 132238 424226
rect 132294 424170 132362 424226
rect 132418 424170 132486 424226
rect 132542 424170 132638 424226
rect 132018 424102 132638 424170
rect 132018 424046 132114 424102
rect 132170 424046 132238 424102
rect 132294 424046 132362 424102
rect 132418 424046 132486 424102
rect 132542 424046 132638 424102
rect 132018 423978 132638 424046
rect 132018 423922 132114 423978
rect 132170 423922 132238 423978
rect 132294 423922 132362 423978
rect 132418 423922 132486 423978
rect 132542 423922 132638 423978
rect 132018 406350 132638 423922
rect 132018 406294 132114 406350
rect 132170 406294 132238 406350
rect 132294 406294 132362 406350
rect 132418 406294 132486 406350
rect 132542 406294 132638 406350
rect 132018 406226 132638 406294
rect 132018 406170 132114 406226
rect 132170 406170 132238 406226
rect 132294 406170 132362 406226
rect 132418 406170 132486 406226
rect 132542 406170 132638 406226
rect 132018 406102 132638 406170
rect 132018 406046 132114 406102
rect 132170 406046 132238 406102
rect 132294 406046 132362 406102
rect 132418 406046 132486 406102
rect 132542 406046 132638 406102
rect 132018 405978 132638 406046
rect 132018 405922 132114 405978
rect 132170 405922 132238 405978
rect 132294 405922 132362 405978
rect 132418 405922 132486 405978
rect 132542 405922 132638 405978
rect 132018 388350 132638 405922
rect 132018 388294 132114 388350
rect 132170 388294 132238 388350
rect 132294 388294 132362 388350
rect 132418 388294 132486 388350
rect 132542 388294 132638 388350
rect 132018 388226 132638 388294
rect 132018 388170 132114 388226
rect 132170 388170 132238 388226
rect 132294 388170 132362 388226
rect 132418 388170 132486 388226
rect 132542 388170 132638 388226
rect 132018 388102 132638 388170
rect 132018 388046 132114 388102
rect 132170 388046 132238 388102
rect 132294 388046 132362 388102
rect 132418 388046 132486 388102
rect 132542 388046 132638 388102
rect 132018 387978 132638 388046
rect 132018 387922 132114 387978
rect 132170 387922 132238 387978
rect 132294 387922 132362 387978
rect 132418 387922 132486 387978
rect 132542 387922 132638 387978
rect 132018 370350 132638 387922
rect 132018 370294 132114 370350
rect 132170 370294 132238 370350
rect 132294 370294 132362 370350
rect 132418 370294 132486 370350
rect 132542 370294 132638 370350
rect 132018 370226 132638 370294
rect 132018 370170 132114 370226
rect 132170 370170 132238 370226
rect 132294 370170 132362 370226
rect 132418 370170 132486 370226
rect 132542 370170 132638 370226
rect 132018 370102 132638 370170
rect 132018 370046 132114 370102
rect 132170 370046 132238 370102
rect 132294 370046 132362 370102
rect 132418 370046 132486 370102
rect 132542 370046 132638 370102
rect 132018 369978 132638 370046
rect 132018 369922 132114 369978
rect 132170 369922 132238 369978
rect 132294 369922 132362 369978
rect 132418 369922 132486 369978
rect 132542 369922 132638 369978
rect 132018 352350 132638 369922
rect 132018 352294 132114 352350
rect 132170 352294 132238 352350
rect 132294 352294 132362 352350
rect 132418 352294 132486 352350
rect 132542 352294 132638 352350
rect 132018 352226 132638 352294
rect 132018 352170 132114 352226
rect 132170 352170 132238 352226
rect 132294 352170 132362 352226
rect 132418 352170 132486 352226
rect 132542 352170 132638 352226
rect 132018 352102 132638 352170
rect 132018 352046 132114 352102
rect 132170 352046 132238 352102
rect 132294 352046 132362 352102
rect 132418 352046 132486 352102
rect 132542 352046 132638 352102
rect 132018 351978 132638 352046
rect 132018 351922 132114 351978
rect 132170 351922 132238 351978
rect 132294 351922 132362 351978
rect 132418 351922 132486 351978
rect 132542 351922 132638 351978
rect 132018 334350 132638 351922
rect 132018 334294 132114 334350
rect 132170 334294 132238 334350
rect 132294 334294 132362 334350
rect 132418 334294 132486 334350
rect 132542 334294 132638 334350
rect 132018 334226 132638 334294
rect 132018 334170 132114 334226
rect 132170 334170 132238 334226
rect 132294 334170 132362 334226
rect 132418 334170 132486 334226
rect 132542 334170 132638 334226
rect 132018 334102 132638 334170
rect 132018 334046 132114 334102
rect 132170 334046 132238 334102
rect 132294 334046 132362 334102
rect 132418 334046 132486 334102
rect 132542 334046 132638 334102
rect 132018 333978 132638 334046
rect 132018 333922 132114 333978
rect 132170 333922 132238 333978
rect 132294 333922 132362 333978
rect 132418 333922 132486 333978
rect 132542 333922 132638 333978
rect 132018 316350 132638 333922
rect 132018 316294 132114 316350
rect 132170 316294 132238 316350
rect 132294 316294 132362 316350
rect 132418 316294 132486 316350
rect 132542 316294 132638 316350
rect 132018 316226 132638 316294
rect 132018 316170 132114 316226
rect 132170 316170 132238 316226
rect 132294 316170 132362 316226
rect 132418 316170 132486 316226
rect 132542 316170 132638 316226
rect 132018 316102 132638 316170
rect 132018 316046 132114 316102
rect 132170 316046 132238 316102
rect 132294 316046 132362 316102
rect 132418 316046 132486 316102
rect 132542 316046 132638 316102
rect 132018 315978 132638 316046
rect 132018 315922 132114 315978
rect 132170 315922 132238 315978
rect 132294 315922 132362 315978
rect 132418 315922 132486 315978
rect 132542 315922 132638 315978
rect 132018 298350 132638 315922
rect 132018 298294 132114 298350
rect 132170 298294 132238 298350
rect 132294 298294 132362 298350
rect 132418 298294 132486 298350
rect 132542 298294 132638 298350
rect 132018 298226 132638 298294
rect 132018 298170 132114 298226
rect 132170 298170 132238 298226
rect 132294 298170 132362 298226
rect 132418 298170 132486 298226
rect 132542 298170 132638 298226
rect 132018 298102 132638 298170
rect 132018 298046 132114 298102
rect 132170 298046 132238 298102
rect 132294 298046 132362 298102
rect 132418 298046 132486 298102
rect 132542 298046 132638 298102
rect 132018 297978 132638 298046
rect 132018 297922 132114 297978
rect 132170 297922 132238 297978
rect 132294 297922 132362 297978
rect 132418 297922 132486 297978
rect 132542 297922 132638 297978
rect 132018 280350 132638 297922
rect 159018 597212 159638 598268
rect 159018 597156 159114 597212
rect 159170 597156 159238 597212
rect 159294 597156 159362 597212
rect 159418 597156 159486 597212
rect 159542 597156 159638 597212
rect 159018 597088 159638 597156
rect 159018 597032 159114 597088
rect 159170 597032 159238 597088
rect 159294 597032 159362 597088
rect 159418 597032 159486 597088
rect 159542 597032 159638 597088
rect 159018 596964 159638 597032
rect 159018 596908 159114 596964
rect 159170 596908 159238 596964
rect 159294 596908 159362 596964
rect 159418 596908 159486 596964
rect 159542 596908 159638 596964
rect 159018 596840 159638 596908
rect 159018 596784 159114 596840
rect 159170 596784 159238 596840
rect 159294 596784 159362 596840
rect 159418 596784 159486 596840
rect 159542 596784 159638 596840
rect 159018 580350 159638 596784
rect 159018 580294 159114 580350
rect 159170 580294 159238 580350
rect 159294 580294 159362 580350
rect 159418 580294 159486 580350
rect 159542 580294 159638 580350
rect 159018 580226 159638 580294
rect 159018 580170 159114 580226
rect 159170 580170 159238 580226
rect 159294 580170 159362 580226
rect 159418 580170 159486 580226
rect 159542 580170 159638 580226
rect 159018 580102 159638 580170
rect 159018 580046 159114 580102
rect 159170 580046 159238 580102
rect 159294 580046 159362 580102
rect 159418 580046 159486 580102
rect 159542 580046 159638 580102
rect 159018 579978 159638 580046
rect 159018 579922 159114 579978
rect 159170 579922 159238 579978
rect 159294 579922 159362 579978
rect 159418 579922 159486 579978
rect 159542 579922 159638 579978
rect 159018 562350 159638 579922
rect 159018 562294 159114 562350
rect 159170 562294 159238 562350
rect 159294 562294 159362 562350
rect 159418 562294 159486 562350
rect 159542 562294 159638 562350
rect 159018 562226 159638 562294
rect 159018 562170 159114 562226
rect 159170 562170 159238 562226
rect 159294 562170 159362 562226
rect 159418 562170 159486 562226
rect 159542 562170 159638 562226
rect 159018 562102 159638 562170
rect 159018 562046 159114 562102
rect 159170 562046 159238 562102
rect 159294 562046 159362 562102
rect 159418 562046 159486 562102
rect 159542 562046 159638 562102
rect 159018 561978 159638 562046
rect 159018 561922 159114 561978
rect 159170 561922 159238 561978
rect 159294 561922 159362 561978
rect 159418 561922 159486 561978
rect 159542 561922 159638 561978
rect 159018 544350 159638 561922
rect 159018 544294 159114 544350
rect 159170 544294 159238 544350
rect 159294 544294 159362 544350
rect 159418 544294 159486 544350
rect 159542 544294 159638 544350
rect 159018 544226 159638 544294
rect 159018 544170 159114 544226
rect 159170 544170 159238 544226
rect 159294 544170 159362 544226
rect 159418 544170 159486 544226
rect 159542 544170 159638 544226
rect 159018 544102 159638 544170
rect 159018 544046 159114 544102
rect 159170 544046 159238 544102
rect 159294 544046 159362 544102
rect 159418 544046 159486 544102
rect 159542 544046 159638 544102
rect 159018 543978 159638 544046
rect 159018 543922 159114 543978
rect 159170 543922 159238 543978
rect 159294 543922 159362 543978
rect 159418 543922 159486 543978
rect 159542 543922 159638 543978
rect 159018 526350 159638 543922
rect 159018 526294 159114 526350
rect 159170 526294 159238 526350
rect 159294 526294 159362 526350
rect 159418 526294 159486 526350
rect 159542 526294 159638 526350
rect 159018 526226 159638 526294
rect 159018 526170 159114 526226
rect 159170 526170 159238 526226
rect 159294 526170 159362 526226
rect 159418 526170 159486 526226
rect 159542 526170 159638 526226
rect 159018 526102 159638 526170
rect 159018 526046 159114 526102
rect 159170 526046 159238 526102
rect 159294 526046 159362 526102
rect 159418 526046 159486 526102
rect 159542 526046 159638 526102
rect 159018 525978 159638 526046
rect 159018 525922 159114 525978
rect 159170 525922 159238 525978
rect 159294 525922 159362 525978
rect 159418 525922 159486 525978
rect 159542 525922 159638 525978
rect 159018 508350 159638 525922
rect 159018 508294 159114 508350
rect 159170 508294 159238 508350
rect 159294 508294 159362 508350
rect 159418 508294 159486 508350
rect 159542 508294 159638 508350
rect 159018 508226 159638 508294
rect 159018 508170 159114 508226
rect 159170 508170 159238 508226
rect 159294 508170 159362 508226
rect 159418 508170 159486 508226
rect 159542 508170 159638 508226
rect 159018 508102 159638 508170
rect 159018 508046 159114 508102
rect 159170 508046 159238 508102
rect 159294 508046 159362 508102
rect 159418 508046 159486 508102
rect 159542 508046 159638 508102
rect 159018 507978 159638 508046
rect 159018 507922 159114 507978
rect 159170 507922 159238 507978
rect 159294 507922 159362 507978
rect 159418 507922 159486 507978
rect 159542 507922 159638 507978
rect 159018 490350 159638 507922
rect 159018 490294 159114 490350
rect 159170 490294 159238 490350
rect 159294 490294 159362 490350
rect 159418 490294 159486 490350
rect 159542 490294 159638 490350
rect 159018 490226 159638 490294
rect 159018 490170 159114 490226
rect 159170 490170 159238 490226
rect 159294 490170 159362 490226
rect 159418 490170 159486 490226
rect 159542 490170 159638 490226
rect 159018 490102 159638 490170
rect 159018 490046 159114 490102
rect 159170 490046 159238 490102
rect 159294 490046 159362 490102
rect 159418 490046 159486 490102
rect 159542 490046 159638 490102
rect 159018 489978 159638 490046
rect 159018 489922 159114 489978
rect 159170 489922 159238 489978
rect 159294 489922 159362 489978
rect 159418 489922 159486 489978
rect 159542 489922 159638 489978
rect 159018 472350 159638 489922
rect 159018 472294 159114 472350
rect 159170 472294 159238 472350
rect 159294 472294 159362 472350
rect 159418 472294 159486 472350
rect 159542 472294 159638 472350
rect 159018 472226 159638 472294
rect 159018 472170 159114 472226
rect 159170 472170 159238 472226
rect 159294 472170 159362 472226
rect 159418 472170 159486 472226
rect 159542 472170 159638 472226
rect 159018 472102 159638 472170
rect 159018 472046 159114 472102
rect 159170 472046 159238 472102
rect 159294 472046 159362 472102
rect 159418 472046 159486 472102
rect 159542 472046 159638 472102
rect 159018 471978 159638 472046
rect 159018 471922 159114 471978
rect 159170 471922 159238 471978
rect 159294 471922 159362 471978
rect 159418 471922 159486 471978
rect 159542 471922 159638 471978
rect 159018 454350 159638 471922
rect 159018 454294 159114 454350
rect 159170 454294 159238 454350
rect 159294 454294 159362 454350
rect 159418 454294 159486 454350
rect 159542 454294 159638 454350
rect 159018 454226 159638 454294
rect 159018 454170 159114 454226
rect 159170 454170 159238 454226
rect 159294 454170 159362 454226
rect 159418 454170 159486 454226
rect 159542 454170 159638 454226
rect 159018 454102 159638 454170
rect 159018 454046 159114 454102
rect 159170 454046 159238 454102
rect 159294 454046 159362 454102
rect 159418 454046 159486 454102
rect 159542 454046 159638 454102
rect 159018 453978 159638 454046
rect 159018 453922 159114 453978
rect 159170 453922 159238 453978
rect 159294 453922 159362 453978
rect 159418 453922 159486 453978
rect 159542 453922 159638 453978
rect 159018 436350 159638 453922
rect 159018 436294 159114 436350
rect 159170 436294 159238 436350
rect 159294 436294 159362 436350
rect 159418 436294 159486 436350
rect 159542 436294 159638 436350
rect 159018 436226 159638 436294
rect 159018 436170 159114 436226
rect 159170 436170 159238 436226
rect 159294 436170 159362 436226
rect 159418 436170 159486 436226
rect 159542 436170 159638 436226
rect 159018 436102 159638 436170
rect 159018 436046 159114 436102
rect 159170 436046 159238 436102
rect 159294 436046 159362 436102
rect 159418 436046 159486 436102
rect 159542 436046 159638 436102
rect 159018 435978 159638 436046
rect 159018 435922 159114 435978
rect 159170 435922 159238 435978
rect 159294 435922 159362 435978
rect 159418 435922 159486 435978
rect 159542 435922 159638 435978
rect 159018 418350 159638 435922
rect 159018 418294 159114 418350
rect 159170 418294 159238 418350
rect 159294 418294 159362 418350
rect 159418 418294 159486 418350
rect 159542 418294 159638 418350
rect 159018 418226 159638 418294
rect 159018 418170 159114 418226
rect 159170 418170 159238 418226
rect 159294 418170 159362 418226
rect 159418 418170 159486 418226
rect 159542 418170 159638 418226
rect 159018 418102 159638 418170
rect 159018 418046 159114 418102
rect 159170 418046 159238 418102
rect 159294 418046 159362 418102
rect 159418 418046 159486 418102
rect 159542 418046 159638 418102
rect 159018 417978 159638 418046
rect 159018 417922 159114 417978
rect 159170 417922 159238 417978
rect 159294 417922 159362 417978
rect 159418 417922 159486 417978
rect 159542 417922 159638 417978
rect 159018 400350 159638 417922
rect 159018 400294 159114 400350
rect 159170 400294 159238 400350
rect 159294 400294 159362 400350
rect 159418 400294 159486 400350
rect 159542 400294 159638 400350
rect 159018 400226 159638 400294
rect 159018 400170 159114 400226
rect 159170 400170 159238 400226
rect 159294 400170 159362 400226
rect 159418 400170 159486 400226
rect 159542 400170 159638 400226
rect 159018 400102 159638 400170
rect 159018 400046 159114 400102
rect 159170 400046 159238 400102
rect 159294 400046 159362 400102
rect 159418 400046 159486 400102
rect 159542 400046 159638 400102
rect 159018 399978 159638 400046
rect 159018 399922 159114 399978
rect 159170 399922 159238 399978
rect 159294 399922 159362 399978
rect 159418 399922 159486 399978
rect 159542 399922 159638 399978
rect 159018 382350 159638 399922
rect 159018 382294 159114 382350
rect 159170 382294 159238 382350
rect 159294 382294 159362 382350
rect 159418 382294 159486 382350
rect 159542 382294 159638 382350
rect 159018 382226 159638 382294
rect 159018 382170 159114 382226
rect 159170 382170 159238 382226
rect 159294 382170 159362 382226
rect 159418 382170 159486 382226
rect 159542 382170 159638 382226
rect 159018 382102 159638 382170
rect 159018 382046 159114 382102
rect 159170 382046 159238 382102
rect 159294 382046 159362 382102
rect 159418 382046 159486 382102
rect 159542 382046 159638 382102
rect 159018 381978 159638 382046
rect 159018 381922 159114 381978
rect 159170 381922 159238 381978
rect 159294 381922 159362 381978
rect 159418 381922 159486 381978
rect 159542 381922 159638 381978
rect 159018 364350 159638 381922
rect 159018 364294 159114 364350
rect 159170 364294 159238 364350
rect 159294 364294 159362 364350
rect 159418 364294 159486 364350
rect 159542 364294 159638 364350
rect 159018 364226 159638 364294
rect 159018 364170 159114 364226
rect 159170 364170 159238 364226
rect 159294 364170 159362 364226
rect 159418 364170 159486 364226
rect 159542 364170 159638 364226
rect 159018 364102 159638 364170
rect 159018 364046 159114 364102
rect 159170 364046 159238 364102
rect 159294 364046 159362 364102
rect 159418 364046 159486 364102
rect 159542 364046 159638 364102
rect 159018 363978 159638 364046
rect 159018 363922 159114 363978
rect 159170 363922 159238 363978
rect 159294 363922 159362 363978
rect 159418 363922 159486 363978
rect 159542 363922 159638 363978
rect 159018 346350 159638 363922
rect 159018 346294 159114 346350
rect 159170 346294 159238 346350
rect 159294 346294 159362 346350
rect 159418 346294 159486 346350
rect 159542 346294 159638 346350
rect 159018 346226 159638 346294
rect 159018 346170 159114 346226
rect 159170 346170 159238 346226
rect 159294 346170 159362 346226
rect 159418 346170 159486 346226
rect 159542 346170 159638 346226
rect 159018 346102 159638 346170
rect 159018 346046 159114 346102
rect 159170 346046 159238 346102
rect 159294 346046 159362 346102
rect 159418 346046 159486 346102
rect 159542 346046 159638 346102
rect 159018 345978 159638 346046
rect 159018 345922 159114 345978
rect 159170 345922 159238 345978
rect 159294 345922 159362 345978
rect 159418 345922 159486 345978
rect 159542 345922 159638 345978
rect 159018 328350 159638 345922
rect 159018 328294 159114 328350
rect 159170 328294 159238 328350
rect 159294 328294 159362 328350
rect 159418 328294 159486 328350
rect 159542 328294 159638 328350
rect 159018 328226 159638 328294
rect 159018 328170 159114 328226
rect 159170 328170 159238 328226
rect 159294 328170 159362 328226
rect 159418 328170 159486 328226
rect 159542 328170 159638 328226
rect 159018 328102 159638 328170
rect 159018 328046 159114 328102
rect 159170 328046 159238 328102
rect 159294 328046 159362 328102
rect 159418 328046 159486 328102
rect 159542 328046 159638 328102
rect 159018 327978 159638 328046
rect 159018 327922 159114 327978
rect 159170 327922 159238 327978
rect 159294 327922 159362 327978
rect 159418 327922 159486 327978
rect 159542 327922 159638 327978
rect 159018 310350 159638 327922
rect 159018 310294 159114 310350
rect 159170 310294 159238 310350
rect 159294 310294 159362 310350
rect 159418 310294 159486 310350
rect 159542 310294 159638 310350
rect 159018 310226 159638 310294
rect 159018 310170 159114 310226
rect 159170 310170 159238 310226
rect 159294 310170 159362 310226
rect 159418 310170 159486 310226
rect 159542 310170 159638 310226
rect 159018 310102 159638 310170
rect 159018 310046 159114 310102
rect 159170 310046 159238 310102
rect 159294 310046 159362 310102
rect 159418 310046 159486 310102
rect 159542 310046 159638 310102
rect 159018 309978 159638 310046
rect 159018 309922 159114 309978
rect 159170 309922 159238 309978
rect 159294 309922 159362 309978
rect 159418 309922 159486 309978
rect 159542 309922 159638 309978
rect 132018 280294 132114 280350
rect 132170 280294 132238 280350
rect 132294 280294 132362 280350
rect 132418 280294 132486 280350
rect 132542 280294 132638 280350
rect 132018 280226 132638 280294
rect 132018 280170 132114 280226
rect 132170 280170 132238 280226
rect 132294 280170 132362 280226
rect 132418 280170 132486 280226
rect 132542 280170 132638 280226
rect 132018 280102 132638 280170
rect 132018 280046 132114 280102
rect 132170 280046 132238 280102
rect 132294 280046 132362 280102
rect 132418 280046 132486 280102
rect 132542 280046 132638 280102
rect 132018 279978 132638 280046
rect 132018 279922 132114 279978
rect 132170 279922 132238 279978
rect 132294 279922 132362 279978
rect 132418 279922 132486 279978
rect 132542 279922 132638 279978
rect 132018 262350 132638 279922
rect 150332 296548 150388 296558
rect 132018 262294 132114 262350
rect 132170 262294 132238 262350
rect 132294 262294 132362 262350
rect 132418 262294 132486 262350
rect 132542 262294 132638 262350
rect 132018 262226 132638 262294
rect 132018 262170 132114 262226
rect 132170 262170 132238 262226
rect 132294 262170 132362 262226
rect 132418 262170 132486 262226
rect 132542 262170 132638 262226
rect 132018 262102 132638 262170
rect 132018 262046 132114 262102
rect 132170 262046 132238 262102
rect 132294 262046 132362 262102
rect 132418 262046 132486 262102
rect 132542 262046 132638 262102
rect 132018 261978 132638 262046
rect 132018 261922 132114 261978
rect 132170 261922 132238 261978
rect 132294 261922 132362 261978
rect 132418 261922 132486 261978
rect 132542 261922 132638 261978
rect 132018 244350 132638 261922
rect 132018 244294 132114 244350
rect 132170 244294 132238 244350
rect 132294 244294 132362 244350
rect 132418 244294 132486 244350
rect 132542 244294 132638 244350
rect 132018 244226 132638 244294
rect 132018 244170 132114 244226
rect 132170 244170 132238 244226
rect 132294 244170 132362 244226
rect 132418 244170 132486 244226
rect 132542 244170 132638 244226
rect 132018 244102 132638 244170
rect 132018 244046 132114 244102
rect 132170 244046 132238 244102
rect 132294 244046 132362 244102
rect 132418 244046 132486 244102
rect 132542 244046 132638 244102
rect 132018 243978 132638 244046
rect 132018 243922 132114 243978
rect 132170 243922 132238 243978
rect 132294 243922 132362 243978
rect 132418 243922 132486 243978
rect 132542 243922 132638 243978
rect 132018 226350 132638 243922
rect 145292 271460 145348 271470
rect 132018 226294 132114 226350
rect 132170 226294 132238 226350
rect 132294 226294 132362 226350
rect 132418 226294 132486 226350
rect 132542 226294 132638 226350
rect 132018 226226 132638 226294
rect 132018 226170 132114 226226
rect 132170 226170 132238 226226
rect 132294 226170 132362 226226
rect 132418 226170 132486 226226
rect 132542 226170 132638 226226
rect 132018 226102 132638 226170
rect 132018 226046 132114 226102
rect 132170 226046 132238 226102
rect 132294 226046 132362 226102
rect 132418 226046 132486 226102
rect 132542 226046 132638 226102
rect 132018 225978 132638 226046
rect 132018 225922 132114 225978
rect 132170 225922 132238 225978
rect 132294 225922 132362 225978
rect 132418 225922 132486 225978
rect 132542 225922 132638 225978
rect 132018 208350 132638 225922
rect 132018 208294 132114 208350
rect 132170 208294 132238 208350
rect 132294 208294 132362 208350
rect 132418 208294 132486 208350
rect 132542 208294 132638 208350
rect 132018 208226 132638 208294
rect 132018 208170 132114 208226
rect 132170 208170 132238 208226
rect 132294 208170 132362 208226
rect 132418 208170 132486 208226
rect 132542 208170 132638 208226
rect 132018 208102 132638 208170
rect 132018 208046 132114 208102
rect 132170 208046 132238 208102
rect 132294 208046 132362 208102
rect 132418 208046 132486 208102
rect 132542 208046 132638 208102
rect 132018 207978 132638 208046
rect 132018 207922 132114 207978
rect 132170 207922 132238 207978
rect 132294 207922 132362 207978
rect 132418 207922 132486 207978
rect 132542 207922 132638 207978
rect 132018 190350 132638 207922
rect 136892 242788 136948 242798
rect 132018 190294 132114 190350
rect 132170 190294 132238 190350
rect 132294 190294 132362 190350
rect 132418 190294 132486 190350
rect 132542 190294 132638 190350
rect 132018 190226 132638 190294
rect 132018 190170 132114 190226
rect 132170 190170 132238 190226
rect 132294 190170 132362 190226
rect 132418 190170 132486 190226
rect 132542 190170 132638 190226
rect 132018 190102 132638 190170
rect 132018 190046 132114 190102
rect 132170 190046 132238 190102
rect 132294 190046 132362 190102
rect 132418 190046 132486 190102
rect 132542 190046 132638 190102
rect 132018 189978 132638 190046
rect 132018 189922 132114 189978
rect 132170 189922 132238 189978
rect 132294 189922 132362 189978
rect 132418 189922 132486 189978
rect 132542 189922 132638 189978
rect 132018 172350 132638 189922
rect 132018 172294 132114 172350
rect 132170 172294 132238 172350
rect 132294 172294 132362 172350
rect 132418 172294 132486 172350
rect 132542 172294 132638 172350
rect 132018 172226 132638 172294
rect 132018 172170 132114 172226
rect 132170 172170 132238 172226
rect 132294 172170 132362 172226
rect 132418 172170 132486 172226
rect 132542 172170 132638 172226
rect 132018 172102 132638 172170
rect 132018 172046 132114 172102
rect 132170 172046 132238 172102
rect 132294 172046 132362 172102
rect 132418 172046 132486 172102
rect 132542 172046 132638 172102
rect 132018 171978 132638 172046
rect 132018 171922 132114 171978
rect 132170 171922 132238 171978
rect 132294 171922 132362 171978
rect 132418 171922 132486 171978
rect 132542 171922 132638 171978
rect 132018 154350 132638 171922
rect 135212 205380 135268 205390
rect 132018 154294 132114 154350
rect 132170 154294 132238 154350
rect 132294 154294 132362 154350
rect 132418 154294 132486 154350
rect 132542 154294 132638 154350
rect 132018 154226 132638 154294
rect 132018 154170 132114 154226
rect 132170 154170 132238 154226
rect 132294 154170 132362 154226
rect 132418 154170 132486 154226
rect 132542 154170 132638 154226
rect 132018 154102 132638 154170
rect 132018 154046 132114 154102
rect 132170 154046 132238 154102
rect 132294 154046 132362 154102
rect 132418 154046 132486 154102
rect 132542 154046 132638 154102
rect 132018 153978 132638 154046
rect 132018 153922 132114 153978
rect 132170 153922 132238 153978
rect 132294 153922 132362 153978
rect 132418 153922 132486 153978
rect 132542 153922 132638 153978
rect 132018 136350 132638 153922
rect 132018 136294 132114 136350
rect 132170 136294 132238 136350
rect 132294 136294 132362 136350
rect 132418 136294 132486 136350
rect 132542 136294 132638 136350
rect 132018 136226 132638 136294
rect 132018 136170 132114 136226
rect 132170 136170 132238 136226
rect 132294 136170 132362 136226
rect 132418 136170 132486 136226
rect 132542 136170 132638 136226
rect 132018 136102 132638 136170
rect 132018 136046 132114 136102
rect 132170 136046 132238 136102
rect 132294 136046 132362 136102
rect 132418 136046 132486 136102
rect 132542 136046 132638 136102
rect 132018 135978 132638 136046
rect 132018 135922 132114 135978
rect 132170 135922 132238 135978
rect 132294 135922 132362 135978
rect 132418 135922 132486 135978
rect 132542 135922 132638 135978
rect 128298 112294 128394 112350
rect 128450 112294 128518 112350
rect 128574 112294 128642 112350
rect 128698 112294 128766 112350
rect 128822 112294 128918 112350
rect 128298 112226 128918 112294
rect 128298 112170 128394 112226
rect 128450 112170 128518 112226
rect 128574 112170 128642 112226
rect 128698 112170 128766 112226
rect 128822 112170 128918 112226
rect 128298 112102 128918 112170
rect 128298 112046 128394 112102
rect 128450 112046 128518 112102
rect 128574 112046 128642 112102
rect 128698 112046 128766 112102
rect 128822 112046 128918 112102
rect 128298 111978 128918 112046
rect 128298 111922 128394 111978
rect 128450 111922 128518 111978
rect 128574 111922 128642 111978
rect 128698 111922 128766 111978
rect 128822 111922 128918 111978
rect 128298 94350 128918 111922
rect 128298 94294 128394 94350
rect 128450 94294 128518 94350
rect 128574 94294 128642 94350
rect 128698 94294 128766 94350
rect 128822 94294 128918 94350
rect 128298 94226 128918 94294
rect 128298 94170 128394 94226
rect 128450 94170 128518 94226
rect 128574 94170 128642 94226
rect 128698 94170 128766 94226
rect 128822 94170 128918 94226
rect 128298 94102 128918 94170
rect 128298 94046 128394 94102
rect 128450 94046 128518 94102
rect 128574 94046 128642 94102
rect 128698 94046 128766 94102
rect 128822 94046 128918 94102
rect 128298 93978 128918 94046
rect 128298 93922 128394 93978
rect 128450 93922 128518 93978
rect 128574 93922 128642 93978
rect 128698 93922 128766 93978
rect 128822 93922 128918 93978
rect 128298 76350 128918 93922
rect 128298 76294 128394 76350
rect 128450 76294 128518 76350
rect 128574 76294 128642 76350
rect 128698 76294 128766 76350
rect 128822 76294 128918 76350
rect 128298 76226 128918 76294
rect 128298 76170 128394 76226
rect 128450 76170 128518 76226
rect 128574 76170 128642 76226
rect 128698 76170 128766 76226
rect 128822 76170 128918 76226
rect 128298 76102 128918 76170
rect 128298 76046 128394 76102
rect 128450 76046 128518 76102
rect 128574 76046 128642 76102
rect 128698 76046 128766 76102
rect 128822 76046 128918 76102
rect 128298 75978 128918 76046
rect 128298 75922 128394 75978
rect 128450 75922 128518 75978
rect 128574 75922 128642 75978
rect 128698 75922 128766 75978
rect 128822 75922 128918 75978
rect 128298 58350 128918 75922
rect 128298 58294 128394 58350
rect 128450 58294 128518 58350
rect 128574 58294 128642 58350
rect 128698 58294 128766 58350
rect 128822 58294 128918 58350
rect 128298 58226 128918 58294
rect 128298 58170 128394 58226
rect 128450 58170 128518 58226
rect 128574 58170 128642 58226
rect 128698 58170 128766 58226
rect 128822 58170 128918 58226
rect 128298 58102 128918 58170
rect 128298 58046 128394 58102
rect 128450 58046 128518 58102
rect 128574 58046 128642 58102
rect 128698 58046 128766 58102
rect 128822 58046 128918 58102
rect 128298 57978 128918 58046
rect 128298 57922 128394 57978
rect 128450 57922 128518 57978
rect 128574 57922 128642 57978
rect 128698 57922 128766 57978
rect 128822 57922 128918 57978
rect 127596 47908 127652 47918
rect 127596 46340 127652 47852
rect 127596 46274 127652 46284
rect 127260 34626 127316 34636
rect 128298 40350 128918 57922
rect 128298 40294 128394 40350
rect 128450 40294 128518 40350
rect 128574 40294 128642 40350
rect 128698 40294 128766 40350
rect 128822 40294 128918 40350
rect 128298 40226 128918 40294
rect 128298 40170 128394 40226
rect 128450 40170 128518 40226
rect 128574 40170 128642 40226
rect 128698 40170 128766 40226
rect 128822 40170 128918 40226
rect 128298 40102 128918 40170
rect 128298 40046 128394 40102
rect 128450 40046 128518 40102
rect 128574 40046 128642 40102
rect 128698 40046 128766 40102
rect 128822 40046 128918 40102
rect 128298 39978 128918 40046
rect 128298 39922 128394 39978
rect 128450 39922 128518 39978
rect 128574 39922 128642 39978
rect 128698 39922 128766 39978
rect 128822 39922 128918 39978
rect 127036 33684 127092 33694
rect 126812 17154 126868 17164
rect 126924 30436 126980 30446
rect 126924 5572 126980 30380
rect 127036 11396 127092 33628
rect 127372 32788 127428 32798
rect 127036 11330 127092 11340
rect 127148 32004 127204 32014
rect 127148 8484 127204 31948
rect 127260 31108 127316 31118
rect 127260 14308 127316 31052
rect 127372 23044 127428 32732
rect 127372 22978 127428 22988
rect 127484 30324 127540 30334
rect 127484 20132 127540 30268
rect 127484 20066 127540 20076
rect 128298 22350 128918 39922
rect 129052 126084 129108 126094
rect 129052 31780 129108 126028
rect 132018 118350 132638 135922
rect 132018 118294 132114 118350
rect 132170 118294 132238 118350
rect 132294 118294 132362 118350
rect 132418 118294 132486 118350
rect 132542 118294 132638 118350
rect 132018 118226 132638 118294
rect 132018 118170 132114 118226
rect 132170 118170 132238 118226
rect 132294 118170 132362 118226
rect 132418 118170 132486 118226
rect 132542 118170 132638 118226
rect 132018 118102 132638 118170
rect 132018 118046 132114 118102
rect 132170 118046 132238 118102
rect 132294 118046 132362 118102
rect 132418 118046 132486 118102
rect 132542 118046 132638 118102
rect 132018 117978 132638 118046
rect 132018 117922 132114 117978
rect 132170 117922 132238 117978
rect 132294 117922 132362 117978
rect 132418 117922 132486 117978
rect 132542 117922 132638 117978
rect 132018 100350 132638 117922
rect 132018 100294 132114 100350
rect 132170 100294 132238 100350
rect 132294 100294 132362 100350
rect 132418 100294 132486 100350
rect 132542 100294 132638 100350
rect 132018 100226 132638 100294
rect 132018 100170 132114 100226
rect 132170 100170 132238 100226
rect 132294 100170 132362 100226
rect 132418 100170 132486 100226
rect 132542 100170 132638 100226
rect 132018 100102 132638 100170
rect 132018 100046 132114 100102
rect 132170 100046 132238 100102
rect 132294 100046 132362 100102
rect 132418 100046 132486 100102
rect 132542 100046 132638 100102
rect 132018 99978 132638 100046
rect 132018 99922 132114 99978
rect 132170 99922 132238 99978
rect 132294 99922 132362 99978
rect 132418 99922 132486 99978
rect 132542 99922 132638 99978
rect 132018 82350 132638 99922
rect 132018 82294 132114 82350
rect 132170 82294 132238 82350
rect 132294 82294 132362 82350
rect 132418 82294 132486 82350
rect 132542 82294 132638 82350
rect 132018 82226 132638 82294
rect 132018 82170 132114 82226
rect 132170 82170 132238 82226
rect 132294 82170 132362 82226
rect 132418 82170 132486 82226
rect 132542 82170 132638 82226
rect 132018 82102 132638 82170
rect 132018 82046 132114 82102
rect 132170 82046 132238 82102
rect 132294 82046 132362 82102
rect 132418 82046 132486 82102
rect 132542 82046 132638 82102
rect 132018 81978 132638 82046
rect 132018 81922 132114 81978
rect 132170 81922 132238 81978
rect 132294 81922 132362 81978
rect 132418 81922 132486 81978
rect 132542 81922 132638 81978
rect 129052 31714 129108 31724
rect 130172 73220 130228 73230
rect 130172 30324 130228 73164
rect 130172 30258 130228 30268
rect 132018 64350 132638 81922
rect 132018 64294 132114 64350
rect 132170 64294 132238 64350
rect 132294 64294 132362 64350
rect 132418 64294 132486 64350
rect 132542 64294 132638 64350
rect 132018 64226 132638 64294
rect 132018 64170 132114 64226
rect 132170 64170 132238 64226
rect 132294 64170 132362 64226
rect 132418 64170 132486 64226
rect 132542 64170 132638 64226
rect 132018 64102 132638 64170
rect 132018 64046 132114 64102
rect 132170 64046 132238 64102
rect 132294 64046 132362 64102
rect 132418 64046 132486 64102
rect 132542 64046 132638 64102
rect 132018 63978 132638 64046
rect 132018 63922 132114 63978
rect 132170 63922 132238 63978
rect 132294 63922 132362 63978
rect 132418 63922 132486 63978
rect 132542 63922 132638 63978
rect 132018 46350 132638 63922
rect 132018 46294 132114 46350
rect 132170 46294 132238 46350
rect 132294 46294 132362 46350
rect 132418 46294 132486 46350
rect 132542 46294 132638 46350
rect 132018 46226 132638 46294
rect 132018 46170 132114 46226
rect 132170 46170 132238 46226
rect 132294 46170 132362 46226
rect 132418 46170 132486 46226
rect 132542 46170 132638 46226
rect 132018 46102 132638 46170
rect 132018 46046 132114 46102
rect 132170 46046 132238 46102
rect 132294 46046 132362 46102
rect 132418 46046 132486 46102
rect 132542 46046 132638 46102
rect 132018 45978 132638 46046
rect 132018 45922 132114 45978
rect 132170 45922 132238 45978
rect 132294 45922 132362 45978
rect 132418 45922 132486 45978
rect 132542 45922 132638 45978
rect 132018 28350 132638 45922
rect 133532 163828 133588 163838
rect 132018 28294 132114 28350
rect 132170 28294 132238 28350
rect 132294 28294 132362 28350
rect 132418 28294 132486 28350
rect 132542 28294 132638 28350
rect 132018 28226 132638 28294
rect 132018 28170 132114 28226
rect 132170 28170 132238 28226
rect 132294 28170 132362 28226
rect 132418 28170 132486 28226
rect 132542 28170 132638 28226
rect 132018 28102 132638 28170
rect 132018 28046 132114 28102
rect 132170 28046 132238 28102
rect 132294 28046 132362 28102
rect 132418 28046 132486 28102
rect 132542 28046 132638 28102
rect 132018 27978 132638 28046
rect 132018 27922 132114 27978
rect 132170 27922 132238 27978
rect 132294 27922 132362 27978
rect 132418 27922 132486 27978
rect 132542 27922 132638 27978
rect 128298 22294 128394 22350
rect 128450 22294 128518 22350
rect 128574 22294 128642 22350
rect 128698 22294 128766 22350
rect 128822 22294 128918 22350
rect 128298 22226 128918 22294
rect 128298 22170 128394 22226
rect 128450 22170 128518 22226
rect 128574 22170 128642 22226
rect 128698 22170 128766 22226
rect 128822 22170 128918 22226
rect 128298 22102 128918 22170
rect 128298 22046 128394 22102
rect 128450 22046 128518 22102
rect 128574 22046 128642 22102
rect 128698 22046 128766 22102
rect 128822 22046 128918 22102
rect 128298 21978 128918 22046
rect 128298 21922 128394 21978
rect 128450 21922 128518 21978
rect 128574 21922 128642 21978
rect 128698 21922 128766 21978
rect 128822 21922 128918 21978
rect 127260 14242 127316 14252
rect 127148 8418 127204 8428
rect 126924 5506 126980 5516
rect 126028 4162 126084 4172
rect 128298 4350 128918 21922
rect 128298 4294 128394 4350
rect 128450 4294 128518 4350
rect 128574 4294 128642 4350
rect 128698 4294 128766 4350
rect 128822 4294 128918 4350
rect 128298 4226 128918 4294
rect 128298 4170 128394 4226
rect 128450 4170 128518 4226
rect 128574 4170 128642 4226
rect 128698 4170 128766 4226
rect 128822 4170 128918 4226
rect 123452 3266 123508 3276
rect 128298 4102 128918 4170
rect 128298 4046 128394 4102
rect 128450 4046 128518 4102
rect 128574 4046 128642 4102
rect 128698 4046 128766 4102
rect 128822 4046 128918 4102
rect 128298 3978 128918 4046
rect 128298 3922 128394 3978
rect 128450 3922 128518 3978
rect 128574 3922 128642 3978
rect 128698 3922 128766 3978
rect 128822 3922 128918 3978
rect 121772 2482 121828 2492
rect 117964 2458 118020 2468
rect 117964 2100 118020 2402
rect 117964 2034 118020 2044
rect 101298 -1176 101394 -1120
rect 101450 -1176 101518 -1120
rect 101574 -1176 101642 -1120
rect 101698 -1176 101766 -1120
rect 101822 -1176 101918 -1120
rect 101298 -1244 101918 -1176
rect 101298 -1300 101394 -1244
rect 101450 -1300 101518 -1244
rect 101574 -1300 101642 -1244
rect 101698 -1300 101766 -1244
rect 101822 -1300 101918 -1244
rect 101298 -1368 101918 -1300
rect 101298 -1424 101394 -1368
rect 101450 -1424 101518 -1368
rect 101574 -1424 101642 -1368
rect 101698 -1424 101766 -1368
rect 101822 -1424 101918 -1368
rect 101298 -1492 101918 -1424
rect 101298 -1548 101394 -1492
rect 101450 -1548 101518 -1492
rect 101574 -1548 101642 -1492
rect 101698 -1548 101766 -1492
rect 101822 -1548 101918 -1492
rect 101298 -1644 101918 -1548
rect 128298 -160 128918 3922
rect 130172 23604 130228 23614
rect 130172 1198 130228 23548
rect 131292 14338 131348 14348
rect 131292 4228 131348 14282
rect 131292 4162 131348 4172
rect 132018 10350 132638 27922
rect 132018 10294 132114 10350
rect 132170 10294 132238 10350
rect 132294 10294 132362 10350
rect 132418 10294 132486 10350
rect 132542 10294 132638 10350
rect 132018 10226 132638 10294
rect 132018 10170 132114 10226
rect 132170 10170 132238 10226
rect 132294 10170 132362 10226
rect 132418 10170 132486 10226
rect 132542 10170 132638 10226
rect 132018 10102 132638 10170
rect 132018 10046 132114 10102
rect 132170 10046 132238 10102
rect 132294 10046 132362 10102
rect 132418 10046 132486 10102
rect 132542 10046 132638 10102
rect 132018 9978 132638 10046
rect 132018 9922 132114 9978
rect 132170 9922 132238 9978
rect 132294 9922 132362 9978
rect 132418 9922 132486 9978
rect 132542 9922 132638 9978
rect 130172 1132 130228 1142
rect 128298 -216 128394 -160
rect 128450 -216 128518 -160
rect 128574 -216 128642 -160
rect 128698 -216 128766 -160
rect 128822 -216 128918 -160
rect 128298 -284 128918 -216
rect 128298 -340 128394 -284
rect 128450 -340 128518 -284
rect 128574 -340 128642 -284
rect 128698 -340 128766 -284
rect 128822 -340 128918 -284
rect 128298 -408 128918 -340
rect 128298 -464 128394 -408
rect 128450 -464 128518 -408
rect 128574 -464 128642 -408
rect 128698 -464 128766 -408
rect 128822 -464 128918 -408
rect 128298 -532 128918 -464
rect 128298 -588 128394 -532
rect 128450 -588 128518 -532
rect 128574 -588 128642 -532
rect 128698 -588 128766 -532
rect 128822 -588 128918 -532
rect 128298 -1644 128918 -588
rect 132018 -1120 132638 9922
rect 132748 44578 132804 44588
rect 132748 4228 132804 44522
rect 133532 40516 133588 163772
rect 133532 40450 133588 40460
rect 134428 51238 134484 51248
rect 132748 4162 132804 4172
rect 134428 4228 134484 51182
rect 135212 49252 135268 205324
rect 136892 57988 136948 242732
rect 141932 192164 141988 192174
rect 140252 152516 140308 152526
rect 136892 57922 136948 57932
rect 138572 112868 138628 112878
rect 135212 49186 135268 49196
rect 138572 28868 138628 112812
rect 140252 37604 140308 152460
rect 141932 47908 141988 192108
rect 145292 63812 145348 271404
rect 145292 63746 145348 63756
rect 148652 231924 148708 231934
rect 148652 55076 148708 231868
rect 150332 69636 150388 296492
rect 150332 69570 150388 69580
rect 159018 292350 159638 309922
rect 159018 292294 159114 292350
rect 159170 292294 159238 292350
rect 159294 292294 159362 292350
rect 159418 292294 159486 292350
rect 159542 292294 159638 292350
rect 159018 292226 159638 292294
rect 159018 292170 159114 292226
rect 159170 292170 159238 292226
rect 159294 292170 159362 292226
rect 159418 292170 159486 292226
rect 159542 292170 159638 292226
rect 159018 292102 159638 292170
rect 159018 292046 159114 292102
rect 159170 292046 159238 292102
rect 159294 292046 159362 292102
rect 159418 292046 159486 292102
rect 159542 292046 159638 292102
rect 159018 291978 159638 292046
rect 159018 291922 159114 291978
rect 159170 291922 159238 291978
rect 159294 291922 159362 291978
rect 159418 291922 159486 291978
rect 159542 291922 159638 291978
rect 159018 274350 159638 291922
rect 159018 274294 159114 274350
rect 159170 274294 159238 274350
rect 159294 274294 159362 274350
rect 159418 274294 159486 274350
rect 159542 274294 159638 274350
rect 159018 274226 159638 274294
rect 159018 274170 159114 274226
rect 159170 274170 159238 274226
rect 159294 274170 159362 274226
rect 159418 274170 159486 274226
rect 159542 274170 159638 274226
rect 159018 274102 159638 274170
rect 159018 274046 159114 274102
rect 159170 274046 159238 274102
rect 159294 274046 159362 274102
rect 159418 274046 159486 274102
rect 159542 274046 159638 274102
rect 159018 273978 159638 274046
rect 159018 273922 159114 273978
rect 159170 273922 159238 273978
rect 159294 273922 159362 273978
rect 159418 273922 159486 273978
rect 159542 273922 159638 273978
rect 159018 256350 159638 273922
rect 159018 256294 159114 256350
rect 159170 256294 159238 256350
rect 159294 256294 159362 256350
rect 159418 256294 159486 256350
rect 159542 256294 159638 256350
rect 159018 256226 159638 256294
rect 159018 256170 159114 256226
rect 159170 256170 159238 256226
rect 159294 256170 159362 256226
rect 159418 256170 159486 256226
rect 159542 256170 159638 256226
rect 159018 256102 159638 256170
rect 159018 256046 159114 256102
rect 159170 256046 159238 256102
rect 159294 256046 159362 256102
rect 159418 256046 159486 256102
rect 159542 256046 159638 256102
rect 159018 255978 159638 256046
rect 159018 255922 159114 255978
rect 159170 255922 159238 255978
rect 159294 255922 159362 255978
rect 159418 255922 159486 255978
rect 159542 255922 159638 255978
rect 159018 238350 159638 255922
rect 159018 238294 159114 238350
rect 159170 238294 159238 238350
rect 159294 238294 159362 238350
rect 159418 238294 159486 238350
rect 159542 238294 159638 238350
rect 159018 238226 159638 238294
rect 159018 238170 159114 238226
rect 159170 238170 159238 238226
rect 159294 238170 159362 238226
rect 159418 238170 159486 238226
rect 159542 238170 159638 238226
rect 159018 238102 159638 238170
rect 159018 238046 159114 238102
rect 159170 238046 159238 238102
rect 159294 238046 159362 238102
rect 159418 238046 159486 238102
rect 159542 238046 159638 238102
rect 159018 237978 159638 238046
rect 159018 237922 159114 237978
rect 159170 237922 159238 237978
rect 159294 237922 159362 237978
rect 159418 237922 159486 237978
rect 159542 237922 159638 237978
rect 159018 220350 159638 237922
rect 159018 220294 159114 220350
rect 159170 220294 159238 220350
rect 159294 220294 159362 220350
rect 159418 220294 159486 220350
rect 159542 220294 159638 220350
rect 159018 220226 159638 220294
rect 159018 220170 159114 220226
rect 159170 220170 159238 220226
rect 159294 220170 159362 220226
rect 159418 220170 159486 220226
rect 159542 220170 159638 220226
rect 159018 220102 159638 220170
rect 159018 220046 159114 220102
rect 159170 220046 159238 220102
rect 159294 220046 159362 220102
rect 159418 220046 159486 220102
rect 159542 220046 159638 220102
rect 159018 219978 159638 220046
rect 159018 219922 159114 219978
rect 159170 219922 159238 219978
rect 159294 219922 159362 219978
rect 159418 219922 159486 219978
rect 159542 219922 159638 219978
rect 159018 202350 159638 219922
rect 159018 202294 159114 202350
rect 159170 202294 159238 202350
rect 159294 202294 159362 202350
rect 159418 202294 159486 202350
rect 159542 202294 159638 202350
rect 159018 202226 159638 202294
rect 159018 202170 159114 202226
rect 159170 202170 159238 202226
rect 159294 202170 159362 202226
rect 159418 202170 159486 202226
rect 159542 202170 159638 202226
rect 159018 202102 159638 202170
rect 159018 202046 159114 202102
rect 159170 202046 159238 202102
rect 159294 202046 159362 202102
rect 159418 202046 159486 202102
rect 159542 202046 159638 202102
rect 159018 201978 159638 202046
rect 159018 201922 159114 201978
rect 159170 201922 159238 201978
rect 159294 201922 159362 201978
rect 159418 201922 159486 201978
rect 159542 201922 159638 201978
rect 159018 184350 159638 201922
rect 159018 184294 159114 184350
rect 159170 184294 159238 184350
rect 159294 184294 159362 184350
rect 159418 184294 159486 184350
rect 159542 184294 159638 184350
rect 159018 184226 159638 184294
rect 159018 184170 159114 184226
rect 159170 184170 159238 184226
rect 159294 184170 159362 184226
rect 159418 184170 159486 184226
rect 159542 184170 159638 184226
rect 159018 184102 159638 184170
rect 159018 184046 159114 184102
rect 159170 184046 159238 184102
rect 159294 184046 159362 184102
rect 159418 184046 159486 184102
rect 159542 184046 159638 184102
rect 159018 183978 159638 184046
rect 159018 183922 159114 183978
rect 159170 183922 159238 183978
rect 159294 183922 159362 183978
rect 159418 183922 159486 183978
rect 159542 183922 159638 183978
rect 159018 166350 159638 183922
rect 159018 166294 159114 166350
rect 159170 166294 159238 166350
rect 159294 166294 159362 166350
rect 159418 166294 159486 166350
rect 159542 166294 159638 166350
rect 159018 166226 159638 166294
rect 159018 166170 159114 166226
rect 159170 166170 159238 166226
rect 159294 166170 159362 166226
rect 159418 166170 159486 166226
rect 159542 166170 159638 166226
rect 159018 166102 159638 166170
rect 159018 166046 159114 166102
rect 159170 166046 159238 166102
rect 159294 166046 159362 166102
rect 159418 166046 159486 166102
rect 159542 166046 159638 166102
rect 159018 165978 159638 166046
rect 159018 165922 159114 165978
rect 159170 165922 159238 165978
rect 159294 165922 159362 165978
rect 159418 165922 159486 165978
rect 159542 165922 159638 165978
rect 159018 148350 159638 165922
rect 159018 148294 159114 148350
rect 159170 148294 159238 148350
rect 159294 148294 159362 148350
rect 159418 148294 159486 148350
rect 159542 148294 159638 148350
rect 159018 148226 159638 148294
rect 159018 148170 159114 148226
rect 159170 148170 159238 148226
rect 159294 148170 159362 148226
rect 159418 148170 159486 148226
rect 159542 148170 159638 148226
rect 159018 148102 159638 148170
rect 159018 148046 159114 148102
rect 159170 148046 159238 148102
rect 159294 148046 159362 148102
rect 159418 148046 159486 148102
rect 159542 148046 159638 148102
rect 159018 147978 159638 148046
rect 159018 147922 159114 147978
rect 159170 147922 159238 147978
rect 159294 147922 159362 147978
rect 159418 147922 159486 147978
rect 159542 147922 159638 147978
rect 159018 130350 159638 147922
rect 159018 130294 159114 130350
rect 159170 130294 159238 130350
rect 159294 130294 159362 130350
rect 159418 130294 159486 130350
rect 159542 130294 159638 130350
rect 159018 130226 159638 130294
rect 159018 130170 159114 130226
rect 159170 130170 159238 130226
rect 159294 130170 159362 130226
rect 159418 130170 159486 130226
rect 159542 130170 159638 130226
rect 159018 130102 159638 130170
rect 159018 130046 159114 130102
rect 159170 130046 159238 130102
rect 159294 130046 159362 130102
rect 159418 130046 159486 130102
rect 159542 130046 159638 130102
rect 159018 129978 159638 130046
rect 159018 129922 159114 129978
rect 159170 129922 159238 129978
rect 159294 129922 159362 129978
rect 159418 129922 159486 129978
rect 159542 129922 159638 129978
rect 159018 112350 159638 129922
rect 159018 112294 159114 112350
rect 159170 112294 159238 112350
rect 159294 112294 159362 112350
rect 159418 112294 159486 112350
rect 159542 112294 159638 112350
rect 159018 112226 159638 112294
rect 159018 112170 159114 112226
rect 159170 112170 159238 112226
rect 159294 112170 159362 112226
rect 159418 112170 159486 112226
rect 159542 112170 159638 112226
rect 159018 112102 159638 112170
rect 159018 112046 159114 112102
rect 159170 112046 159238 112102
rect 159294 112046 159362 112102
rect 159418 112046 159486 112102
rect 159542 112046 159638 112102
rect 159018 111978 159638 112046
rect 159018 111922 159114 111978
rect 159170 111922 159238 111978
rect 159294 111922 159362 111978
rect 159418 111922 159486 111978
rect 159542 111922 159638 111978
rect 159018 94350 159638 111922
rect 159018 94294 159114 94350
rect 159170 94294 159238 94350
rect 159294 94294 159362 94350
rect 159418 94294 159486 94350
rect 159542 94294 159638 94350
rect 159018 94226 159638 94294
rect 159018 94170 159114 94226
rect 159170 94170 159238 94226
rect 159294 94170 159362 94226
rect 159418 94170 159486 94226
rect 159542 94170 159638 94226
rect 159018 94102 159638 94170
rect 159018 94046 159114 94102
rect 159170 94046 159238 94102
rect 159294 94046 159362 94102
rect 159418 94046 159486 94102
rect 159542 94046 159638 94102
rect 159018 93978 159638 94046
rect 159018 93922 159114 93978
rect 159170 93922 159238 93978
rect 159294 93922 159362 93978
rect 159418 93922 159486 93978
rect 159542 93922 159638 93978
rect 159018 76350 159638 93922
rect 159018 76294 159114 76350
rect 159170 76294 159238 76350
rect 159294 76294 159362 76350
rect 159418 76294 159486 76350
rect 159542 76294 159638 76350
rect 159018 76226 159638 76294
rect 159018 76170 159114 76226
rect 159170 76170 159238 76226
rect 159294 76170 159362 76226
rect 159418 76170 159486 76226
rect 159542 76170 159638 76226
rect 159018 76102 159638 76170
rect 159018 76046 159114 76102
rect 159170 76046 159238 76102
rect 159294 76046 159362 76102
rect 159418 76046 159486 76102
rect 159542 76046 159638 76102
rect 159018 75978 159638 76046
rect 159018 75922 159114 75978
rect 159170 75922 159238 75978
rect 159294 75922 159362 75978
rect 159418 75922 159486 75978
rect 159542 75922 159638 75978
rect 148652 55010 148708 55020
rect 159018 58350 159638 75922
rect 159018 58294 159114 58350
rect 159170 58294 159238 58350
rect 159294 58294 159362 58350
rect 159418 58294 159486 58350
rect 159542 58294 159638 58350
rect 159018 58226 159638 58294
rect 159018 58170 159114 58226
rect 159170 58170 159238 58226
rect 159294 58170 159362 58226
rect 159418 58170 159486 58226
rect 159542 58170 159638 58226
rect 159018 58102 159638 58170
rect 159018 58046 159114 58102
rect 159170 58046 159238 58102
rect 159294 58046 159362 58102
rect 159418 58046 159486 58102
rect 159542 58046 159638 58102
rect 159018 57978 159638 58046
rect 159018 57922 159114 57978
rect 159170 57922 159238 57978
rect 159294 57922 159362 57978
rect 159418 57922 159486 57978
rect 159542 57922 159638 57978
rect 141932 47842 141988 47852
rect 140252 37538 140308 37548
rect 147868 41158 147924 41168
rect 138572 28802 138628 28812
rect 142828 29278 142884 29288
rect 134428 4162 134484 4172
rect 137788 19198 137844 19208
rect 137788 4228 137844 19142
rect 137788 4162 137844 4172
rect 139468 12538 139524 12548
rect 139468 4228 139524 12482
rect 139468 4162 139524 4172
rect 142828 4228 142884 29222
rect 144508 24418 144564 24428
rect 144508 20188 144564 24362
rect 144508 20132 144676 20188
rect 142828 4162 142884 4172
rect 144620 4228 144676 20132
rect 144620 4162 144676 4172
rect 146188 15958 146244 15968
rect 146188 4228 146244 15902
rect 146188 4162 146244 4172
rect 147868 4228 147924 41102
rect 159018 40350 159638 57922
rect 159018 40294 159114 40350
rect 159170 40294 159238 40350
rect 159294 40294 159362 40350
rect 159418 40294 159486 40350
rect 159542 40294 159638 40350
rect 159018 40226 159638 40294
rect 159018 40170 159114 40226
rect 159170 40170 159238 40226
rect 159294 40170 159362 40226
rect 159418 40170 159486 40226
rect 159542 40170 159638 40226
rect 159018 40102 159638 40170
rect 159018 40046 159114 40102
rect 159170 40046 159238 40102
rect 159294 40046 159362 40102
rect 159418 40046 159486 40102
rect 159542 40046 159638 40102
rect 159018 39978 159638 40046
rect 159018 39922 159114 39978
rect 159170 39922 159238 39978
rect 159294 39922 159362 39978
rect 159418 39922 159486 39978
rect 159542 39922 159638 39978
rect 151228 37738 151284 37748
rect 147868 4162 147924 4172
rect 149548 17578 149604 17588
rect 149548 4228 149604 17522
rect 149548 4162 149604 4172
rect 151228 4228 151284 37682
rect 154588 30898 154644 30908
rect 151228 4162 151284 4172
rect 152908 24238 152964 24248
rect 152908 4228 152964 24182
rect 152908 4162 152964 4172
rect 154588 4228 154644 30842
rect 159018 22350 159638 39922
rect 159018 22294 159114 22350
rect 159170 22294 159238 22350
rect 159294 22294 159362 22350
rect 159418 22294 159486 22350
rect 159542 22294 159638 22350
rect 159018 22226 159638 22294
rect 159018 22170 159114 22226
rect 159170 22170 159238 22226
rect 159294 22170 159362 22226
rect 159418 22170 159486 22226
rect 159542 22170 159638 22226
rect 159018 22102 159638 22170
rect 159018 22046 159114 22102
rect 159170 22046 159238 22102
rect 159294 22046 159362 22102
rect 159418 22046 159486 22102
rect 159542 22046 159638 22102
rect 159018 21978 159638 22046
rect 159018 21922 159114 21978
rect 159170 21922 159238 21978
rect 159294 21922 159362 21978
rect 159418 21922 159486 21978
rect 159542 21922 159638 21978
rect 154588 4162 154644 4172
rect 157948 19018 158004 19028
rect 157948 4228 158004 18962
rect 157948 4162 158004 4172
rect 159018 4350 159638 21922
rect 162738 598172 163358 598268
rect 162738 598116 162834 598172
rect 162890 598116 162958 598172
rect 163014 598116 163082 598172
rect 163138 598116 163206 598172
rect 163262 598116 163358 598172
rect 162738 598048 163358 598116
rect 162738 597992 162834 598048
rect 162890 597992 162958 598048
rect 163014 597992 163082 598048
rect 163138 597992 163206 598048
rect 163262 597992 163358 598048
rect 162738 597924 163358 597992
rect 162738 597868 162834 597924
rect 162890 597868 162958 597924
rect 163014 597868 163082 597924
rect 163138 597868 163206 597924
rect 163262 597868 163358 597924
rect 162738 597800 163358 597868
rect 162738 597744 162834 597800
rect 162890 597744 162958 597800
rect 163014 597744 163082 597800
rect 163138 597744 163206 597800
rect 163262 597744 163358 597800
rect 162738 586350 163358 597744
rect 189738 597212 190358 598268
rect 189738 597156 189834 597212
rect 189890 597156 189958 597212
rect 190014 597156 190082 597212
rect 190138 597156 190206 597212
rect 190262 597156 190358 597212
rect 189738 597088 190358 597156
rect 189738 597032 189834 597088
rect 189890 597032 189958 597088
rect 190014 597032 190082 597088
rect 190138 597032 190206 597088
rect 190262 597032 190358 597088
rect 189738 596964 190358 597032
rect 189738 596908 189834 596964
rect 189890 596908 189958 596964
rect 190014 596908 190082 596964
rect 190138 596908 190206 596964
rect 190262 596908 190358 596964
rect 189738 596840 190358 596908
rect 189738 596784 189834 596840
rect 189890 596784 189958 596840
rect 190014 596784 190082 596840
rect 190138 596784 190206 596840
rect 190262 596784 190358 596840
rect 162738 586294 162834 586350
rect 162890 586294 162958 586350
rect 163014 586294 163082 586350
rect 163138 586294 163206 586350
rect 163262 586294 163358 586350
rect 162738 586226 163358 586294
rect 162738 586170 162834 586226
rect 162890 586170 162958 586226
rect 163014 586170 163082 586226
rect 163138 586170 163206 586226
rect 163262 586170 163358 586226
rect 162738 586102 163358 586170
rect 162738 586046 162834 586102
rect 162890 586046 162958 586102
rect 163014 586046 163082 586102
rect 163138 586046 163206 586102
rect 163262 586046 163358 586102
rect 162738 585978 163358 586046
rect 162738 585922 162834 585978
rect 162890 585922 162958 585978
rect 163014 585922 163082 585978
rect 163138 585922 163206 585978
rect 163262 585922 163358 585978
rect 162738 568350 163358 585922
rect 162738 568294 162834 568350
rect 162890 568294 162958 568350
rect 163014 568294 163082 568350
rect 163138 568294 163206 568350
rect 163262 568294 163358 568350
rect 162738 568226 163358 568294
rect 162738 568170 162834 568226
rect 162890 568170 162958 568226
rect 163014 568170 163082 568226
rect 163138 568170 163206 568226
rect 163262 568170 163358 568226
rect 162738 568102 163358 568170
rect 162738 568046 162834 568102
rect 162890 568046 162958 568102
rect 163014 568046 163082 568102
rect 163138 568046 163206 568102
rect 163262 568046 163358 568102
rect 162738 567978 163358 568046
rect 162738 567922 162834 567978
rect 162890 567922 162958 567978
rect 163014 567922 163082 567978
rect 163138 567922 163206 567978
rect 163262 567922 163358 567978
rect 162738 550350 163358 567922
rect 162738 550294 162834 550350
rect 162890 550294 162958 550350
rect 163014 550294 163082 550350
rect 163138 550294 163206 550350
rect 163262 550294 163358 550350
rect 162738 550226 163358 550294
rect 162738 550170 162834 550226
rect 162890 550170 162958 550226
rect 163014 550170 163082 550226
rect 163138 550170 163206 550226
rect 163262 550170 163358 550226
rect 162738 550102 163358 550170
rect 162738 550046 162834 550102
rect 162890 550046 162958 550102
rect 163014 550046 163082 550102
rect 163138 550046 163206 550102
rect 163262 550046 163358 550102
rect 162738 549978 163358 550046
rect 162738 549922 162834 549978
rect 162890 549922 162958 549978
rect 163014 549922 163082 549978
rect 163138 549922 163206 549978
rect 163262 549922 163358 549978
rect 162738 532350 163358 549922
rect 162738 532294 162834 532350
rect 162890 532294 162958 532350
rect 163014 532294 163082 532350
rect 163138 532294 163206 532350
rect 163262 532294 163358 532350
rect 162738 532226 163358 532294
rect 162738 532170 162834 532226
rect 162890 532170 162958 532226
rect 163014 532170 163082 532226
rect 163138 532170 163206 532226
rect 163262 532170 163358 532226
rect 162738 532102 163358 532170
rect 162738 532046 162834 532102
rect 162890 532046 162958 532102
rect 163014 532046 163082 532102
rect 163138 532046 163206 532102
rect 163262 532046 163358 532102
rect 162738 531978 163358 532046
rect 162738 531922 162834 531978
rect 162890 531922 162958 531978
rect 163014 531922 163082 531978
rect 163138 531922 163206 531978
rect 163262 531922 163358 531978
rect 162738 514350 163358 531922
rect 162738 514294 162834 514350
rect 162890 514294 162958 514350
rect 163014 514294 163082 514350
rect 163138 514294 163206 514350
rect 163262 514294 163358 514350
rect 162738 514226 163358 514294
rect 162738 514170 162834 514226
rect 162890 514170 162958 514226
rect 163014 514170 163082 514226
rect 163138 514170 163206 514226
rect 163262 514170 163358 514226
rect 162738 514102 163358 514170
rect 162738 514046 162834 514102
rect 162890 514046 162958 514102
rect 163014 514046 163082 514102
rect 163138 514046 163206 514102
rect 163262 514046 163358 514102
rect 162738 513978 163358 514046
rect 162738 513922 162834 513978
rect 162890 513922 162958 513978
rect 163014 513922 163082 513978
rect 163138 513922 163206 513978
rect 163262 513922 163358 513978
rect 162738 496350 163358 513922
rect 162738 496294 162834 496350
rect 162890 496294 162958 496350
rect 163014 496294 163082 496350
rect 163138 496294 163206 496350
rect 163262 496294 163358 496350
rect 162738 496226 163358 496294
rect 162738 496170 162834 496226
rect 162890 496170 162958 496226
rect 163014 496170 163082 496226
rect 163138 496170 163206 496226
rect 163262 496170 163358 496226
rect 162738 496102 163358 496170
rect 162738 496046 162834 496102
rect 162890 496046 162958 496102
rect 163014 496046 163082 496102
rect 163138 496046 163206 496102
rect 163262 496046 163358 496102
rect 162738 495978 163358 496046
rect 162738 495922 162834 495978
rect 162890 495922 162958 495978
rect 163014 495922 163082 495978
rect 163138 495922 163206 495978
rect 163262 495922 163358 495978
rect 162738 478350 163358 495922
rect 162738 478294 162834 478350
rect 162890 478294 162958 478350
rect 163014 478294 163082 478350
rect 163138 478294 163206 478350
rect 163262 478294 163358 478350
rect 162738 478226 163358 478294
rect 162738 478170 162834 478226
rect 162890 478170 162958 478226
rect 163014 478170 163082 478226
rect 163138 478170 163206 478226
rect 163262 478170 163358 478226
rect 162738 478102 163358 478170
rect 162738 478046 162834 478102
rect 162890 478046 162958 478102
rect 163014 478046 163082 478102
rect 163138 478046 163206 478102
rect 163262 478046 163358 478102
rect 162738 477978 163358 478046
rect 162738 477922 162834 477978
rect 162890 477922 162958 477978
rect 163014 477922 163082 477978
rect 163138 477922 163206 477978
rect 163262 477922 163358 477978
rect 162738 460350 163358 477922
rect 162738 460294 162834 460350
rect 162890 460294 162958 460350
rect 163014 460294 163082 460350
rect 163138 460294 163206 460350
rect 163262 460294 163358 460350
rect 162738 460226 163358 460294
rect 162738 460170 162834 460226
rect 162890 460170 162958 460226
rect 163014 460170 163082 460226
rect 163138 460170 163206 460226
rect 163262 460170 163358 460226
rect 162738 460102 163358 460170
rect 162738 460046 162834 460102
rect 162890 460046 162958 460102
rect 163014 460046 163082 460102
rect 163138 460046 163206 460102
rect 163262 460046 163358 460102
rect 162738 459978 163358 460046
rect 162738 459922 162834 459978
rect 162890 459922 162958 459978
rect 163014 459922 163082 459978
rect 163138 459922 163206 459978
rect 163262 459922 163358 459978
rect 162738 442350 163358 459922
rect 162738 442294 162834 442350
rect 162890 442294 162958 442350
rect 163014 442294 163082 442350
rect 163138 442294 163206 442350
rect 163262 442294 163358 442350
rect 162738 442226 163358 442294
rect 162738 442170 162834 442226
rect 162890 442170 162958 442226
rect 163014 442170 163082 442226
rect 163138 442170 163206 442226
rect 163262 442170 163358 442226
rect 162738 442102 163358 442170
rect 162738 442046 162834 442102
rect 162890 442046 162958 442102
rect 163014 442046 163082 442102
rect 163138 442046 163206 442102
rect 163262 442046 163358 442102
rect 162738 441978 163358 442046
rect 162738 441922 162834 441978
rect 162890 441922 162958 441978
rect 163014 441922 163082 441978
rect 163138 441922 163206 441978
rect 163262 441922 163358 441978
rect 162738 424350 163358 441922
rect 162738 424294 162834 424350
rect 162890 424294 162958 424350
rect 163014 424294 163082 424350
rect 163138 424294 163206 424350
rect 163262 424294 163358 424350
rect 162738 424226 163358 424294
rect 162738 424170 162834 424226
rect 162890 424170 162958 424226
rect 163014 424170 163082 424226
rect 163138 424170 163206 424226
rect 163262 424170 163358 424226
rect 162738 424102 163358 424170
rect 162738 424046 162834 424102
rect 162890 424046 162958 424102
rect 163014 424046 163082 424102
rect 163138 424046 163206 424102
rect 163262 424046 163358 424102
rect 162738 423978 163358 424046
rect 162738 423922 162834 423978
rect 162890 423922 162958 423978
rect 163014 423922 163082 423978
rect 163138 423922 163206 423978
rect 163262 423922 163358 423978
rect 162738 406350 163358 423922
rect 162738 406294 162834 406350
rect 162890 406294 162958 406350
rect 163014 406294 163082 406350
rect 163138 406294 163206 406350
rect 163262 406294 163358 406350
rect 162738 406226 163358 406294
rect 162738 406170 162834 406226
rect 162890 406170 162958 406226
rect 163014 406170 163082 406226
rect 163138 406170 163206 406226
rect 163262 406170 163358 406226
rect 162738 406102 163358 406170
rect 162738 406046 162834 406102
rect 162890 406046 162958 406102
rect 163014 406046 163082 406102
rect 163138 406046 163206 406102
rect 163262 406046 163358 406102
rect 162738 405978 163358 406046
rect 162738 405922 162834 405978
rect 162890 405922 162958 405978
rect 163014 405922 163082 405978
rect 163138 405922 163206 405978
rect 163262 405922 163358 405978
rect 162738 388350 163358 405922
rect 162738 388294 162834 388350
rect 162890 388294 162958 388350
rect 163014 388294 163082 388350
rect 163138 388294 163206 388350
rect 163262 388294 163358 388350
rect 162738 388226 163358 388294
rect 162738 388170 162834 388226
rect 162890 388170 162958 388226
rect 163014 388170 163082 388226
rect 163138 388170 163206 388226
rect 163262 388170 163358 388226
rect 162738 388102 163358 388170
rect 162738 388046 162834 388102
rect 162890 388046 162958 388102
rect 163014 388046 163082 388102
rect 163138 388046 163206 388102
rect 163262 388046 163358 388102
rect 162738 387978 163358 388046
rect 162738 387922 162834 387978
rect 162890 387922 162958 387978
rect 163014 387922 163082 387978
rect 163138 387922 163206 387978
rect 163262 387922 163358 387978
rect 162738 370350 163358 387922
rect 162738 370294 162834 370350
rect 162890 370294 162958 370350
rect 163014 370294 163082 370350
rect 163138 370294 163206 370350
rect 163262 370294 163358 370350
rect 162738 370226 163358 370294
rect 162738 370170 162834 370226
rect 162890 370170 162958 370226
rect 163014 370170 163082 370226
rect 163138 370170 163206 370226
rect 163262 370170 163358 370226
rect 162738 370102 163358 370170
rect 162738 370046 162834 370102
rect 162890 370046 162958 370102
rect 163014 370046 163082 370102
rect 163138 370046 163206 370102
rect 163262 370046 163358 370102
rect 162738 369978 163358 370046
rect 162738 369922 162834 369978
rect 162890 369922 162958 369978
rect 163014 369922 163082 369978
rect 163138 369922 163206 369978
rect 163262 369922 163358 369978
rect 162738 352350 163358 369922
rect 162738 352294 162834 352350
rect 162890 352294 162958 352350
rect 163014 352294 163082 352350
rect 163138 352294 163206 352350
rect 163262 352294 163358 352350
rect 162738 352226 163358 352294
rect 162738 352170 162834 352226
rect 162890 352170 162958 352226
rect 163014 352170 163082 352226
rect 163138 352170 163206 352226
rect 163262 352170 163358 352226
rect 162738 352102 163358 352170
rect 162738 352046 162834 352102
rect 162890 352046 162958 352102
rect 163014 352046 163082 352102
rect 163138 352046 163206 352102
rect 163262 352046 163358 352102
rect 162738 351978 163358 352046
rect 162738 351922 162834 351978
rect 162890 351922 162958 351978
rect 163014 351922 163082 351978
rect 163138 351922 163206 351978
rect 163262 351922 163358 351978
rect 162738 334350 163358 351922
rect 162738 334294 162834 334350
rect 162890 334294 162958 334350
rect 163014 334294 163082 334350
rect 163138 334294 163206 334350
rect 163262 334294 163358 334350
rect 162738 334226 163358 334294
rect 162738 334170 162834 334226
rect 162890 334170 162958 334226
rect 163014 334170 163082 334226
rect 163138 334170 163206 334226
rect 163262 334170 163358 334226
rect 162738 334102 163358 334170
rect 162738 334046 162834 334102
rect 162890 334046 162958 334102
rect 163014 334046 163082 334102
rect 163138 334046 163206 334102
rect 163262 334046 163358 334102
rect 162738 333978 163358 334046
rect 162738 333922 162834 333978
rect 162890 333922 162958 333978
rect 163014 333922 163082 333978
rect 163138 333922 163206 333978
rect 163262 333922 163358 333978
rect 162738 316350 163358 333922
rect 162738 316294 162834 316350
rect 162890 316294 162958 316350
rect 163014 316294 163082 316350
rect 163138 316294 163206 316350
rect 163262 316294 163358 316350
rect 162738 316226 163358 316294
rect 162738 316170 162834 316226
rect 162890 316170 162958 316226
rect 163014 316170 163082 316226
rect 163138 316170 163206 316226
rect 163262 316170 163358 316226
rect 162738 316102 163358 316170
rect 162738 316046 162834 316102
rect 162890 316046 162958 316102
rect 163014 316046 163082 316102
rect 163138 316046 163206 316102
rect 163262 316046 163358 316102
rect 162738 315978 163358 316046
rect 162738 315922 162834 315978
rect 162890 315922 162958 315978
rect 163014 315922 163082 315978
rect 163138 315922 163206 315978
rect 163262 315922 163358 315978
rect 162738 298350 163358 315922
rect 162738 298294 162834 298350
rect 162890 298294 162958 298350
rect 163014 298294 163082 298350
rect 163138 298294 163206 298350
rect 163262 298294 163358 298350
rect 162738 298226 163358 298294
rect 162738 298170 162834 298226
rect 162890 298170 162958 298226
rect 163014 298170 163082 298226
rect 163138 298170 163206 298226
rect 163262 298170 163358 298226
rect 162738 298102 163358 298170
rect 162738 298046 162834 298102
rect 162890 298046 162958 298102
rect 163014 298046 163082 298102
rect 163138 298046 163206 298102
rect 163262 298046 163358 298102
rect 162738 297978 163358 298046
rect 162738 297922 162834 297978
rect 162890 297922 162958 297978
rect 163014 297922 163082 297978
rect 163138 297922 163206 297978
rect 163262 297922 163358 297978
rect 162738 280350 163358 297922
rect 162738 280294 162834 280350
rect 162890 280294 162958 280350
rect 163014 280294 163082 280350
rect 163138 280294 163206 280350
rect 163262 280294 163358 280350
rect 162738 280226 163358 280294
rect 162738 280170 162834 280226
rect 162890 280170 162958 280226
rect 163014 280170 163082 280226
rect 163138 280170 163206 280226
rect 163262 280170 163358 280226
rect 162738 280102 163358 280170
rect 162738 280046 162834 280102
rect 162890 280046 162958 280102
rect 163014 280046 163082 280102
rect 163138 280046 163206 280102
rect 163262 280046 163358 280102
rect 162738 279978 163358 280046
rect 162738 279922 162834 279978
rect 162890 279922 162958 279978
rect 163014 279922 163082 279978
rect 163138 279922 163206 279978
rect 163262 279922 163358 279978
rect 162738 262350 163358 279922
rect 162738 262294 162834 262350
rect 162890 262294 162958 262350
rect 163014 262294 163082 262350
rect 163138 262294 163206 262350
rect 163262 262294 163358 262350
rect 162738 262226 163358 262294
rect 162738 262170 162834 262226
rect 162890 262170 162958 262226
rect 163014 262170 163082 262226
rect 163138 262170 163206 262226
rect 163262 262170 163358 262226
rect 162738 262102 163358 262170
rect 162738 262046 162834 262102
rect 162890 262046 162958 262102
rect 163014 262046 163082 262102
rect 163138 262046 163206 262102
rect 163262 262046 163358 262102
rect 162738 261978 163358 262046
rect 162738 261922 162834 261978
rect 162890 261922 162958 261978
rect 163014 261922 163082 261978
rect 163138 261922 163206 261978
rect 163262 261922 163358 261978
rect 162738 244350 163358 261922
rect 162738 244294 162834 244350
rect 162890 244294 162958 244350
rect 163014 244294 163082 244350
rect 163138 244294 163206 244350
rect 163262 244294 163358 244350
rect 162738 244226 163358 244294
rect 162738 244170 162834 244226
rect 162890 244170 162958 244226
rect 163014 244170 163082 244226
rect 163138 244170 163206 244226
rect 163262 244170 163358 244226
rect 162738 244102 163358 244170
rect 162738 244046 162834 244102
rect 162890 244046 162958 244102
rect 163014 244046 163082 244102
rect 163138 244046 163206 244102
rect 163262 244046 163358 244102
rect 162738 243978 163358 244046
rect 162738 243922 162834 243978
rect 162890 243922 162958 243978
rect 163014 243922 163082 243978
rect 163138 243922 163206 243978
rect 163262 243922 163358 243978
rect 162738 226350 163358 243922
rect 162738 226294 162834 226350
rect 162890 226294 162958 226350
rect 163014 226294 163082 226350
rect 163138 226294 163206 226350
rect 163262 226294 163358 226350
rect 162738 226226 163358 226294
rect 162738 226170 162834 226226
rect 162890 226170 162958 226226
rect 163014 226170 163082 226226
rect 163138 226170 163206 226226
rect 163262 226170 163358 226226
rect 162738 226102 163358 226170
rect 162738 226046 162834 226102
rect 162890 226046 162958 226102
rect 163014 226046 163082 226102
rect 163138 226046 163206 226102
rect 163262 226046 163358 226102
rect 162738 225978 163358 226046
rect 162738 225922 162834 225978
rect 162890 225922 162958 225978
rect 163014 225922 163082 225978
rect 163138 225922 163206 225978
rect 163262 225922 163358 225978
rect 162738 208350 163358 225922
rect 162738 208294 162834 208350
rect 162890 208294 162958 208350
rect 163014 208294 163082 208350
rect 163138 208294 163206 208350
rect 163262 208294 163358 208350
rect 162738 208226 163358 208294
rect 162738 208170 162834 208226
rect 162890 208170 162958 208226
rect 163014 208170 163082 208226
rect 163138 208170 163206 208226
rect 163262 208170 163358 208226
rect 162738 208102 163358 208170
rect 162738 208046 162834 208102
rect 162890 208046 162958 208102
rect 163014 208046 163082 208102
rect 163138 208046 163206 208102
rect 163262 208046 163358 208102
rect 162738 207978 163358 208046
rect 162738 207922 162834 207978
rect 162890 207922 162958 207978
rect 163014 207922 163082 207978
rect 163138 207922 163206 207978
rect 163262 207922 163358 207978
rect 162738 190350 163358 207922
rect 162738 190294 162834 190350
rect 162890 190294 162958 190350
rect 163014 190294 163082 190350
rect 163138 190294 163206 190350
rect 163262 190294 163358 190350
rect 162738 190226 163358 190294
rect 162738 190170 162834 190226
rect 162890 190170 162958 190226
rect 163014 190170 163082 190226
rect 163138 190170 163206 190226
rect 163262 190170 163358 190226
rect 162738 190102 163358 190170
rect 162738 190046 162834 190102
rect 162890 190046 162958 190102
rect 163014 190046 163082 190102
rect 163138 190046 163206 190102
rect 163262 190046 163358 190102
rect 162738 189978 163358 190046
rect 162738 189922 162834 189978
rect 162890 189922 162958 189978
rect 163014 189922 163082 189978
rect 163138 189922 163206 189978
rect 163262 189922 163358 189978
rect 162738 172350 163358 189922
rect 162738 172294 162834 172350
rect 162890 172294 162958 172350
rect 163014 172294 163082 172350
rect 163138 172294 163206 172350
rect 163262 172294 163358 172350
rect 162738 172226 163358 172294
rect 162738 172170 162834 172226
rect 162890 172170 162958 172226
rect 163014 172170 163082 172226
rect 163138 172170 163206 172226
rect 163262 172170 163358 172226
rect 162738 172102 163358 172170
rect 162738 172046 162834 172102
rect 162890 172046 162958 172102
rect 163014 172046 163082 172102
rect 163138 172046 163206 172102
rect 163262 172046 163358 172102
rect 162738 171978 163358 172046
rect 162738 171922 162834 171978
rect 162890 171922 162958 171978
rect 163014 171922 163082 171978
rect 163138 171922 163206 171978
rect 163262 171922 163358 171978
rect 162738 154350 163358 171922
rect 162738 154294 162834 154350
rect 162890 154294 162958 154350
rect 163014 154294 163082 154350
rect 163138 154294 163206 154350
rect 163262 154294 163358 154350
rect 162738 154226 163358 154294
rect 162738 154170 162834 154226
rect 162890 154170 162958 154226
rect 163014 154170 163082 154226
rect 163138 154170 163206 154226
rect 163262 154170 163358 154226
rect 162738 154102 163358 154170
rect 162738 154046 162834 154102
rect 162890 154046 162958 154102
rect 163014 154046 163082 154102
rect 163138 154046 163206 154102
rect 163262 154046 163358 154102
rect 162738 153978 163358 154046
rect 162738 153922 162834 153978
rect 162890 153922 162958 153978
rect 163014 153922 163082 153978
rect 163138 153922 163206 153978
rect 163262 153922 163358 153978
rect 162738 136350 163358 153922
rect 162738 136294 162834 136350
rect 162890 136294 162958 136350
rect 163014 136294 163082 136350
rect 163138 136294 163206 136350
rect 163262 136294 163358 136350
rect 162738 136226 163358 136294
rect 162738 136170 162834 136226
rect 162890 136170 162958 136226
rect 163014 136170 163082 136226
rect 163138 136170 163206 136226
rect 163262 136170 163358 136226
rect 162738 136102 163358 136170
rect 162738 136046 162834 136102
rect 162890 136046 162958 136102
rect 163014 136046 163082 136102
rect 163138 136046 163206 136102
rect 163262 136046 163358 136102
rect 162738 135978 163358 136046
rect 162738 135922 162834 135978
rect 162890 135922 162958 135978
rect 163014 135922 163082 135978
rect 163138 135922 163206 135978
rect 163262 135922 163358 135978
rect 162738 118350 163358 135922
rect 162738 118294 162834 118350
rect 162890 118294 162958 118350
rect 163014 118294 163082 118350
rect 163138 118294 163206 118350
rect 163262 118294 163358 118350
rect 162738 118226 163358 118294
rect 162738 118170 162834 118226
rect 162890 118170 162958 118226
rect 163014 118170 163082 118226
rect 163138 118170 163206 118226
rect 163262 118170 163358 118226
rect 162738 118102 163358 118170
rect 162738 118046 162834 118102
rect 162890 118046 162958 118102
rect 163014 118046 163082 118102
rect 163138 118046 163206 118102
rect 163262 118046 163358 118102
rect 162738 117978 163358 118046
rect 162738 117922 162834 117978
rect 162890 117922 162958 117978
rect 163014 117922 163082 117978
rect 163138 117922 163206 117978
rect 163262 117922 163358 117978
rect 162738 100350 163358 117922
rect 162738 100294 162834 100350
rect 162890 100294 162958 100350
rect 163014 100294 163082 100350
rect 163138 100294 163206 100350
rect 163262 100294 163358 100350
rect 162738 100226 163358 100294
rect 162738 100170 162834 100226
rect 162890 100170 162958 100226
rect 163014 100170 163082 100226
rect 163138 100170 163206 100226
rect 163262 100170 163358 100226
rect 162738 100102 163358 100170
rect 162738 100046 162834 100102
rect 162890 100046 162958 100102
rect 163014 100046 163082 100102
rect 163138 100046 163206 100102
rect 163262 100046 163358 100102
rect 162738 99978 163358 100046
rect 162738 99922 162834 99978
rect 162890 99922 162958 99978
rect 163014 99922 163082 99978
rect 163138 99922 163206 99978
rect 163262 99922 163358 99978
rect 162738 82350 163358 99922
rect 162738 82294 162834 82350
rect 162890 82294 162958 82350
rect 163014 82294 163082 82350
rect 163138 82294 163206 82350
rect 163262 82294 163358 82350
rect 162738 82226 163358 82294
rect 162738 82170 162834 82226
rect 162890 82170 162958 82226
rect 163014 82170 163082 82226
rect 163138 82170 163206 82226
rect 163262 82170 163358 82226
rect 162738 82102 163358 82170
rect 162738 82046 162834 82102
rect 162890 82046 162958 82102
rect 163014 82046 163082 82102
rect 163138 82046 163206 82102
rect 163262 82046 163358 82102
rect 162738 81978 163358 82046
rect 162738 81922 162834 81978
rect 162890 81922 162958 81978
rect 163014 81922 163082 81978
rect 163138 81922 163206 81978
rect 163262 81922 163358 81978
rect 162738 64350 163358 81922
rect 164668 590212 164724 590222
rect 164668 74998 164724 590156
rect 186508 590212 186564 590222
rect 164668 74932 164724 74942
rect 173852 284676 173908 284686
rect 173852 66724 173908 284620
rect 186508 74818 186564 590156
rect 186508 74752 186564 74762
rect 189738 580350 190358 596784
rect 189738 580294 189834 580350
rect 189890 580294 189958 580350
rect 190014 580294 190082 580350
rect 190138 580294 190206 580350
rect 190262 580294 190358 580350
rect 189738 580226 190358 580294
rect 189738 580170 189834 580226
rect 189890 580170 189958 580226
rect 190014 580170 190082 580226
rect 190138 580170 190206 580226
rect 190262 580170 190358 580226
rect 189738 580102 190358 580170
rect 189738 580046 189834 580102
rect 189890 580046 189958 580102
rect 190014 580046 190082 580102
rect 190138 580046 190206 580102
rect 190262 580046 190358 580102
rect 189738 579978 190358 580046
rect 189738 579922 189834 579978
rect 189890 579922 189958 579978
rect 190014 579922 190082 579978
rect 190138 579922 190206 579978
rect 190262 579922 190358 579978
rect 189738 562350 190358 579922
rect 189738 562294 189834 562350
rect 189890 562294 189958 562350
rect 190014 562294 190082 562350
rect 190138 562294 190206 562350
rect 190262 562294 190358 562350
rect 189738 562226 190358 562294
rect 189738 562170 189834 562226
rect 189890 562170 189958 562226
rect 190014 562170 190082 562226
rect 190138 562170 190206 562226
rect 190262 562170 190358 562226
rect 189738 562102 190358 562170
rect 189738 562046 189834 562102
rect 189890 562046 189958 562102
rect 190014 562046 190082 562102
rect 190138 562046 190206 562102
rect 190262 562046 190358 562102
rect 189738 561978 190358 562046
rect 189738 561922 189834 561978
rect 189890 561922 189958 561978
rect 190014 561922 190082 561978
rect 190138 561922 190206 561978
rect 190262 561922 190358 561978
rect 189738 544350 190358 561922
rect 189738 544294 189834 544350
rect 189890 544294 189958 544350
rect 190014 544294 190082 544350
rect 190138 544294 190206 544350
rect 190262 544294 190358 544350
rect 189738 544226 190358 544294
rect 189738 544170 189834 544226
rect 189890 544170 189958 544226
rect 190014 544170 190082 544226
rect 190138 544170 190206 544226
rect 190262 544170 190358 544226
rect 189738 544102 190358 544170
rect 189738 544046 189834 544102
rect 189890 544046 189958 544102
rect 190014 544046 190082 544102
rect 190138 544046 190206 544102
rect 190262 544046 190358 544102
rect 189738 543978 190358 544046
rect 189738 543922 189834 543978
rect 189890 543922 189958 543978
rect 190014 543922 190082 543978
rect 190138 543922 190206 543978
rect 190262 543922 190358 543978
rect 189738 526350 190358 543922
rect 189738 526294 189834 526350
rect 189890 526294 189958 526350
rect 190014 526294 190082 526350
rect 190138 526294 190206 526350
rect 190262 526294 190358 526350
rect 189738 526226 190358 526294
rect 189738 526170 189834 526226
rect 189890 526170 189958 526226
rect 190014 526170 190082 526226
rect 190138 526170 190206 526226
rect 190262 526170 190358 526226
rect 189738 526102 190358 526170
rect 189738 526046 189834 526102
rect 189890 526046 189958 526102
rect 190014 526046 190082 526102
rect 190138 526046 190206 526102
rect 190262 526046 190358 526102
rect 189738 525978 190358 526046
rect 189738 525922 189834 525978
rect 189890 525922 189958 525978
rect 190014 525922 190082 525978
rect 190138 525922 190206 525978
rect 190262 525922 190358 525978
rect 189738 508350 190358 525922
rect 189738 508294 189834 508350
rect 189890 508294 189958 508350
rect 190014 508294 190082 508350
rect 190138 508294 190206 508350
rect 190262 508294 190358 508350
rect 189738 508226 190358 508294
rect 189738 508170 189834 508226
rect 189890 508170 189958 508226
rect 190014 508170 190082 508226
rect 190138 508170 190206 508226
rect 190262 508170 190358 508226
rect 189738 508102 190358 508170
rect 189738 508046 189834 508102
rect 189890 508046 189958 508102
rect 190014 508046 190082 508102
rect 190138 508046 190206 508102
rect 190262 508046 190358 508102
rect 189738 507978 190358 508046
rect 189738 507922 189834 507978
rect 189890 507922 189958 507978
rect 190014 507922 190082 507978
rect 190138 507922 190206 507978
rect 190262 507922 190358 507978
rect 189738 490350 190358 507922
rect 189738 490294 189834 490350
rect 189890 490294 189958 490350
rect 190014 490294 190082 490350
rect 190138 490294 190206 490350
rect 190262 490294 190358 490350
rect 189738 490226 190358 490294
rect 189738 490170 189834 490226
rect 189890 490170 189958 490226
rect 190014 490170 190082 490226
rect 190138 490170 190206 490226
rect 190262 490170 190358 490226
rect 189738 490102 190358 490170
rect 189738 490046 189834 490102
rect 189890 490046 189958 490102
rect 190014 490046 190082 490102
rect 190138 490046 190206 490102
rect 190262 490046 190358 490102
rect 189738 489978 190358 490046
rect 189738 489922 189834 489978
rect 189890 489922 189958 489978
rect 190014 489922 190082 489978
rect 190138 489922 190206 489978
rect 190262 489922 190358 489978
rect 189738 472350 190358 489922
rect 189738 472294 189834 472350
rect 189890 472294 189958 472350
rect 190014 472294 190082 472350
rect 190138 472294 190206 472350
rect 190262 472294 190358 472350
rect 189738 472226 190358 472294
rect 189738 472170 189834 472226
rect 189890 472170 189958 472226
rect 190014 472170 190082 472226
rect 190138 472170 190206 472226
rect 190262 472170 190358 472226
rect 189738 472102 190358 472170
rect 189738 472046 189834 472102
rect 189890 472046 189958 472102
rect 190014 472046 190082 472102
rect 190138 472046 190206 472102
rect 190262 472046 190358 472102
rect 189738 471978 190358 472046
rect 189738 471922 189834 471978
rect 189890 471922 189958 471978
rect 190014 471922 190082 471978
rect 190138 471922 190206 471978
rect 190262 471922 190358 471978
rect 189738 454350 190358 471922
rect 189738 454294 189834 454350
rect 189890 454294 189958 454350
rect 190014 454294 190082 454350
rect 190138 454294 190206 454350
rect 190262 454294 190358 454350
rect 189738 454226 190358 454294
rect 189738 454170 189834 454226
rect 189890 454170 189958 454226
rect 190014 454170 190082 454226
rect 190138 454170 190206 454226
rect 190262 454170 190358 454226
rect 189738 454102 190358 454170
rect 189738 454046 189834 454102
rect 189890 454046 189958 454102
rect 190014 454046 190082 454102
rect 190138 454046 190206 454102
rect 190262 454046 190358 454102
rect 189738 453978 190358 454046
rect 189738 453922 189834 453978
rect 189890 453922 189958 453978
rect 190014 453922 190082 453978
rect 190138 453922 190206 453978
rect 190262 453922 190358 453978
rect 189738 436350 190358 453922
rect 189738 436294 189834 436350
rect 189890 436294 189958 436350
rect 190014 436294 190082 436350
rect 190138 436294 190206 436350
rect 190262 436294 190358 436350
rect 189738 436226 190358 436294
rect 189738 436170 189834 436226
rect 189890 436170 189958 436226
rect 190014 436170 190082 436226
rect 190138 436170 190206 436226
rect 190262 436170 190358 436226
rect 189738 436102 190358 436170
rect 189738 436046 189834 436102
rect 189890 436046 189958 436102
rect 190014 436046 190082 436102
rect 190138 436046 190206 436102
rect 190262 436046 190358 436102
rect 189738 435978 190358 436046
rect 189738 435922 189834 435978
rect 189890 435922 189958 435978
rect 190014 435922 190082 435978
rect 190138 435922 190206 435978
rect 190262 435922 190358 435978
rect 189738 418350 190358 435922
rect 189738 418294 189834 418350
rect 189890 418294 189958 418350
rect 190014 418294 190082 418350
rect 190138 418294 190206 418350
rect 190262 418294 190358 418350
rect 189738 418226 190358 418294
rect 189738 418170 189834 418226
rect 189890 418170 189958 418226
rect 190014 418170 190082 418226
rect 190138 418170 190206 418226
rect 190262 418170 190358 418226
rect 189738 418102 190358 418170
rect 189738 418046 189834 418102
rect 189890 418046 189958 418102
rect 190014 418046 190082 418102
rect 190138 418046 190206 418102
rect 190262 418046 190358 418102
rect 189738 417978 190358 418046
rect 189738 417922 189834 417978
rect 189890 417922 189958 417978
rect 190014 417922 190082 417978
rect 190138 417922 190206 417978
rect 190262 417922 190358 417978
rect 189738 400350 190358 417922
rect 189738 400294 189834 400350
rect 189890 400294 189958 400350
rect 190014 400294 190082 400350
rect 190138 400294 190206 400350
rect 190262 400294 190358 400350
rect 189738 400226 190358 400294
rect 189738 400170 189834 400226
rect 189890 400170 189958 400226
rect 190014 400170 190082 400226
rect 190138 400170 190206 400226
rect 190262 400170 190358 400226
rect 189738 400102 190358 400170
rect 189738 400046 189834 400102
rect 189890 400046 189958 400102
rect 190014 400046 190082 400102
rect 190138 400046 190206 400102
rect 190262 400046 190358 400102
rect 189738 399978 190358 400046
rect 189738 399922 189834 399978
rect 189890 399922 189958 399978
rect 190014 399922 190082 399978
rect 190138 399922 190206 399978
rect 190262 399922 190358 399978
rect 189738 382350 190358 399922
rect 189738 382294 189834 382350
rect 189890 382294 189958 382350
rect 190014 382294 190082 382350
rect 190138 382294 190206 382350
rect 190262 382294 190358 382350
rect 189738 382226 190358 382294
rect 189738 382170 189834 382226
rect 189890 382170 189958 382226
rect 190014 382170 190082 382226
rect 190138 382170 190206 382226
rect 190262 382170 190358 382226
rect 189738 382102 190358 382170
rect 189738 382046 189834 382102
rect 189890 382046 189958 382102
rect 190014 382046 190082 382102
rect 190138 382046 190206 382102
rect 190262 382046 190358 382102
rect 189738 381978 190358 382046
rect 189738 381922 189834 381978
rect 189890 381922 189958 381978
rect 190014 381922 190082 381978
rect 190138 381922 190206 381978
rect 190262 381922 190358 381978
rect 189738 364350 190358 381922
rect 189738 364294 189834 364350
rect 189890 364294 189958 364350
rect 190014 364294 190082 364350
rect 190138 364294 190206 364350
rect 190262 364294 190358 364350
rect 189738 364226 190358 364294
rect 189738 364170 189834 364226
rect 189890 364170 189958 364226
rect 190014 364170 190082 364226
rect 190138 364170 190206 364226
rect 190262 364170 190358 364226
rect 189738 364102 190358 364170
rect 189738 364046 189834 364102
rect 189890 364046 189958 364102
rect 190014 364046 190082 364102
rect 190138 364046 190206 364102
rect 190262 364046 190358 364102
rect 189738 363978 190358 364046
rect 189738 363922 189834 363978
rect 189890 363922 189958 363978
rect 190014 363922 190082 363978
rect 190138 363922 190206 363978
rect 190262 363922 190358 363978
rect 189738 346350 190358 363922
rect 189738 346294 189834 346350
rect 189890 346294 189958 346350
rect 190014 346294 190082 346350
rect 190138 346294 190206 346350
rect 190262 346294 190358 346350
rect 189738 346226 190358 346294
rect 189738 346170 189834 346226
rect 189890 346170 189958 346226
rect 190014 346170 190082 346226
rect 190138 346170 190206 346226
rect 190262 346170 190358 346226
rect 189738 346102 190358 346170
rect 189738 346046 189834 346102
rect 189890 346046 189958 346102
rect 190014 346046 190082 346102
rect 190138 346046 190206 346102
rect 190262 346046 190358 346102
rect 189738 345978 190358 346046
rect 189738 345922 189834 345978
rect 189890 345922 189958 345978
rect 190014 345922 190082 345978
rect 190138 345922 190206 345978
rect 190262 345922 190358 345978
rect 189738 328350 190358 345922
rect 189738 328294 189834 328350
rect 189890 328294 189958 328350
rect 190014 328294 190082 328350
rect 190138 328294 190206 328350
rect 190262 328294 190358 328350
rect 189738 328226 190358 328294
rect 189738 328170 189834 328226
rect 189890 328170 189958 328226
rect 190014 328170 190082 328226
rect 190138 328170 190206 328226
rect 190262 328170 190358 328226
rect 189738 328102 190358 328170
rect 189738 328046 189834 328102
rect 189890 328046 189958 328102
rect 190014 328046 190082 328102
rect 190138 328046 190206 328102
rect 190262 328046 190358 328102
rect 189738 327978 190358 328046
rect 189738 327922 189834 327978
rect 189890 327922 189958 327978
rect 190014 327922 190082 327978
rect 190138 327922 190206 327978
rect 190262 327922 190358 327978
rect 189738 310350 190358 327922
rect 189738 310294 189834 310350
rect 189890 310294 189958 310350
rect 190014 310294 190082 310350
rect 190138 310294 190206 310350
rect 190262 310294 190358 310350
rect 189738 310226 190358 310294
rect 189738 310170 189834 310226
rect 189890 310170 189958 310226
rect 190014 310170 190082 310226
rect 190138 310170 190206 310226
rect 190262 310170 190358 310226
rect 189738 310102 190358 310170
rect 189738 310046 189834 310102
rect 189890 310046 189958 310102
rect 190014 310046 190082 310102
rect 190138 310046 190206 310102
rect 190262 310046 190358 310102
rect 189738 309978 190358 310046
rect 189738 309922 189834 309978
rect 189890 309922 189958 309978
rect 190014 309922 190082 309978
rect 190138 309922 190206 309978
rect 190262 309922 190358 309978
rect 189738 292350 190358 309922
rect 189738 292294 189834 292350
rect 189890 292294 189958 292350
rect 190014 292294 190082 292350
rect 190138 292294 190206 292350
rect 190262 292294 190358 292350
rect 189738 292226 190358 292294
rect 189738 292170 189834 292226
rect 189890 292170 189958 292226
rect 190014 292170 190082 292226
rect 190138 292170 190206 292226
rect 190262 292170 190358 292226
rect 189738 292102 190358 292170
rect 189738 292046 189834 292102
rect 189890 292046 189958 292102
rect 190014 292046 190082 292102
rect 190138 292046 190206 292102
rect 190262 292046 190358 292102
rect 189738 291978 190358 292046
rect 189738 291922 189834 291978
rect 189890 291922 189958 291978
rect 190014 291922 190082 291978
rect 190138 291922 190206 291978
rect 190262 291922 190358 291978
rect 189738 274350 190358 291922
rect 189738 274294 189834 274350
rect 189890 274294 189958 274350
rect 190014 274294 190082 274350
rect 190138 274294 190206 274350
rect 190262 274294 190358 274350
rect 189738 274226 190358 274294
rect 189738 274170 189834 274226
rect 189890 274170 189958 274226
rect 190014 274170 190082 274226
rect 190138 274170 190206 274226
rect 190262 274170 190358 274226
rect 189738 274102 190358 274170
rect 189738 274046 189834 274102
rect 189890 274046 189958 274102
rect 190014 274046 190082 274102
rect 190138 274046 190206 274102
rect 190262 274046 190358 274102
rect 189738 273978 190358 274046
rect 189738 273922 189834 273978
rect 189890 273922 189958 273978
rect 190014 273922 190082 273978
rect 190138 273922 190206 273978
rect 190262 273922 190358 273978
rect 189738 256350 190358 273922
rect 189738 256294 189834 256350
rect 189890 256294 189958 256350
rect 190014 256294 190082 256350
rect 190138 256294 190206 256350
rect 190262 256294 190358 256350
rect 189738 256226 190358 256294
rect 189738 256170 189834 256226
rect 189890 256170 189958 256226
rect 190014 256170 190082 256226
rect 190138 256170 190206 256226
rect 190262 256170 190358 256226
rect 189738 256102 190358 256170
rect 189738 256046 189834 256102
rect 189890 256046 189958 256102
rect 190014 256046 190082 256102
rect 190138 256046 190206 256102
rect 190262 256046 190358 256102
rect 189738 255978 190358 256046
rect 189738 255922 189834 255978
rect 189890 255922 189958 255978
rect 190014 255922 190082 255978
rect 190138 255922 190206 255978
rect 190262 255922 190358 255978
rect 189738 238350 190358 255922
rect 189738 238294 189834 238350
rect 189890 238294 189958 238350
rect 190014 238294 190082 238350
rect 190138 238294 190206 238350
rect 190262 238294 190358 238350
rect 189738 238226 190358 238294
rect 189738 238170 189834 238226
rect 189890 238170 189958 238226
rect 190014 238170 190082 238226
rect 190138 238170 190206 238226
rect 190262 238170 190358 238226
rect 189738 238102 190358 238170
rect 189738 238046 189834 238102
rect 189890 238046 189958 238102
rect 190014 238046 190082 238102
rect 190138 238046 190206 238102
rect 190262 238046 190358 238102
rect 189738 237978 190358 238046
rect 189738 237922 189834 237978
rect 189890 237922 189958 237978
rect 190014 237922 190082 237978
rect 190138 237922 190206 237978
rect 190262 237922 190358 237978
rect 189738 220350 190358 237922
rect 189738 220294 189834 220350
rect 189890 220294 189958 220350
rect 190014 220294 190082 220350
rect 190138 220294 190206 220350
rect 190262 220294 190358 220350
rect 189738 220226 190358 220294
rect 189738 220170 189834 220226
rect 189890 220170 189958 220226
rect 190014 220170 190082 220226
rect 190138 220170 190206 220226
rect 190262 220170 190358 220226
rect 189738 220102 190358 220170
rect 189738 220046 189834 220102
rect 189890 220046 189958 220102
rect 190014 220046 190082 220102
rect 190138 220046 190206 220102
rect 190262 220046 190358 220102
rect 189738 219978 190358 220046
rect 189738 219922 189834 219978
rect 189890 219922 189958 219978
rect 190014 219922 190082 219978
rect 190138 219922 190206 219978
rect 190262 219922 190358 219978
rect 189738 202350 190358 219922
rect 189738 202294 189834 202350
rect 189890 202294 189958 202350
rect 190014 202294 190082 202350
rect 190138 202294 190206 202350
rect 190262 202294 190358 202350
rect 189738 202226 190358 202294
rect 189738 202170 189834 202226
rect 189890 202170 189958 202226
rect 190014 202170 190082 202226
rect 190138 202170 190206 202226
rect 190262 202170 190358 202226
rect 189738 202102 190358 202170
rect 189738 202046 189834 202102
rect 189890 202046 189958 202102
rect 190014 202046 190082 202102
rect 190138 202046 190206 202102
rect 190262 202046 190358 202102
rect 189738 201978 190358 202046
rect 189738 201922 189834 201978
rect 189890 201922 189958 201978
rect 190014 201922 190082 201978
rect 190138 201922 190206 201978
rect 190262 201922 190358 201978
rect 189738 184350 190358 201922
rect 189738 184294 189834 184350
rect 189890 184294 189958 184350
rect 190014 184294 190082 184350
rect 190138 184294 190206 184350
rect 190262 184294 190358 184350
rect 189738 184226 190358 184294
rect 189738 184170 189834 184226
rect 189890 184170 189958 184226
rect 190014 184170 190082 184226
rect 190138 184170 190206 184226
rect 190262 184170 190358 184226
rect 189738 184102 190358 184170
rect 189738 184046 189834 184102
rect 189890 184046 189958 184102
rect 190014 184046 190082 184102
rect 190138 184046 190206 184102
rect 190262 184046 190358 184102
rect 189738 183978 190358 184046
rect 189738 183922 189834 183978
rect 189890 183922 189958 183978
rect 190014 183922 190082 183978
rect 190138 183922 190206 183978
rect 190262 183922 190358 183978
rect 189738 166350 190358 183922
rect 189738 166294 189834 166350
rect 189890 166294 189958 166350
rect 190014 166294 190082 166350
rect 190138 166294 190206 166350
rect 190262 166294 190358 166350
rect 189738 166226 190358 166294
rect 189738 166170 189834 166226
rect 189890 166170 189958 166226
rect 190014 166170 190082 166226
rect 190138 166170 190206 166226
rect 190262 166170 190358 166226
rect 189738 166102 190358 166170
rect 189738 166046 189834 166102
rect 189890 166046 189958 166102
rect 190014 166046 190082 166102
rect 190138 166046 190206 166102
rect 190262 166046 190358 166102
rect 189738 165978 190358 166046
rect 189738 165922 189834 165978
rect 189890 165922 189958 165978
rect 190014 165922 190082 165978
rect 190138 165922 190206 165978
rect 190262 165922 190358 165978
rect 189738 148350 190358 165922
rect 189738 148294 189834 148350
rect 189890 148294 189958 148350
rect 190014 148294 190082 148350
rect 190138 148294 190206 148350
rect 190262 148294 190358 148350
rect 189738 148226 190358 148294
rect 189738 148170 189834 148226
rect 189890 148170 189958 148226
rect 190014 148170 190082 148226
rect 190138 148170 190206 148226
rect 190262 148170 190358 148226
rect 189738 148102 190358 148170
rect 189738 148046 189834 148102
rect 189890 148046 189958 148102
rect 190014 148046 190082 148102
rect 190138 148046 190206 148102
rect 190262 148046 190358 148102
rect 189738 147978 190358 148046
rect 189738 147922 189834 147978
rect 189890 147922 189958 147978
rect 190014 147922 190082 147978
rect 190138 147922 190206 147978
rect 190262 147922 190358 147978
rect 189738 130350 190358 147922
rect 189738 130294 189834 130350
rect 189890 130294 189958 130350
rect 190014 130294 190082 130350
rect 190138 130294 190206 130350
rect 190262 130294 190358 130350
rect 189738 130226 190358 130294
rect 189738 130170 189834 130226
rect 189890 130170 189958 130226
rect 190014 130170 190082 130226
rect 190138 130170 190206 130226
rect 190262 130170 190358 130226
rect 189738 130102 190358 130170
rect 189738 130046 189834 130102
rect 189890 130046 189958 130102
rect 190014 130046 190082 130102
rect 190138 130046 190206 130102
rect 190262 130046 190358 130102
rect 189738 129978 190358 130046
rect 189738 129922 189834 129978
rect 189890 129922 189958 129978
rect 190014 129922 190082 129978
rect 190138 129922 190206 129978
rect 190262 129922 190358 129978
rect 189738 112350 190358 129922
rect 189738 112294 189834 112350
rect 189890 112294 189958 112350
rect 190014 112294 190082 112350
rect 190138 112294 190206 112350
rect 190262 112294 190358 112350
rect 189738 112226 190358 112294
rect 189738 112170 189834 112226
rect 189890 112170 189958 112226
rect 190014 112170 190082 112226
rect 190138 112170 190206 112226
rect 190262 112170 190358 112226
rect 189738 112102 190358 112170
rect 189738 112046 189834 112102
rect 189890 112046 189958 112102
rect 190014 112046 190082 112102
rect 190138 112046 190206 112102
rect 190262 112046 190358 112102
rect 189738 111978 190358 112046
rect 189738 111922 189834 111978
rect 189890 111922 189958 111978
rect 190014 111922 190082 111978
rect 190138 111922 190206 111978
rect 190262 111922 190358 111978
rect 189738 94350 190358 111922
rect 189738 94294 189834 94350
rect 189890 94294 189958 94350
rect 190014 94294 190082 94350
rect 190138 94294 190206 94350
rect 190262 94294 190358 94350
rect 189738 94226 190358 94294
rect 189738 94170 189834 94226
rect 189890 94170 189958 94226
rect 190014 94170 190082 94226
rect 190138 94170 190206 94226
rect 190262 94170 190358 94226
rect 189738 94102 190358 94170
rect 189738 94046 189834 94102
rect 189890 94046 189958 94102
rect 190014 94046 190082 94102
rect 190138 94046 190206 94102
rect 190262 94046 190358 94102
rect 189738 93978 190358 94046
rect 189738 93922 189834 93978
rect 189890 93922 189958 93978
rect 190014 93922 190082 93978
rect 190138 93922 190206 93978
rect 190262 93922 190358 93978
rect 189738 76350 190358 93922
rect 189738 76294 189834 76350
rect 189890 76294 189958 76350
rect 190014 76294 190082 76350
rect 190138 76294 190206 76350
rect 190262 76294 190358 76350
rect 189738 76226 190358 76294
rect 189738 76170 189834 76226
rect 189890 76170 189958 76226
rect 190014 76170 190082 76226
rect 190138 76170 190206 76226
rect 190262 76170 190358 76226
rect 189738 76102 190358 76170
rect 189738 76046 189834 76102
rect 189890 76046 189958 76102
rect 190014 76046 190082 76102
rect 190138 76046 190206 76102
rect 190262 76046 190358 76102
rect 189738 75978 190358 76046
rect 189738 75922 189834 75978
rect 189890 75922 189958 75978
rect 190014 75922 190082 75978
rect 190138 75922 190206 75978
rect 190262 75922 190358 75978
rect 173852 66658 173908 66668
rect 162738 64294 162834 64350
rect 162890 64294 162958 64350
rect 163014 64294 163082 64350
rect 163138 64294 163206 64350
rect 163262 64294 163358 64350
rect 162738 64226 163358 64294
rect 162738 64170 162834 64226
rect 162890 64170 162958 64226
rect 163014 64170 163082 64226
rect 163138 64170 163206 64226
rect 163262 64170 163358 64226
rect 162738 64102 163358 64170
rect 162738 64046 162834 64102
rect 162890 64046 162958 64102
rect 163014 64046 163082 64102
rect 163138 64046 163206 64102
rect 163262 64046 163358 64102
rect 162738 63978 163358 64046
rect 162738 63922 162834 63978
rect 162890 63922 162958 63978
rect 163014 63922 163082 63978
rect 163138 63922 163206 63978
rect 163262 63922 163358 63978
rect 162738 46350 163358 63922
rect 162738 46294 162834 46350
rect 162890 46294 162958 46350
rect 163014 46294 163082 46350
rect 163138 46294 163206 46350
rect 163262 46294 163358 46350
rect 162738 46226 163358 46294
rect 162738 46170 162834 46226
rect 162890 46170 162958 46226
rect 163014 46170 163082 46226
rect 163138 46170 163206 46226
rect 163262 46170 163358 46226
rect 162738 46102 163358 46170
rect 162738 46046 162834 46102
rect 162890 46046 162958 46102
rect 163014 46046 163082 46102
rect 163138 46046 163206 46102
rect 163262 46046 163358 46102
rect 162738 45978 163358 46046
rect 162738 45922 162834 45978
rect 162890 45922 162958 45978
rect 163014 45922 163082 45978
rect 163138 45922 163206 45978
rect 163262 45922 163358 45978
rect 162738 28350 163358 45922
rect 166348 61318 166404 61328
rect 162738 28294 162834 28350
rect 162890 28294 162958 28350
rect 163014 28294 163082 28350
rect 163138 28294 163206 28350
rect 163262 28294 163358 28350
rect 162738 28226 163358 28294
rect 162738 28170 162834 28226
rect 162890 28170 162958 28226
rect 163014 28170 163082 28226
rect 163138 28170 163206 28226
rect 163262 28170 163358 28226
rect 162738 28102 163358 28170
rect 162738 28046 162834 28102
rect 162890 28046 162958 28102
rect 163014 28046 163082 28102
rect 163138 28046 163206 28102
rect 163262 28046 163358 28102
rect 162738 27978 163358 28046
rect 162738 27922 162834 27978
rect 162890 27922 162958 27978
rect 163014 27922 163082 27978
rect 163138 27922 163206 27978
rect 163262 27922 163358 27978
rect 159018 4294 159114 4350
rect 159170 4294 159238 4350
rect 159294 4294 159362 4350
rect 159418 4294 159486 4350
rect 159542 4294 159638 4350
rect 159018 4226 159638 4294
rect 159018 4170 159114 4226
rect 159170 4170 159238 4226
rect 159294 4170 159362 4226
rect 159418 4170 159486 4226
rect 159542 4170 159638 4226
rect 132018 -1176 132114 -1120
rect 132170 -1176 132238 -1120
rect 132294 -1176 132362 -1120
rect 132418 -1176 132486 -1120
rect 132542 -1176 132638 -1120
rect 132018 -1244 132638 -1176
rect 132018 -1300 132114 -1244
rect 132170 -1300 132238 -1244
rect 132294 -1300 132362 -1244
rect 132418 -1300 132486 -1244
rect 132542 -1300 132638 -1244
rect 132018 -1368 132638 -1300
rect 132018 -1424 132114 -1368
rect 132170 -1424 132238 -1368
rect 132294 -1424 132362 -1368
rect 132418 -1424 132486 -1368
rect 132542 -1424 132638 -1368
rect 132018 -1492 132638 -1424
rect 132018 -1548 132114 -1492
rect 132170 -1548 132238 -1492
rect 132294 -1548 132362 -1492
rect 132418 -1548 132486 -1492
rect 132542 -1548 132638 -1492
rect 132018 -1644 132638 -1548
rect 159018 4102 159638 4170
rect 161308 14158 161364 14168
rect 161308 4228 161364 14102
rect 161308 4162 161364 4172
rect 162738 10350 163358 27922
rect 162738 10294 162834 10350
rect 162890 10294 162958 10350
rect 163014 10294 163082 10350
rect 163138 10294 163206 10350
rect 163262 10294 163358 10350
rect 162738 10226 163358 10294
rect 162738 10170 162834 10226
rect 162890 10170 162958 10226
rect 163014 10170 163082 10226
rect 163138 10170 163206 10226
rect 163262 10170 163358 10226
rect 162738 10102 163358 10170
rect 162738 10046 162834 10102
rect 162890 10046 162958 10102
rect 163014 10046 163082 10102
rect 163138 10046 163206 10102
rect 163262 10046 163358 10102
rect 162738 9978 163358 10046
rect 162738 9922 162834 9978
rect 162890 9922 162958 9978
rect 163014 9922 163082 9978
rect 163138 9922 163206 9978
rect 163262 9922 163358 9978
rect 159018 4046 159114 4102
rect 159170 4046 159238 4102
rect 159294 4046 159362 4102
rect 159418 4046 159486 4102
rect 159542 4046 159638 4102
rect 159018 3978 159638 4046
rect 159018 3922 159114 3978
rect 159170 3922 159238 3978
rect 159294 3922 159362 3978
rect 159418 3922 159486 3978
rect 159542 3922 159638 3978
rect 159018 -160 159638 3922
rect 159018 -216 159114 -160
rect 159170 -216 159238 -160
rect 159294 -216 159362 -160
rect 159418 -216 159486 -160
rect 159542 -216 159638 -160
rect 159018 -284 159638 -216
rect 159018 -340 159114 -284
rect 159170 -340 159238 -284
rect 159294 -340 159362 -284
rect 159418 -340 159486 -284
rect 159542 -340 159638 -284
rect 159018 -408 159638 -340
rect 159018 -464 159114 -408
rect 159170 -464 159238 -408
rect 159294 -464 159362 -408
rect 159418 -464 159486 -408
rect 159542 -464 159638 -408
rect 159018 -532 159638 -464
rect 159018 -588 159114 -532
rect 159170 -588 159238 -532
rect 159294 -588 159362 -532
rect 159418 -588 159486 -532
rect 159542 -588 159638 -532
rect 159018 -1644 159638 -588
rect 162738 -1120 163358 9922
rect 164668 29098 164724 29108
rect 163660 9118 163716 9128
rect 163660 4228 163716 9062
rect 163660 4162 163716 4172
rect 164668 4228 164724 29042
rect 164668 4162 164724 4172
rect 166348 4228 166404 61262
rect 189738 58350 190358 75922
rect 189738 58294 189834 58350
rect 189890 58294 189958 58350
rect 190014 58294 190082 58350
rect 190138 58294 190206 58350
rect 190262 58294 190358 58350
rect 189738 58226 190358 58294
rect 189738 58170 189834 58226
rect 189890 58170 189958 58226
rect 190014 58170 190082 58226
rect 190138 58170 190206 58226
rect 190262 58170 190358 58226
rect 189738 58102 190358 58170
rect 189738 58046 189834 58102
rect 189890 58046 189958 58102
rect 190014 58046 190082 58102
rect 190138 58046 190206 58102
rect 190262 58046 190358 58102
rect 189738 57978 190358 58046
rect 189738 57922 189834 57978
rect 189890 57922 189958 57978
rect 190014 57922 190082 57978
rect 190138 57922 190206 57978
rect 190262 57922 190358 57978
rect 189738 40350 190358 57922
rect 193458 598172 194078 598268
rect 193458 598116 193554 598172
rect 193610 598116 193678 598172
rect 193734 598116 193802 598172
rect 193858 598116 193926 598172
rect 193982 598116 194078 598172
rect 193458 598048 194078 598116
rect 193458 597992 193554 598048
rect 193610 597992 193678 598048
rect 193734 597992 193802 598048
rect 193858 597992 193926 598048
rect 193982 597992 194078 598048
rect 193458 597924 194078 597992
rect 193458 597868 193554 597924
rect 193610 597868 193678 597924
rect 193734 597868 193802 597924
rect 193858 597868 193926 597924
rect 193982 597868 194078 597924
rect 193458 597800 194078 597868
rect 193458 597744 193554 597800
rect 193610 597744 193678 597800
rect 193734 597744 193802 597800
rect 193858 597744 193926 597800
rect 193982 597744 194078 597800
rect 193458 586350 194078 597744
rect 193458 586294 193554 586350
rect 193610 586294 193678 586350
rect 193734 586294 193802 586350
rect 193858 586294 193926 586350
rect 193982 586294 194078 586350
rect 193458 586226 194078 586294
rect 193458 586170 193554 586226
rect 193610 586170 193678 586226
rect 193734 586170 193802 586226
rect 193858 586170 193926 586226
rect 193982 586170 194078 586226
rect 193458 586102 194078 586170
rect 193458 586046 193554 586102
rect 193610 586046 193678 586102
rect 193734 586046 193802 586102
rect 193858 586046 193926 586102
rect 193982 586046 194078 586102
rect 193458 585978 194078 586046
rect 193458 585922 193554 585978
rect 193610 585922 193678 585978
rect 193734 585922 193802 585978
rect 193858 585922 193926 585978
rect 193982 585922 194078 585978
rect 193458 568350 194078 585922
rect 193458 568294 193554 568350
rect 193610 568294 193678 568350
rect 193734 568294 193802 568350
rect 193858 568294 193926 568350
rect 193982 568294 194078 568350
rect 193458 568226 194078 568294
rect 193458 568170 193554 568226
rect 193610 568170 193678 568226
rect 193734 568170 193802 568226
rect 193858 568170 193926 568226
rect 193982 568170 194078 568226
rect 193458 568102 194078 568170
rect 193458 568046 193554 568102
rect 193610 568046 193678 568102
rect 193734 568046 193802 568102
rect 193858 568046 193926 568102
rect 193982 568046 194078 568102
rect 193458 567978 194078 568046
rect 193458 567922 193554 567978
rect 193610 567922 193678 567978
rect 193734 567922 193802 567978
rect 193858 567922 193926 567978
rect 193982 567922 194078 567978
rect 193458 550350 194078 567922
rect 193458 550294 193554 550350
rect 193610 550294 193678 550350
rect 193734 550294 193802 550350
rect 193858 550294 193926 550350
rect 193982 550294 194078 550350
rect 193458 550226 194078 550294
rect 193458 550170 193554 550226
rect 193610 550170 193678 550226
rect 193734 550170 193802 550226
rect 193858 550170 193926 550226
rect 193982 550170 194078 550226
rect 193458 550102 194078 550170
rect 193458 550046 193554 550102
rect 193610 550046 193678 550102
rect 193734 550046 193802 550102
rect 193858 550046 193926 550102
rect 193982 550046 194078 550102
rect 193458 549978 194078 550046
rect 193458 549922 193554 549978
rect 193610 549922 193678 549978
rect 193734 549922 193802 549978
rect 193858 549922 193926 549978
rect 193982 549922 194078 549978
rect 193458 532350 194078 549922
rect 193458 532294 193554 532350
rect 193610 532294 193678 532350
rect 193734 532294 193802 532350
rect 193858 532294 193926 532350
rect 193982 532294 194078 532350
rect 193458 532226 194078 532294
rect 193458 532170 193554 532226
rect 193610 532170 193678 532226
rect 193734 532170 193802 532226
rect 193858 532170 193926 532226
rect 193982 532170 194078 532226
rect 193458 532102 194078 532170
rect 193458 532046 193554 532102
rect 193610 532046 193678 532102
rect 193734 532046 193802 532102
rect 193858 532046 193926 532102
rect 193982 532046 194078 532102
rect 193458 531978 194078 532046
rect 193458 531922 193554 531978
rect 193610 531922 193678 531978
rect 193734 531922 193802 531978
rect 193858 531922 193926 531978
rect 193982 531922 194078 531978
rect 193458 514350 194078 531922
rect 193458 514294 193554 514350
rect 193610 514294 193678 514350
rect 193734 514294 193802 514350
rect 193858 514294 193926 514350
rect 193982 514294 194078 514350
rect 193458 514226 194078 514294
rect 193458 514170 193554 514226
rect 193610 514170 193678 514226
rect 193734 514170 193802 514226
rect 193858 514170 193926 514226
rect 193982 514170 194078 514226
rect 193458 514102 194078 514170
rect 193458 514046 193554 514102
rect 193610 514046 193678 514102
rect 193734 514046 193802 514102
rect 193858 514046 193926 514102
rect 193982 514046 194078 514102
rect 193458 513978 194078 514046
rect 193458 513922 193554 513978
rect 193610 513922 193678 513978
rect 193734 513922 193802 513978
rect 193858 513922 193926 513978
rect 193982 513922 194078 513978
rect 193458 496350 194078 513922
rect 193458 496294 193554 496350
rect 193610 496294 193678 496350
rect 193734 496294 193802 496350
rect 193858 496294 193926 496350
rect 193982 496294 194078 496350
rect 193458 496226 194078 496294
rect 193458 496170 193554 496226
rect 193610 496170 193678 496226
rect 193734 496170 193802 496226
rect 193858 496170 193926 496226
rect 193982 496170 194078 496226
rect 193458 496102 194078 496170
rect 193458 496046 193554 496102
rect 193610 496046 193678 496102
rect 193734 496046 193802 496102
rect 193858 496046 193926 496102
rect 193982 496046 194078 496102
rect 193458 495978 194078 496046
rect 193458 495922 193554 495978
rect 193610 495922 193678 495978
rect 193734 495922 193802 495978
rect 193858 495922 193926 495978
rect 193982 495922 194078 495978
rect 193458 478350 194078 495922
rect 193458 478294 193554 478350
rect 193610 478294 193678 478350
rect 193734 478294 193802 478350
rect 193858 478294 193926 478350
rect 193982 478294 194078 478350
rect 193458 478226 194078 478294
rect 193458 478170 193554 478226
rect 193610 478170 193678 478226
rect 193734 478170 193802 478226
rect 193858 478170 193926 478226
rect 193982 478170 194078 478226
rect 193458 478102 194078 478170
rect 193458 478046 193554 478102
rect 193610 478046 193678 478102
rect 193734 478046 193802 478102
rect 193858 478046 193926 478102
rect 193982 478046 194078 478102
rect 193458 477978 194078 478046
rect 193458 477922 193554 477978
rect 193610 477922 193678 477978
rect 193734 477922 193802 477978
rect 193858 477922 193926 477978
rect 193982 477922 194078 477978
rect 193458 460350 194078 477922
rect 193458 460294 193554 460350
rect 193610 460294 193678 460350
rect 193734 460294 193802 460350
rect 193858 460294 193926 460350
rect 193982 460294 194078 460350
rect 193458 460226 194078 460294
rect 193458 460170 193554 460226
rect 193610 460170 193678 460226
rect 193734 460170 193802 460226
rect 193858 460170 193926 460226
rect 193982 460170 194078 460226
rect 193458 460102 194078 460170
rect 193458 460046 193554 460102
rect 193610 460046 193678 460102
rect 193734 460046 193802 460102
rect 193858 460046 193926 460102
rect 193982 460046 194078 460102
rect 193458 459978 194078 460046
rect 193458 459922 193554 459978
rect 193610 459922 193678 459978
rect 193734 459922 193802 459978
rect 193858 459922 193926 459978
rect 193982 459922 194078 459978
rect 193458 442350 194078 459922
rect 193458 442294 193554 442350
rect 193610 442294 193678 442350
rect 193734 442294 193802 442350
rect 193858 442294 193926 442350
rect 193982 442294 194078 442350
rect 193458 442226 194078 442294
rect 193458 442170 193554 442226
rect 193610 442170 193678 442226
rect 193734 442170 193802 442226
rect 193858 442170 193926 442226
rect 193982 442170 194078 442226
rect 193458 442102 194078 442170
rect 193458 442046 193554 442102
rect 193610 442046 193678 442102
rect 193734 442046 193802 442102
rect 193858 442046 193926 442102
rect 193982 442046 194078 442102
rect 193458 441978 194078 442046
rect 193458 441922 193554 441978
rect 193610 441922 193678 441978
rect 193734 441922 193802 441978
rect 193858 441922 193926 441978
rect 193982 441922 194078 441978
rect 193458 424350 194078 441922
rect 193458 424294 193554 424350
rect 193610 424294 193678 424350
rect 193734 424294 193802 424350
rect 193858 424294 193926 424350
rect 193982 424294 194078 424350
rect 193458 424226 194078 424294
rect 193458 424170 193554 424226
rect 193610 424170 193678 424226
rect 193734 424170 193802 424226
rect 193858 424170 193926 424226
rect 193982 424170 194078 424226
rect 193458 424102 194078 424170
rect 193458 424046 193554 424102
rect 193610 424046 193678 424102
rect 193734 424046 193802 424102
rect 193858 424046 193926 424102
rect 193982 424046 194078 424102
rect 193458 423978 194078 424046
rect 193458 423922 193554 423978
rect 193610 423922 193678 423978
rect 193734 423922 193802 423978
rect 193858 423922 193926 423978
rect 193982 423922 194078 423978
rect 193458 406350 194078 423922
rect 193458 406294 193554 406350
rect 193610 406294 193678 406350
rect 193734 406294 193802 406350
rect 193858 406294 193926 406350
rect 193982 406294 194078 406350
rect 193458 406226 194078 406294
rect 193458 406170 193554 406226
rect 193610 406170 193678 406226
rect 193734 406170 193802 406226
rect 193858 406170 193926 406226
rect 193982 406170 194078 406226
rect 193458 406102 194078 406170
rect 193458 406046 193554 406102
rect 193610 406046 193678 406102
rect 193734 406046 193802 406102
rect 193858 406046 193926 406102
rect 193982 406046 194078 406102
rect 193458 405978 194078 406046
rect 193458 405922 193554 405978
rect 193610 405922 193678 405978
rect 193734 405922 193802 405978
rect 193858 405922 193926 405978
rect 193982 405922 194078 405978
rect 193458 388350 194078 405922
rect 193458 388294 193554 388350
rect 193610 388294 193678 388350
rect 193734 388294 193802 388350
rect 193858 388294 193926 388350
rect 193982 388294 194078 388350
rect 193458 388226 194078 388294
rect 193458 388170 193554 388226
rect 193610 388170 193678 388226
rect 193734 388170 193802 388226
rect 193858 388170 193926 388226
rect 193982 388170 194078 388226
rect 193458 388102 194078 388170
rect 193458 388046 193554 388102
rect 193610 388046 193678 388102
rect 193734 388046 193802 388102
rect 193858 388046 193926 388102
rect 193982 388046 194078 388102
rect 193458 387978 194078 388046
rect 193458 387922 193554 387978
rect 193610 387922 193678 387978
rect 193734 387922 193802 387978
rect 193858 387922 193926 387978
rect 193982 387922 194078 387978
rect 193458 370350 194078 387922
rect 193458 370294 193554 370350
rect 193610 370294 193678 370350
rect 193734 370294 193802 370350
rect 193858 370294 193926 370350
rect 193982 370294 194078 370350
rect 193458 370226 194078 370294
rect 193458 370170 193554 370226
rect 193610 370170 193678 370226
rect 193734 370170 193802 370226
rect 193858 370170 193926 370226
rect 193982 370170 194078 370226
rect 193458 370102 194078 370170
rect 193458 370046 193554 370102
rect 193610 370046 193678 370102
rect 193734 370046 193802 370102
rect 193858 370046 193926 370102
rect 193982 370046 194078 370102
rect 193458 369978 194078 370046
rect 193458 369922 193554 369978
rect 193610 369922 193678 369978
rect 193734 369922 193802 369978
rect 193858 369922 193926 369978
rect 193982 369922 194078 369978
rect 193458 352350 194078 369922
rect 193458 352294 193554 352350
rect 193610 352294 193678 352350
rect 193734 352294 193802 352350
rect 193858 352294 193926 352350
rect 193982 352294 194078 352350
rect 193458 352226 194078 352294
rect 193458 352170 193554 352226
rect 193610 352170 193678 352226
rect 193734 352170 193802 352226
rect 193858 352170 193926 352226
rect 193982 352170 194078 352226
rect 193458 352102 194078 352170
rect 193458 352046 193554 352102
rect 193610 352046 193678 352102
rect 193734 352046 193802 352102
rect 193858 352046 193926 352102
rect 193982 352046 194078 352102
rect 193458 351978 194078 352046
rect 193458 351922 193554 351978
rect 193610 351922 193678 351978
rect 193734 351922 193802 351978
rect 193858 351922 193926 351978
rect 193982 351922 194078 351978
rect 193458 334350 194078 351922
rect 193458 334294 193554 334350
rect 193610 334294 193678 334350
rect 193734 334294 193802 334350
rect 193858 334294 193926 334350
rect 193982 334294 194078 334350
rect 193458 334226 194078 334294
rect 193458 334170 193554 334226
rect 193610 334170 193678 334226
rect 193734 334170 193802 334226
rect 193858 334170 193926 334226
rect 193982 334170 194078 334226
rect 193458 334102 194078 334170
rect 193458 334046 193554 334102
rect 193610 334046 193678 334102
rect 193734 334046 193802 334102
rect 193858 334046 193926 334102
rect 193982 334046 194078 334102
rect 193458 333978 194078 334046
rect 193458 333922 193554 333978
rect 193610 333922 193678 333978
rect 193734 333922 193802 333978
rect 193858 333922 193926 333978
rect 193982 333922 194078 333978
rect 193458 316350 194078 333922
rect 193458 316294 193554 316350
rect 193610 316294 193678 316350
rect 193734 316294 193802 316350
rect 193858 316294 193926 316350
rect 193982 316294 194078 316350
rect 193458 316226 194078 316294
rect 193458 316170 193554 316226
rect 193610 316170 193678 316226
rect 193734 316170 193802 316226
rect 193858 316170 193926 316226
rect 193982 316170 194078 316226
rect 193458 316102 194078 316170
rect 193458 316046 193554 316102
rect 193610 316046 193678 316102
rect 193734 316046 193802 316102
rect 193858 316046 193926 316102
rect 193982 316046 194078 316102
rect 193458 315978 194078 316046
rect 193458 315922 193554 315978
rect 193610 315922 193678 315978
rect 193734 315922 193802 315978
rect 193858 315922 193926 315978
rect 193982 315922 194078 315978
rect 193458 298350 194078 315922
rect 193458 298294 193554 298350
rect 193610 298294 193678 298350
rect 193734 298294 193802 298350
rect 193858 298294 193926 298350
rect 193982 298294 194078 298350
rect 193458 298226 194078 298294
rect 193458 298170 193554 298226
rect 193610 298170 193678 298226
rect 193734 298170 193802 298226
rect 193858 298170 193926 298226
rect 193982 298170 194078 298226
rect 193458 298102 194078 298170
rect 193458 298046 193554 298102
rect 193610 298046 193678 298102
rect 193734 298046 193802 298102
rect 193858 298046 193926 298102
rect 193982 298046 194078 298102
rect 193458 297978 194078 298046
rect 193458 297922 193554 297978
rect 193610 297922 193678 297978
rect 193734 297922 193802 297978
rect 193858 297922 193926 297978
rect 193982 297922 194078 297978
rect 193458 280350 194078 297922
rect 193458 280294 193554 280350
rect 193610 280294 193678 280350
rect 193734 280294 193802 280350
rect 193858 280294 193926 280350
rect 193982 280294 194078 280350
rect 193458 280226 194078 280294
rect 193458 280170 193554 280226
rect 193610 280170 193678 280226
rect 193734 280170 193802 280226
rect 193858 280170 193926 280226
rect 193982 280170 194078 280226
rect 193458 280102 194078 280170
rect 193458 280046 193554 280102
rect 193610 280046 193678 280102
rect 193734 280046 193802 280102
rect 193858 280046 193926 280102
rect 193982 280046 194078 280102
rect 193458 279978 194078 280046
rect 193458 279922 193554 279978
rect 193610 279922 193678 279978
rect 193734 279922 193802 279978
rect 193858 279922 193926 279978
rect 193982 279922 194078 279978
rect 193458 262350 194078 279922
rect 193458 262294 193554 262350
rect 193610 262294 193678 262350
rect 193734 262294 193802 262350
rect 193858 262294 193926 262350
rect 193982 262294 194078 262350
rect 193458 262226 194078 262294
rect 193458 262170 193554 262226
rect 193610 262170 193678 262226
rect 193734 262170 193802 262226
rect 193858 262170 193926 262226
rect 193982 262170 194078 262226
rect 193458 262102 194078 262170
rect 193458 262046 193554 262102
rect 193610 262046 193678 262102
rect 193734 262046 193802 262102
rect 193858 262046 193926 262102
rect 193982 262046 194078 262102
rect 193458 261978 194078 262046
rect 193458 261922 193554 261978
rect 193610 261922 193678 261978
rect 193734 261922 193802 261978
rect 193858 261922 193926 261978
rect 193982 261922 194078 261978
rect 193458 244350 194078 261922
rect 193458 244294 193554 244350
rect 193610 244294 193678 244350
rect 193734 244294 193802 244350
rect 193858 244294 193926 244350
rect 193982 244294 194078 244350
rect 193458 244226 194078 244294
rect 193458 244170 193554 244226
rect 193610 244170 193678 244226
rect 193734 244170 193802 244226
rect 193858 244170 193926 244226
rect 193982 244170 194078 244226
rect 193458 244102 194078 244170
rect 193458 244046 193554 244102
rect 193610 244046 193678 244102
rect 193734 244046 193802 244102
rect 193858 244046 193926 244102
rect 193982 244046 194078 244102
rect 193458 243978 194078 244046
rect 193458 243922 193554 243978
rect 193610 243922 193678 243978
rect 193734 243922 193802 243978
rect 193858 243922 193926 243978
rect 193982 243922 194078 243978
rect 193458 226350 194078 243922
rect 193458 226294 193554 226350
rect 193610 226294 193678 226350
rect 193734 226294 193802 226350
rect 193858 226294 193926 226350
rect 193982 226294 194078 226350
rect 193458 226226 194078 226294
rect 193458 226170 193554 226226
rect 193610 226170 193678 226226
rect 193734 226170 193802 226226
rect 193858 226170 193926 226226
rect 193982 226170 194078 226226
rect 193458 226102 194078 226170
rect 193458 226046 193554 226102
rect 193610 226046 193678 226102
rect 193734 226046 193802 226102
rect 193858 226046 193926 226102
rect 193982 226046 194078 226102
rect 193458 225978 194078 226046
rect 193458 225922 193554 225978
rect 193610 225922 193678 225978
rect 193734 225922 193802 225978
rect 193858 225922 193926 225978
rect 193982 225922 194078 225978
rect 193458 208350 194078 225922
rect 193458 208294 193554 208350
rect 193610 208294 193678 208350
rect 193734 208294 193802 208350
rect 193858 208294 193926 208350
rect 193982 208294 194078 208350
rect 193458 208226 194078 208294
rect 193458 208170 193554 208226
rect 193610 208170 193678 208226
rect 193734 208170 193802 208226
rect 193858 208170 193926 208226
rect 193982 208170 194078 208226
rect 193458 208102 194078 208170
rect 193458 208046 193554 208102
rect 193610 208046 193678 208102
rect 193734 208046 193802 208102
rect 193858 208046 193926 208102
rect 193982 208046 194078 208102
rect 193458 207978 194078 208046
rect 193458 207922 193554 207978
rect 193610 207922 193678 207978
rect 193734 207922 193802 207978
rect 193858 207922 193926 207978
rect 193982 207922 194078 207978
rect 193458 190350 194078 207922
rect 193458 190294 193554 190350
rect 193610 190294 193678 190350
rect 193734 190294 193802 190350
rect 193858 190294 193926 190350
rect 193982 190294 194078 190350
rect 193458 190226 194078 190294
rect 193458 190170 193554 190226
rect 193610 190170 193678 190226
rect 193734 190170 193802 190226
rect 193858 190170 193926 190226
rect 193982 190170 194078 190226
rect 193458 190102 194078 190170
rect 193458 190046 193554 190102
rect 193610 190046 193678 190102
rect 193734 190046 193802 190102
rect 193858 190046 193926 190102
rect 193982 190046 194078 190102
rect 193458 189978 194078 190046
rect 193458 189922 193554 189978
rect 193610 189922 193678 189978
rect 193734 189922 193802 189978
rect 193858 189922 193926 189978
rect 193982 189922 194078 189978
rect 193458 172350 194078 189922
rect 193458 172294 193554 172350
rect 193610 172294 193678 172350
rect 193734 172294 193802 172350
rect 193858 172294 193926 172350
rect 193982 172294 194078 172350
rect 193458 172226 194078 172294
rect 193458 172170 193554 172226
rect 193610 172170 193678 172226
rect 193734 172170 193802 172226
rect 193858 172170 193926 172226
rect 193982 172170 194078 172226
rect 193458 172102 194078 172170
rect 193458 172046 193554 172102
rect 193610 172046 193678 172102
rect 193734 172046 193802 172102
rect 193858 172046 193926 172102
rect 193982 172046 194078 172102
rect 193458 171978 194078 172046
rect 193458 171922 193554 171978
rect 193610 171922 193678 171978
rect 193734 171922 193802 171978
rect 193858 171922 193926 171978
rect 193982 171922 194078 171978
rect 193458 154350 194078 171922
rect 193458 154294 193554 154350
rect 193610 154294 193678 154350
rect 193734 154294 193802 154350
rect 193858 154294 193926 154350
rect 193982 154294 194078 154350
rect 193458 154226 194078 154294
rect 193458 154170 193554 154226
rect 193610 154170 193678 154226
rect 193734 154170 193802 154226
rect 193858 154170 193926 154226
rect 193982 154170 194078 154226
rect 193458 154102 194078 154170
rect 193458 154046 193554 154102
rect 193610 154046 193678 154102
rect 193734 154046 193802 154102
rect 193858 154046 193926 154102
rect 193982 154046 194078 154102
rect 193458 153978 194078 154046
rect 193458 153922 193554 153978
rect 193610 153922 193678 153978
rect 193734 153922 193802 153978
rect 193858 153922 193926 153978
rect 193982 153922 194078 153978
rect 193458 136350 194078 153922
rect 193458 136294 193554 136350
rect 193610 136294 193678 136350
rect 193734 136294 193802 136350
rect 193858 136294 193926 136350
rect 193982 136294 194078 136350
rect 193458 136226 194078 136294
rect 193458 136170 193554 136226
rect 193610 136170 193678 136226
rect 193734 136170 193802 136226
rect 193858 136170 193926 136226
rect 193982 136170 194078 136226
rect 193458 136102 194078 136170
rect 193458 136046 193554 136102
rect 193610 136046 193678 136102
rect 193734 136046 193802 136102
rect 193858 136046 193926 136102
rect 193982 136046 194078 136102
rect 193458 135978 194078 136046
rect 193458 135922 193554 135978
rect 193610 135922 193678 135978
rect 193734 135922 193802 135978
rect 193858 135922 193926 135978
rect 193982 135922 194078 135978
rect 193458 118350 194078 135922
rect 193458 118294 193554 118350
rect 193610 118294 193678 118350
rect 193734 118294 193802 118350
rect 193858 118294 193926 118350
rect 193982 118294 194078 118350
rect 193458 118226 194078 118294
rect 193458 118170 193554 118226
rect 193610 118170 193678 118226
rect 193734 118170 193802 118226
rect 193858 118170 193926 118226
rect 193982 118170 194078 118226
rect 193458 118102 194078 118170
rect 193458 118046 193554 118102
rect 193610 118046 193678 118102
rect 193734 118046 193802 118102
rect 193858 118046 193926 118102
rect 193982 118046 194078 118102
rect 193458 117978 194078 118046
rect 193458 117922 193554 117978
rect 193610 117922 193678 117978
rect 193734 117922 193802 117978
rect 193858 117922 193926 117978
rect 193982 117922 194078 117978
rect 193458 100350 194078 117922
rect 193458 100294 193554 100350
rect 193610 100294 193678 100350
rect 193734 100294 193802 100350
rect 193858 100294 193926 100350
rect 193982 100294 194078 100350
rect 193458 100226 194078 100294
rect 193458 100170 193554 100226
rect 193610 100170 193678 100226
rect 193734 100170 193802 100226
rect 193858 100170 193926 100226
rect 193982 100170 194078 100226
rect 193458 100102 194078 100170
rect 193458 100046 193554 100102
rect 193610 100046 193678 100102
rect 193734 100046 193802 100102
rect 193858 100046 193926 100102
rect 193982 100046 194078 100102
rect 193458 99978 194078 100046
rect 193458 99922 193554 99978
rect 193610 99922 193678 99978
rect 193734 99922 193802 99978
rect 193858 99922 193926 99978
rect 193982 99922 194078 99978
rect 193458 82350 194078 99922
rect 193458 82294 193554 82350
rect 193610 82294 193678 82350
rect 193734 82294 193802 82350
rect 193858 82294 193926 82350
rect 193982 82294 194078 82350
rect 193458 82226 194078 82294
rect 193458 82170 193554 82226
rect 193610 82170 193678 82226
rect 193734 82170 193802 82226
rect 193858 82170 193926 82226
rect 193982 82170 194078 82226
rect 193458 82102 194078 82170
rect 193458 82046 193554 82102
rect 193610 82046 193678 82102
rect 193734 82046 193802 82102
rect 193858 82046 193926 82102
rect 193982 82046 194078 82102
rect 193458 81978 194078 82046
rect 193458 81922 193554 81978
rect 193610 81922 193678 81978
rect 193734 81922 193802 81978
rect 193858 81922 193926 81978
rect 193982 81922 194078 81978
rect 193458 64350 194078 81922
rect 220458 597212 221078 598268
rect 220458 597156 220554 597212
rect 220610 597156 220678 597212
rect 220734 597156 220802 597212
rect 220858 597156 220926 597212
rect 220982 597156 221078 597212
rect 220458 597088 221078 597156
rect 220458 597032 220554 597088
rect 220610 597032 220678 597088
rect 220734 597032 220802 597088
rect 220858 597032 220926 597088
rect 220982 597032 221078 597088
rect 220458 596964 221078 597032
rect 220458 596908 220554 596964
rect 220610 596908 220678 596964
rect 220734 596908 220802 596964
rect 220858 596908 220926 596964
rect 220982 596908 221078 596964
rect 220458 596840 221078 596908
rect 220458 596784 220554 596840
rect 220610 596784 220678 596840
rect 220734 596784 220802 596840
rect 220858 596784 220926 596840
rect 220982 596784 221078 596840
rect 220458 580350 221078 596784
rect 220458 580294 220554 580350
rect 220610 580294 220678 580350
rect 220734 580294 220802 580350
rect 220858 580294 220926 580350
rect 220982 580294 221078 580350
rect 220458 580226 221078 580294
rect 220458 580170 220554 580226
rect 220610 580170 220678 580226
rect 220734 580170 220802 580226
rect 220858 580170 220926 580226
rect 220982 580170 221078 580226
rect 220458 580102 221078 580170
rect 220458 580046 220554 580102
rect 220610 580046 220678 580102
rect 220734 580046 220802 580102
rect 220858 580046 220926 580102
rect 220982 580046 221078 580102
rect 220458 579978 221078 580046
rect 220458 579922 220554 579978
rect 220610 579922 220678 579978
rect 220734 579922 220802 579978
rect 220858 579922 220926 579978
rect 220982 579922 221078 579978
rect 220458 562350 221078 579922
rect 220458 562294 220554 562350
rect 220610 562294 220678 562350
rect 220734 562294 220802 562350
rect 220858 562294 220926 562350
rect 220982 562294 221078 562350
rect 220458 562226 221078 562294
rect 220458 562170 220554 562226
rect 220610 562170 220678 562226
rect 220734 562170 220802 562226
rect 220858 562170 220926 562226
rect 220982 562170 221078 562226
rect 220458 562102 221078 562170
rect 220458 562046 220554 562102
rect 220610 562046 220678 562102
rect 220734 562046 220802 562102
rect 220858 562046 220926 562102
rect 220982 562046 221078 562102
rect 220458 561978 221078 562046
rect 220458 561922 220554 561978
rect 220610 561922 220678 561978
rect 220734 561922 220802 561978
rect 220858 561922 220926 561978
rect 220982 561922 221078 561978
rect 220458 544350 221078 561922
rect 220458 544294 220554 544350
rect 220610 544294 220678 544350
rect 220734 544294 220802 544350
rect 220858 544294 220926 544350
rect 220982 544294 221078 544350
rect 220458 544226 221078 544294
rect 220458 544170 220554 544226
rect 220610 544170 220678 544226
rect 220734 544170 220802 544226
rect 220858 544170 220926 544226
rect 220982 544170 221078 544226
rect 220458 544102 221078 544170
rect 220458 544046 220554 544102
rect 220610 544046 220678 544102
rect 220734 544046 220802 544102
rect 220858 544046 220926 544102
rect 220982 544046 221078 544102
rect 220458 543978 221078 544046
rect 220458 543922 220554 543978
rect 220610 543922 220678 543978
rect 220734 543922 220802 543978
rect 220858 543922 220926 543978
rect 220982 543922 221078 543978
rect 220458 526350 221078 543922
rect 220458 526294 220554 526350
rect 220610 526294 220678 526350
rect 220734 526294 220802 526350
rect 220858 526294 220926 526350
rect 220982 526294 221078 526350
rect 220458 526226 221078 526294
rect 220458 526170 220554 526226
rect 220610 526170 220678 526226
rect 220734 526170 220802 526226
rect 220858 526170 220926 526226
rect 220982 526170 221078 526226
rect 220458 526102 221078 526170
rect 220458 526046 220554 526102
rect 220610 526046 220678 526102
rect 220734 526046 220802 526102
rect 220858 526046 220926 526102
rect 220982 526046 221078 526102
rect 220458 525978 221078 526046
rect 220458 525922 220554 525978
rect 220610 525922 220678 525978
rect 220734 525922 220802 525978
rect 220858 525922 220926 525978
rect 220982 525922 221078 525978
rect 220458 508350 221078 525922
rect 220458 508294 220554 508350
rect 220610 508294 220678 508350
rect 220734 508294 220802 508350
rect 220858 508294 220926 508350
rect 220982 508294 221078 508350
rect 220458 508226 221078 508294
rect 220458 508170 220554 508226
rect 220610 508170 220678 508226
rect 220734 508170 220802 508226
rect 220858 508170 220926 508226
rect 220982 508170 221078 508226
rect 220458 508102 221078 508170
rect 220458 508046 220554 508102
rect 220610 508046 220678 508102
rect 220734 508046 220802 508102
rect 220858 508046 220926 508102
rect 220982 508046 221078 508102
rect 220458 507978 221078 508046
rect 220458 507922 220554 507978
rect 220610 507922 220678 507978
rect 220734 507922 220802 507978
rect 220858 507922 220926 507978
rect 220982 507922 221078 507978
rect 220458 490350 221078 507922
rect 220458 490294 220554 490350
rect 220610 490294 220678 490350
rect 220734 490294 220802 490350
rect 220858 490294 220926 490350
rect 220982 490294 221078 490350
rect 220458 490226 221078 490294
rect 220458 490170 220554 490226
rect 220610 490170 220678 490226
rect 220734 490170 220802 490226
rect 220858 490170 220926 490226
rect 220982 490170 221078 490226
rect 220458 490102 221078 490170
rect 220458 490046 220554 490102
rect 220610 490046 220678 490102
rect 220734 490046 220802 490102
rect 220858 490046 220926 490102
rect 220982 490046 221078 490102
rect 220458 489978 221078 490046
rect 220458 489922 220554 489978
rect 220610 489922 220678 489978
rect 220734 489922 220802 489978
rect 220858 489922 220926 489978
rect 220982 489922 221078 489978
rect 220458 472350 221078 489922
rect 220458 472294 220554 472350
rect 220610 472294 220678 472350
rect 220734 472294 220802 472350
rect 220858 472294 220926 472350
rect 220982 472294 221078 472350
rect 220458 472226 221078 472294
rect 220458 472170 220554 472226
rect 220610 472170 220678 472226
rect 220734 472170 220802 472226
rect 220858 472170 220926 472226
rect 220982 472170 221078 472226
rect 220458 472102 221078 472170
rect 220458 472046 220554 472102
rect 220610 472046 220678 472102
rect 220734 472046 220802 472102
rect 220858 472046 220926 472102
rect 220982 472046 221078 472102
rect 220458 471978 221078 472046
rect 220458 471922 220554 471978
rect 220610 471922 220678 471978
rect 220734 471922 220802 471978
rect 220858 471922 220926 471978
rect 220982 471922 221078 471978
rect 220458 454350 221078 471922
rect 220458 454294 220554 454350
rect 220610 454294 220678 454350
rect 220734 454294 220802 454350
rect 220858 454294 220926 454350
rect 220982 454294 221078 454350
rect 220458 454226 221078 454294
rect 220458 454170 220554 454226
rect 220610 454170 220678 454226
rect 220734 454170 220802 454226
rect 220858 454170 220926 454226
rect 220982 454170 221078 454226
rect 220458 454102 221078 454170
rect 220458 454046 220554 454102
rect 220610 454046 220678 454102
rect 220734 454046 220802 454102
rect 220858 454046 220926 454102
rect 220982 454046 221078 454102
rect 220458 453978 221078 454046
rect 220458 453922 220554 453978
rect 220610 453922 220678 453978
rect 220734 453922 220802 453978
rect 220858 453922 220926 453978
rect 220982 453922 221078 453978
rect 220458 436350 221078 453922
rect 220458 436294 220554 436350
rect 220610 436294 220678 436350
rect 220734 436294 220802 436350
rect 220858 436294 220926 436350
rect 220982 436294 221078 436350
rect 220458 436226 221078 436294
rect 220458 436170 220554 436226
rect 220610 436170 220678 436226
rect 220734 436170 220802 436226
rect 220858 436170 220926 436226
rect 220982 436170 221078 436226
rect 220458 436102 221078 436170
rect 220458 436046 220554 436102
rect 220610 436046 220678 436102
rect 220734 436046 220802 436102
rect 220858 436046 220926 436102
rect 220982 436046 221078 436102
rect 220458 435978 221078 436046
rect 220458 435922 220554 435978
rect 220610 435922 220678 435978
rect 220734 435922 220802 435978
rect 220858 435922 220926 435978
rect 220982 435922 221078 435978
rect 220458 418350 221078 435922
rect 220458 418294 220554 418350
rect 220610 418294 220678 418350
rect 220734 418294 220802 418350
rect 220858 418294 220926 418350
rect 220982 418294 221078 418350
rect 220458 418226 221078 418294
rect 220458 418170 220554 418226
rect 220610 418170 220678 418226
rect 220734 418170 220802 418226
rect 220858 418170 220926 418226
rect 220982 418170 221078 418226
rect 220458 418102 221078 418170
rect 220458 418046 220554 418102
rect 220610 418046 220678 418102
rect 220734 418046 220802 418102
rect 220858 418046 220926 418102
rect 220982 418046 221078 418102
rect 220458 417978 221078 418046
rect 220458 417922 220554 417978
rect 220610 417922 220678 417978
rect 220734 417922 220802 417978
rect 220858 417922 220926 417978
rect 220982 417922 221078 417978
rect 220458 400350 221078 417922
rect 220458 400294 220554 400350
rect 220610 400294 220678 400350
rect 220734 400294 220802 400350
rect 220858 400294 220926 400350
rect 220982 400294 221078 400350
rect 220458 400226 221078 400294
rect 220458 400170 220554 400226
rect 220610 400170 220678 400226
rect 220734 400170 220802 400226
rect 220858 400170 220926 400226
rect 220982 400170 221078 400226
rect 220458 400102 221078 400170
rect 220458 400046 220554 400102
rect 220610 400046 220678 400102
rect 220734 400046 220802 400102
rect 220858 400046 220926 400102
rect 220982 400046 221078 400102
rect 220458 399978 221078 400046
rect 220458 399922 220554 399978
rect 220610 399922 220678 399978
rect 220734 399922 220802 399978
rect 220858 399922 220926 399978
rect 220982 399922 221078 399978
rect 220458 382350 221078 399922
rect 220458 382294 220554 382350
rect 220610 382294 220678 382350
rect 220734 382294 220802 382350
rect 220858 382294 220926 382350
rect 220982 382294 221078 382350
rect 220458 382226 221078 382294
rect 220458 382170 220554 382226
rect 220610 382170 220678 382226
rect 220734 382170 220802 382226
rect 220858 382170 220926 382226
rect 220982 382170 221078 382226
rect 220458 382102 221078 382170
rect 220458 382046 220554 382102
rect 220610 382046 220678 382102
rect 220734 382046 220802 382102
rect 220858 382046 220926 382102
rect 220982 382046 221078 382102
rect 220458 381978 221078 382046
rect 220458 381922 220554 381978
rect 220610 381922 220678 381978
rect 220734 381922 220802 381978
rect 220858 381922 220926 381978
rect 220982 381922 221078 381978
rect 220458 364350 221078 381922
rect 220458 364294 220554 364350
rect 220610 364294 220678 364350
rect 220734 364294 220802 364350
rect 220858 364294 220926 364350
rect 220982 364294 221078 364350
rect 220458 364226 221078 364294
rect 220458 364170 220554 364226
rect 220610 364170 220678 364226
rect 220734 364170 220802 364226
rect 220858 364170 220926 364226
rect 220982 364170 221078 364226
rect 220458 364102 221078 364170
rect 220458 364046 220554 364102
rect 220610 364046 220678 364102
rect 220734 364046 220802 364102
rect 220858 364046 220926 364102
rect 220982 364046 221078 364102
rect 220458 363978 221078 364046
rect 220458 363922 220554 363978
rect 220610 363922 220678 363978
rect 220734 363922 220802 363978
rect 220858 363922 220926 363978
rect 220982 363922 221078 363978
rect 220458 346350 221078 363922
rect 220458 346294 220554 346350
rect 220610 346294 220678 346350
rect 220734 346294 220802 346350
rect 220858 346294 220926 346350
rect 220982 346294 221078 346350
rect 220458 346226 221078 346294
rect 220458 346170 220554 346226
rect 220610 346170 220678 346226
rect 220734 346170 220802 346226
rect 220858 346170 220926 346226
rect 220982 346170 221078 346226
rect 220458 346102 221078 346170
rect 220458 346046 220554 346102
rect 220610 346046 220678 346102
rect 220734 346046 220802 346102
rect 220858 346046 220926 346102
rect 220982 346046 221078 346102
rect 220458 345978 221078 346046
rect 220458 345922 220554 345978
rect 220610 345922 220678 345978
rect 220734 345922 220802 345978
rect 220858 345922 220926 345978
rect 220982 345922 221078 345978
rect 220458 328350 221078 345922
rect 220458 328294 220554 328350
rect 220610 328294 220678 328350
rect 220734 328294 220802 328350
rect 220858 328294 220926 328350
rect 220982 328294 221078 328350
rect 220458 328226 221078 328294
rect 220458 328170 220554 328226
rect 220610 328170 220678 328226
rect 220734 328170 220802 328226
rect 220858 328170 220926 328226
rect 220982 328170 221078 328226
rect 220458 328102 221078 328170
rect 220458 328046 220554 328102
rect 220610 328046 220678 328102
rect 220734 328046 220802 328102
rect 220858 328046 220926 328102
rect 220982 328046 221078 328102
rect 220458 327978 221078 328046
rect 220458 327922 220554 327978
rect 220610 327922 220678 327978
rect 220734 327922 220802 327978
rect 220858 327922 220926 327978
rect 220982 327922 221078 327978
rect 220458 310350 221078 327922
rect 220458 310294 220554 310350
rect 220610 310294 220678 310350
rect 220734 310294 220802 310350
rect 220858 310294 220926 310350
rect 220982 310294 221078 310350
rect 220458 310226 221078 310294
rect 220458 310170 220554 310226
rect 220610 310170 220678 310226
rect 220734 310170 220802 310226
rect 220858 310170 220926 310226
rect 220982 310170 221078 310226
rect 220458 310102 221078 310170
rect 220458 310046 220554 310102
rect 220610 310046 220678 310102
rect 220734 310046 220802 310102
rect 220858 310046 220926 310102
rect 220982 310046 221078 310102
rect 220458 309978 221078 310046
rect 220458 309922 220554 309978
rect 220610 309922 220678 309978
rect 220734 309922 220802 309978
rect 220858 309922 220926 309978
rect 220982 309922 221078 309978
rect 220458 292350 221078 309922
rect 220458 292294 220554 292350
rect 220610 292294 220678 292350
rect 220734 292294 220802 292350
rect 220858 292294 220926 292350
rect 220982 292294 221078 292350
rect 220458 292226 221078 292294
rect 220458 292170 220554 292226
rect 220610 292170 220678 292226
rect 220734 292170 220802 292226
rect 220858 292170 220926 292226
rect 220982 292170 221078 292226
rect 220458 292102 221078 292170
rect 220458 292046 220554 292102
rect 220610 292046 220678 292102
rect 220734 292046 220802 292102
rect 220858 292046 220926 292102
rect 220982 292046 221078 292102
rect 220458 291978 221078 292046
rect 220458 291922 220554 291978
rect 220610 291922 220678 291978
rect 220734 291922 220802 291978
rect 220858 291922 220926 291978
rect 220982 291922 221078 291978
rect 220458 274350 221078 291922
rect 220458 274294 220554 274350
rect 220610 274294 220678 274350
rect 220734 274294 220802 274350
rect 220858 274294 220926 274350
rect 220982 274294 221078 274350
rect 220458 274226 221078 274294
rect 220458 274170 220554 274226
rect 220610 274170 220678 274226
rect 220734 274170 220802 274226
rect 220858 274170 220926 274226
rect 220982 274170 221078 274226
rect 220458 274102 221078 274170
rect 220458 274046 220554 274102
rect 220610 274046 220678 274102
rect 220734 274046 220802 274102
rect 220858 274046 220926 274102
rect 220982 274046 221078 274102
rect 220458 273978 221078 274046
rect 220458 273922 220554 273978
rect 220610 273922 220678 273978
rect 220734 273922 220802 273978
rect 220858 273922 220926 273978
rect 220982 273922 221078 273978
rect 220458 256350 221078 273922
rect 220458 256294 220554 256350
rect 220610 256294 220678 256350
rect 220734 256294 220802 256350
rect 220858 256294 220926 256350
rect 220982 256294 221078 256350
rect 220458 256226 221078 256294
rect 220458 256170 220554 256226
rect 220610 256170 220678 256226
rect 220734 256170 220802 256226
rect 220858 256170 220926 256226
rect 220982 256170 221078 256226
rect 220458 256102 221078 256170
rect 220458 256046 220554 256102
rect 220610 256046 220678 256102
rect 220734 256046 220802 256102
rect 220858 256046 220926 256102
rect 220982 256046 221078 256102
rect 220458 255978 221078 256046
rect 220458 255922 220554 255978
rect 220610 255922 220678 255978
rect 220734 255922 220802 255978
rect 220858 255922 220926 255978
rect 220982 255922 221078 255978
rect 220458 238350 221078 255922
rect 220458 238294 220554 238350
rect 220610 238294 220678 238350
rect 220734 238294 220802 238350
rect 220858 238294 220926 238350
rect 220982 238294 221078 238350
rect 220458 238226 221078 238294
rect 220458 238170 220554 238226
rect 220610 238170 220678 238226
rect 220734 238170 220802 238226
rect 220858 238170 220926 238226
rect 220982 238170 221078 238226
rect 220458 238102 221078 238170
rect 220458 238046 220554 238102
rect 220610 238046 220678 238102
rect 220734 238046 220802 238102
rect 220858 238046 220926 238102
rect 220982 238046 221078 238102
rect 220458 237978 221078 238046
rect 220458 237922 220554 237978
rect 220610 237922 220678 237978
rect 220734 237922 220802 237978
rect 220858 237922 220926 237978
rect 220982 237922 221078 237978
rect 220458 220350 221078 237922
rect 220458 220294 220554 220350
rect 220610 220294 220678 220350
rect 220734 220294 220802 220350
rect 220858 220294 220926 220350
rect 220982 220294 221078 220350
rect 220458 220226 221078 220294
rect 220458 220170 220554 220226
rect 220610 220170 220678 220226
rect 220734 220170 220802 220226
rect 220858 220170 220926 220226
rect 220982 220170 221078 220226
rect 220458 220102 221078 220170
rect 220458 220046 220554 220102
rect 220610 220046 220678 220102
rect 220734 220046 220802 220102
rect 220858 220046 220926 220102
rect 220982 220046 221078 220102
rect 220458 219978 221078 220046
rect 220458 219922 220554 219978
rect 220610 219922 220678 219978
rect 220734 219922 220802 219978
rect 220858 219922 220926 219978
rect 220982 219922 221078 219978
rect 220458 202350 221078 219922
rect 220458 202294 220554 202350
rect 220610 202294 220678 202350
rect 220734 202294 220802 202350
rect 220858 202294 220926 202350
rect 220982 202294 221078 202350
rect 220458 202226 221078 202294
rect 220458 202170 220554 202226
rect 220610 202170 220678 202226
rect 220734 202170 220802 202226
rect 220858 202170 220926 202226
rect 220982 202170 221078 202226
rect 220458 202102 221078 202170
rect 220458 202046 220554 202102
rect 220610 202046 220678 202102
rect 220734 202046 220802 202102
rect 220858 202046 220926 202102
rect 220982 202046 221078 202102
rect 220458 201978 221078 202046
rect 220458 201922 220554 201978
rect 220610 201922 220678 201978
rect 220734 201922 220802 201978
rect 220858 201922 220926 201978
rect 220982 201922 221078 201978
rect 220458 184350 221078 201922
rect 220458 184294 220554 184350
rect 220610 184294 220678 184350
rect 220734 184294 220802 184350
rect 220858 184294 220926 184350
rect 220982 184294 221078 184350
rect 220458 184226 221078 184294
rect 220458 184170 220554 184226
rect 220610 184170 220678 184226
rect 220734 184170 220802 184226
rect 220858 184170 220926 184226
rect 220982 184170 221078 184226
rect 220458 184102 221078 184170
rect 220458 184046 220554 184102
rect 220610 184046 220678 184102
rect 220734 184046 220802 184102
rect 220858 184046 220926 184102
rect 220982 184046 221078 184102
rect 220458 183978 221078 184046
rect 220458 183922 220554 183978
rect 220610 183922 220678 183978
rect 220734 183922 220802 183978
rect 220858 183922 220926 183978
rect 220982 183922 221078 183978
rect 220458 166350 221078 183922
rect 220458 166294 220554 166350
rect 220610 166294 220678 166350
rect 220734 166294 220802 166350
rect 220858 166294 220926 166350
rect 220982 166294 221078 166350
rect 220458 166226 221078 166294
rect 220458 166170 220554 166226
rect 220610 166170 220678 166226
rect 220734 166170 220802 166226
rect 220858 166170 220926 166226
rect 220982 166170 221078 166226
rect 220458 166102 221078 166170
rect 220458 166046 220554 166102
rect 220610 166046 220678 166102
rect 220734 166046 220802 166102
rect 220858 166046 220926 166102
rect 220982 166046 221078 166102
rect 220458 165978 221078 166046
rect 220458 165922 220554 165978
rect 220610 165922 220678 165978
rect 220734 165922 220802 165978
rect 220858 165922 220926 165978
rect 220982 165922 221078 165978
rect 220458 148350 221078 165922
rect 220458 148294 220554 148350
rect 220610 148294 220678 148350
rect 220734 148294 220802 148350
rect 220858 148294 220926 148350
rect 220982 148294 221078 148350
rect 220458 148226 221078 148294
rect 220458 148170 220554 148226
rect 220610 148170 220678 148226
rect 220734 148170 220802 148226
rect 220858 148170 220926 148226
rect 220982 148170 221078 148226
rect 220458 148102 221078 148170
rect 220458 148046 220554 148102
rect 220610 148046 220678 148102
rect 220734 148046 220802 148102
rect 220858 148046 220926 148102
rect 220982 148046 221078 148102
rect 220458 147978 221078 148046
rect 220458 147922 220554 147978
rect 220610 147922 220678 147978
rect 220734 147922 220802 147978
rect 220858 147922 220926 147978
rect 220982 147922 221078 147978
rect 220458 130350 221078 147922
rect 220458 130294 220554 130350
rect 220610 130294 220678 130350
rect 220734 130294 220802 130350
rect 220858 130294 220926 130350
rect 220982 130294 221078 130350
rect 220458 130226 221078 130294
rect 220458 130170 220554 130226
rect 220610 130170 220678 130226
rect 220734 130170 220802 130226
rect 220858 130170 220926 130226
rect 220982 130170 221078 130226
rect 220458 130102 221078 130170
rect 220458 130046 220554 130102
rect 220610 130046 220678 130102
rect 220734 130046 220802 130102
rect 220858 130046 220926 130102
rect 220982 130046 221078 130102
rect 220458 129978 221078 130046
rect 220458 129922 220554 129978
rect 220610 129922 220678 129978
rect 220734 129922 220802 129978
rect 220858 129922 220926 129978
rect 220982 129922 221078 129978
rect 220458 112350 221078 129922
rect 220458 112294 220554 112350
rect 220610 112294 220678 112350
rect 220734 112294 220802 112350
rect 220858 112294 220926 112350
rect 220982 112294 221078 112350
rect 220458 112226 221078 112294
rect 220458 112170 220554 112226
rect 220610 112170 220678 112226
rect 220734 112170 220802 112226
rect 220858 112170 220926 112226
rect 220982 112170 221078 112226
rect 220458 112102 221078 112170
rect 220458 112046 220554 112102
rect 220610 112046 220678 112102
rect 220734 112046 220802 112102
rect 220858 112046 220926 112102
rect 220982 112046 221078 112102
rect 220458 111978 221078 112046
rect 220458 111922 220554 111978
rect 220610 111922 220678 111978
rect 220734 111922 220802 111978
rect 220858 111922 220926 111978
rect 220982 111922 221078 111978
rect 220458 94350 221078 111922
rect 220458 94294 220554 94350
rect 220610 94294 220678 94350
rect 220734 94294 220802 94350
rect 220858 94294 220926 94350
rect 220982 94294 221078 94350
rect 220458 94226 221078 94294
rect 220458 94170 220554 94226
rect 220610 94170 220678 94226
rect 220734 94170 220802 94226
rect 220858 94170 220926 94226
rect 220982 94170 221078 94226
rect 220458 94102 221078 94170
rect 220458 94046 220554 94102
rect 220610 94046 220678 94102
rect 220734 94046 220802 94102
rect 220858 94046 220926 94102
rect 220982 94046 221078 94102
rect 220458 93978 221078 94046
rect 220458 93922 220554 93978
rect 220610 93922 220678 93978
rect 220734 93922 220802 93978
rect 220858 93922 220926 93978
rect 220982 93922 221078 93978
rect 220458 76350 221078 93922
rect 220458 76294 220554 76350
rect 220610 76294 220678 76350
rect 220734 76294 220802 76350
rect 220858 76294 220926 76350
rect 220982 76294 221078 76350
rect 220458 76226 221078 76294
rect 220458 76170 220554 76226
rect 220610 76170 220678 76226
rect 220734 76170 220802 76226
rect 220858 76170 220926 76226
rect 220982 76170 221078 76226
rect 220458 76102 221078 76170
rect 220458 76046 220554 76102
rect 220610 76046 220678 76102
rect 220734 76046 220802 76102
rect 220858 76046 220926 76102
rect 220982 76046 221078 76102
rect 220458 75978 221078 76046
rect 220458 75922 220554 75978
rect 220610 75922 220678 75978
rect 220734 75922 220802 75978
rect 220858 75922 220926 75978
rect 220982 75922 221078 75978
rect 193458 64294 193554 64350
rect 193610 64294 193678 64350
rect 193734 64294 193802 64350
rect 193858 64294 193926 64350
rect 193982 64294 194078 64350
rect 193458 64226 194078 64294
rect 193458 64170 193554 64226
rect 193610 64170 193678 64226
rect 193734 64170 193802 64226
rect 193858 64170 193926 64226
rect 193982 64170 194078 64226
rect 193458 64102 194078 64170
rect 193458 64046 193554 64102
rect 193610 64046 193678 64102
rect 193734 64046 193802 64102
rect 193858 64046 193926 64102
rect 193982 64046 194078 64102
rect 193458 63978 194078 64046
rect 193458 63922 193554 63978
rect 193610 63922 193678 63978
rect 193734 63922 193802 63978
rect 193858 63922 193926 63978
rect 193982 63922 194078 63978
rect 193458 46350 194078 63922
rect 193458 46294 193554 46350
rect 193610 46294 193678 46350
rect 193734 46294 193802 46350
rect 193858 46294 193926 46350
rect 193982 46294 194078 46350
rect 193458 46226 194078 46294
rect 193458 46170 193554 46226
rect 193610 46170 193678 46226
rect 193734 46170 193802 46226
rect 193858 46170 193926 46226
rect 193982 46170 194078 46226
rect 193458 46102 194078 46170
rect 193458 46046 193554 46102
rect 193610 46046 193678 46102
rect 193734 46046 193802 46102
rect 193858 46046 193926 46102
rect 193982 46046 194078 46102
rect 193458 45978 194078 46046
rect 193458 45922 193554 45978
rect 193610 45922 193678 45978
rect 193734 45922 193802 45978
rect 193858 45922 193926 45978
rect 193982 45922 194078 45978
rect 189738 40294 189834 40350
rect 189890 40294 189958 40350
rect 190014 40294 190082 40350
rect 190138 40294 190206 40350
rect 190262 40294 190358 40350
rect 189738 40226 190358 40294
rect 189738 40170 189834 40226
rect 189890 40170 189958 40226
rect 190014 40170 190082 40226
rect 190138 40170 190206 40226
rect 190262 40170 190358 40226
rect 189738 40102 190358 40170
rect 189738 40046 189834 40102
rect 189890 40046 189958 40102
rect 190014 40046 190082 40102
rect 190138 40046 190206 40102
rect 190262 40046 190358 40102
rect 189738 39978 190358 40046
rect 189738 39922 189834 39978
rect 189890 39922 189958 39978
rect 190014 39922 190082 39978
rect 190138 39922 190206 39978
rect 190262 39922 190358 39978
rect 178108 32518 178164 32528
rect 173068 26938 173124 26948
rect 173068 20188 173124 26882
rect 174748 20638 174804 20648
rect 173068 20132 173236 20188
rect 166348 4162 166404 4172
rect 169372 8938 169428 8948
rect 169372 4228 169428 8882
rect 169372 4162 169428 4172
rect 173180 4228 173236 20132
rect 173180 4162 173236 4172
rect 174748 4228 174804 20582
rect 174748 4162 174804 4172
rect 178108 4228 178164 32462
rect 189738 22350 190358 39922
rect 189738 22294 189834 22350
rect 189890 22294 189958 22350
rect 190014 22294 190082 22350
rect 190138 22294 190206 22350
rect 190262 22294 190358 22350
rect 189738 22226 190358 22294
rect 189738 22170 189834 22226
rect 189890 22170 189958 22226
rect 190014 22170 190082 22226
rect 190138 22170 190206 22226
rect 190262 22170 190358 22226
rect 189738 22102 190358 22170
rect 189738 22046 189834 22102
rect 189890 22046 189958 22102
rect 190014 22046 190082 22102
rect 190138 22046 190206 22102
rect 190262 22046 190358 22102
rect 189738 21978 190358 22046
rect 189738 21922 189834 21978
rect 189890 21922 189958 21978
rect 190014 21922 190082 21978
rect 190138 21922 190206 21978
rect 190262 21922 190358 21978
rect 183148 17398 183204 17408
rect 178108 4162 178164 4172
rect 179788 13978 179844 13988
rect 179788 4228 179844 13922
rect 179788 4162 179844 4172
rect 183148 4228 183204 17342
rect 183148 4162 183204 4172
rect 189738 4350 190358 21922
rect 189738 4294 189834 4350
rect 189890 4294 189958 4350
rect 190014 4294 190082 4350
rect 190138 4294 190206 4350
rect 190262 4294 190358 4350
rect 189738 4226 190358 4294
rect 189738 4170 189834 4226
rect 189890 4170 189958 4226
rect 190014 4170 190082 4226
rect 190138 4170 190206 4226
rect 190262 4170 190358 4226
rect 162738 -1176 162834 -1120
rect 162890 -1176 162958 -1120
rect 163014 -1176 163082 -1120
rect 163138 -1176 163206 -1120
rect 163262 -1176 163358 -1120
rect 162738 -1244 163358 -1176
rect 162738 -1300 162834 -1244
rect 162890 -1300 162958 -1244
rect 163014 -1300 163082 -1244
rect 163138 -1300 163206 -1244
rect 163262 -1300 163358 -1244
rect 162738 -1368 163358 -1300
rect 162738 -1424 162834 -1368
rect 162890 -1424 162958 -1368
rect 163014 -1424 163082 -1368
rect 163138 -1424 163206 -1368
rect 163262 -1424 163358 -1368
rect 162738 -1492 163358 -1424
rect 162738 -1548 162834 -1492
rect 162890 -1548 162958 -1492
rect 163014 -1548 163082 -1492
rect 163138 -1548 163206 -1492
rect 163262 -1548 163358 -1492
rect 162738 -1644 163358 -1548
rect 189738 4102 190358 4170
rect 190428 45478 190484 45488
rect 190428 4228 190484 45422
rect 193458 28350 194078 45922
rect 193458 28294 193554 28350
rect 193610 28294 193678 28350
rect 193734 28294 193802 28350
rect 193858 28294 193926 28350
rect 193982 28294 194078 28350
rect 193458 28226 194078 28294
rect 193458 28170 193554 28226
rect 193610 28170 193678 28226
rect 193734 28170 193802 28226
rect 193858 28170 193926 28226
rect 193982 28170 194078 28226
rect 193458 28102 194078 28170
rect 193458 28046 193554 28102
rect 193610 28046 193678 28102
rect 193734 28046 193802 28102
rect 193858 28046 193926 28102
rect 193982 28046 194078 28102
rect 193458 27978 194078 28046
rect 193458 27922 193554 27978
rect 193610 27922 193678 27978
rect 193734 27922 193802 27978
rect 193858 27922 193926 27978
rect 193982 27922 194078 27978
rect 190428 4162 190484 4172
rect 191548 18838 191604 18848
rect 191548 4228 191604 18782
rect 191548 4162 191604 4172
rect 193458 10350 194078 27922
rect 206668 71398 206724 71408
rect 193458 10294 193554 10350
rect 193610 10294 193678 10350
rect 193734 10294 193802 10350
rect 193858 10294 193926 10350
rect 193982 10294 194078 10350
rect 193458 10226 194078 10294
rect 193458 10170 193554 10226
rect 193610 10170 193678 10226
rect 193734 10170 193802 10226
rect 193858 10170 193926 10226
rect 193982 10170 194078 10226
rect 193458 10102 194078 10170
rect 193458 10046 193554 10102
rect 193610 10046 193678 10102
rect 193734 10046 193802 10102
rect 193858 10046 193926 10102
rect 193982 10046 194078 10102
rect 193458 9978 194078 10046
rect 193458 9922 193554 9978
rect 193610 9922 193678 9978
rect 193734 9922 193802 9978
rect 193858 9922 193926 9978
rect 193982 9922 194078 9978
rect 189738 4046 189834 4102
rect 189890 4046 189958 4102
rect 190014 4046 190082 4102
rect 190138 4046 190206 4102
rect 190262 4046 190358 4102
rect 189738 3978 190358 4046
rect 189738 3922 189834 3978
rect 189890 3922 189958 3978
rect 190014 3922 190082 3978
rect 190138 3922 190206 3978
rect 190262 3922 190358 3978
rect 189738 -160 190358 3922
rect 193228 3538 193284 3548
rect 193228 3444 193284 3482
rect 193228 3378 193284 3388
rect 189738 -216 189834 -160
rect 189890 -216 189958 -160
rect 190014 -216 190082 -160
rect 190138 -216 190206 -160
rect 190262 -216 190358 -160
rect 189738 -284 190358 -216
rect 189738 -340 189834 -284
rect 189890 -340 189958 -284
rect 190014 -340 190082 -284
rect 190138 -340 190206 -284
rect 190262 -340 190358 -284
rect 189738 -408 190358 -340
rect 189738 -464 189834 -408
rect 189890 -464 189958 -408
rect 190014 -464 190082 -408
rect 190138 -464 190206 -408
rect 190262 -464 190358 -408
rect 189738 -532 190358 -464
rect 189738 -588 189834 -532
rect 189890 -588 189958 -532
rect 190014 -588 190082 -532
rect 190138 -588 190206 -532
rect 190262 -588 190358 -532
rect 189738 -1644 190358 -588
rect 193458 -1120 194078 9922
rect 194908 20458 194964 20468
rect 194908 4228 194964 20402
rect 194908 4162 194964 4172
rect 201740 15778 201796 15788
rect 201740 4228 201796 15722
rect 201740 4162 201796 4172
rect 203644 10918 203700 10928
rect 203644 4228 203700 10862
rect 203644 4162 203700 4172
rect 206668 4228 206724 71342
rect 216748 61138 216804 61148
rect 215068 37558 215124 37568
rect 206668 4162 206724 4172
rect 209356 7318 209412 7328
rect 209356 3668 209412 7262
rect 215068 4228 215124 37502
rect 216748 20188 216804 61082
rect 220458 58350 221078 75922
rect 224178 598172 224798 598268
rect 224178 598116 224274 598172
rect 224330 598116 224398 598172
rect 224454 598116 224522 598172
rect 224578 598116 224646 598172
rect 224702 598116 224798 598172
rect 224178 598048 224798 598116
rect 224178 597992 224274 598048
rect 224330 597992 224398 598048
rect 224454 597992 224522 598048
rect 224578 597992 224646 598048
rect 224702 597992 224798 598048
rect 224178 597924 224798 597992
rect 224178 597868 224274 597924
rect 224330 597868 224398 597924
rect 224454 597868 224522 597924
rect 224578 597868 224646 597924
rect 224702 597868 224798 597924
rect 224178 597800 224798 597868
rect 224178 597744 224274 597800
rect 224330 597744 224398 597800
rect 224454 597744 224522 597800
rect 224578 597744 224646 597800
rect 224702 597744 224798 597800
rect 224178 586350 224798 597744
rect 224178 586294 224274 586350
rect 224330 586294 224398 586350
rect 224454 586294 224522 586350
rect 224578 586294 224646 586350
rect 224702 586294 224798 586350
rect 224178 586226 224798 586294
rect 224178 586170 224274 586226
rect 224330 586170 224398 586226
rect 224454 586170 224522 586226
rect 224578 586170 224646 586226
rect 224702 586170 224798 586226
rect 224178 586102 224798 586170
rect 224178 586046 224274 586102
rect 224330 586046 224398 586102
rect 224454 586046 224522 586102
rect 224578 586046 224646 586102
rect 224702 586046 224798 586102
rect 224178 585978 224798 586046
rect 224178 585922 224274 585978
rect 224330 585922 224398 585978
rect 224454 585922 224522 585978
rect 224578 585922 224646 585978
rect 224702 585922 224798 585978
rect 224178 568350 224798 585922
rect 224178 568294 224274 568350
rect 224330 568294 224398 568350
rect 224454 568294 224522 568350
rect 224578 568294 224646 568350
rect 224702 568294 224798 568350
rect 224178 568226 224798 568294
rect 224178 568170 224274 568226
rect 224330 568170 224398 568226
rect 224454 568170 224522 568226
rect 224578 568170 224646 568226
rect 224702 568170 224798 568226
rect 224178 568102 224798 568170
rect 224178 568046 224274 568102
rect 224330 568046 224398 568102
rect 224454 568046 224522 568102
rect 224578 568046 224646 568102
rect 224702 568046 224798 568102
rect 224178 567978 224798 568046
rect 224178 567922 224274 567978
rect 224330 567922 224398 567978
rect 224454 567922 224522 567978
rect 224578 567922 224646 567978
rect 224702 567922 224798 567978
rect 224178 550350 224798 567922
rect 224178 550294 224274 550350
rect 224330 550294 224398 550350
rect 224454 550294 224522 550350
rect 224578 550294 224646 550350
rect 224702 550294 224798 550350
rect 224178 550226 224798 550294
rect 224178 550170 224274 550226
rect 224330 550170 224398 550226
rect 224454 550170 224522 550226
rect 224578 550170 224646 550226
rect 224702 550170 224798 550226
rect 224178 550102 224798 550170
rect 224178 550046 224274 550102
rect 224330 550046 224398 550102
rect 224454 550046 224522 550102
rect 224578 550046 224646 550102
rect 224702 550046 224798 550102
rect 224178 549978 224798 550046
rect 224178 549922 224274 549978
rect 224330 549922 224398 549978
rect 224454 549922 224522 549978
rect 224578 549922 224646 549978
rect 224702 549922 224798 549978
rect 224178 532350 224798 549922
rect 224178 532294 224274 532350
rect 224330 532294 224398 532350
rect 224454 532294 224522 532350
rect 224578 532294 224646 532350
rect 224702 532294 224798 532350
rect 224178 532226 224798 532294
rect 224178 532170 224274 532226
rect 224330 532170 224398 532226
rect 224454 532170 224522 532226
rect 224578 532170 224646 532226
rect 224702 532170 224798 532226
rect 224178 532102 224798 532170
rect 224178 532046 224274 532102
rect 224330 532046 224398 532102
rect 224454 532046 224522 532102
rect 224578 532046 224646 532102
rect 224702 532046 224798 532102
rect 224178 531978 224798 532046
rect 224178 531922 224274 531978
rect 224330 531922 224398 531978
rect 224454 531922 224522 531978
rect 224578 531922 224646 531978
rect 224702 531922 224798 531978
rect 224178 514350 224798 531922
rect 224178 514294 224274 514350
rect 224330 514294 224398 514350
rect 224454 514294 224522 514350
rect 224578 514294 224646 514350
rect 224702 514294 224798 514350
rect 224178 514226 224798 514294
rect 224178 514170 224274 514226
rect 224330 514170 224398 514226
rect 224454 514170 224522 514226
rect 224578 514170 224646 514226
rect 224702 514170 224798 514226
rect 224178 514102 224798 514170
rect 224178 514046 224274 514102
rect 224330 514046 224398 514102
rect 224454 514046 224522 514102
rect 224578 514046 224646 514102
rect 224702 514046 224798 514102
rect 224178 513978 224798 514046
rect 224178 513922 224274 513978
rect 224330 513922 224398 513978
rect 224454 513922 224522 513978
rect 224578 513922 224646 513978
rect 224702 513922 224798 513978
rect 224178 496350 224798 513922
rect 224178 496294 224274 496350
rect 224330 496294 224398 496350
rect 224454 496294 224522 496350
rect 224578 496294 224646 496350
rect 224702 496294 224798 496350
rect 224178 496226 224798 496294
rect 224178 496170 224274 496226
rect 224330 496170 224398 496226
rect 224454 496170 224522 496226
rect 224578 496170 224646 496226
rect 224702 496170 224798 496226
rect 224178 496102 224798 496170
rect 224178 496046 224274 496102
rect 224330 496046 224398 496102
rect 224454 496046 224522 496102
rect 224578 496046 224646 496102
rect 224702 496046 224798 496102
rect 224178 495978 224798 496046
rect 224178 495922 224274 495978
rect 224330 495922 224398 495978
rect 224454 495922 224522 495978
rect 224578 495922 224646 495978
rect 224702 495922 224798 495978
rect 224178 478350 224798 495922
rect 224178 478294 224274 478350
rect 224330 478294 224398 478350
rect 224454 478294 224522 478350
rect 224578 478294 224646 478350
rect 224702 478294 224798 478350
rect 224178 478226 224798 478294
rect 224178 478170 224274 478226
rect 224330 478170 224398 478226
rect 224454 478170 224522 478226
rect 224578 478170 224646 478226
rect 224702 478170 224798 478226
rect 224178 478102 224798 478170
rect 224178 478046 224274 478102
rect 224330 478046 224398 478102
rect 224454 478046 224522 478102
rect 224578 478046 224646 478102
rect 224702 478046 224798 478102
rect 224178 477978 224798 478046
rect 224178 477922 224274 477978
rect 224330 477922 224398 477978
rect 224454 477922 224522 477978
rect 224578 477922 224646 477978
rect 224702 477922 224798 477978
rect 224178 460350 224798 477922
rect 224178 460294 224274 460350
rect 224330 460294 224398 460350
rect 224454 460294 224522 460350
rect 224578 460294 224646 460350
rect 224702 460294 224798 460350
rect 224178 460226 224798 460294
rect 224178 460170 224274 460226
rect 224330 460170 224398 460226
rect 224454 460170 224522 460226
rect 224578 460170 224646 460226
rect 224702 460170 224798 460226
rect 224178 460102 224798 460170
rect 224178 460046 224274 460102
rect 224330 460046 224398 460102
rect 224454 460046 224522 460102
rect 224578 460046 224646 460102
rect 224702 460046 224798 460102
rect 224178 459978 224798 460046
rect 224178 459922 224274 459978
rect 224330 459922 224398 459978
rect 224454 459922 224522 459978
rect 224578 459922 224646 459978
rect 224702 459922 224798 459978
rect 224178 442350 224798 459922
rect 224178 442294 224274 442350
rect 224330 442294 224398 442350
rect 224454 442294 224522 442350
rect 224578 442294 224646 442350
rect 224702 442294 224798 442350
rect 224178 442226 224798 442294
rect 224178 442170 224274 442226
rect 224330 442170 224398 442226
rect 224454 442170 224522 442226
rect 224578 442170 224646 442226
rect 224702 442170 224798 442226
rect 224178 442102 224798 442170
rect 224178 442046 224274 442102
rect 224330 442046 224398 442102
rect 224454 442046 224522 442102
rect 224578 442046 224646 442102
rect 224702 442046 224798 442102
rect 224178 441978 224798 442046
rect 224178 441922 224274 441978
rect 224330 441922 224398 441978
rect 224454 441922 224522 441978
rect 224578 441922 224646 441978
rect 224702 441922 224798 441978
rect 224178 424350 224798 441922
rect 224178 424294 224274 424350
rect 224330 424294 224398 424350
rect 224454 424294 224522 424350
rect 224578 424294 224646 424350
rect 224702 424294 224798 424350
rect 224178 424226 224798 424294
rect 224178 424170 224274 424226
rect 224330 424170 224398 424226
rect 224454 424170 224522 424226
rect 224578 424170 224646 424226
rect 224702 424170 224798 424226
rect 224178 424102 224798 424170
rect 224178 424046 224274 424102
rect 224330 424046 224398 424102
rect 224454 424046 224522 424102
rect 224578 424046 224646 424102
rect 224702 424046 224798 424102
rect 224178 423978 224798 424046
rect 224178 423922 224274 423978
rect 224330 423922 224398 423978
rect 224454 423922 224522 423978
rect 224578 423922 224646 423978
rect 224702 423922 224798 423978
rect 224178 406350 224798 423922
rect 224178 406294 224274 406350
rect 224330 406294 224398 406350
rect 224454 406294 224522 406350
rect 224578 406294 224646 406350
rect 224702 406294 224798 406350
rect 224178 406226 224798 406294
rect 224178 406170 224274 406226
rect 224330 406170 224398 406226
rect 224454 406170 224522 406226
rect 224578 406170 224646 406226
rect 224702 406170 224798 406226
rect 224178 406102 224798 406170
rect 224178 406046 224274 406102
rect 224330 406046 224398 406102
rect 224454 406046 224522 406102
rect 224578 406046 224646 406102
rect 224702 406046 224798 406102
rect 224178 405978 224798 406046
rect 224178 405922 224274 405978
rect 224330 405922 224398 405978
rect 224454 405922 224522 405978
rect 224578 405922 224646 405978
rect 224702 405922 224798 405978
rect 224178 388350 224798 405922
rect 224178 388294 224274 388350
rect 224330 388294 224398 388350
rect 224454 388294 224522 388350
rect 224578 388294 224646 388350
rect 224702 388294 224798 388350
rect 224178 388226 224798 388294
rect 224178 388170 224274 388226
rect 224330 388170 224398 388226
rect 224454 388170 224522 388226
rect 224578 388170 224646 388226
rect 224702 388170 224798 388226
rect 224178 388102 224798 388170
rect 224178 388046 224274 388102
rect 224330 388046 224398 388102
rect 224454 388046 224522 388102
rect 224578 388046 224646 388102
rect 224702 388046 224798 388102
rect 224178 387978 224798 388046
rect 224178 387922 224274 387978
rect 224330 387922 224398 387978
rect 224454 387922 224522 387978
rect 224578 387922 224646 387978
rect 224702 387922 224798 387978
rect 224178 370350 224798 387922
rect 224178 370294 224274 370350
rect 224330 370294 224398 370350
rect 224454 370294 224522 370350
rect 224578 370294 224646 370350
rect 224702 370294 224798 370350
rect 224178 370226 224798 370294
rect 224178 370170 224274 370226
rect 224330 370170 224398 370226
rect 224454 370170 224522 370226
rect 224578 370170 224646 370226
rect 224702 370170 224798 370226
rect 224178 370102 224798 370170
rect 224178 370046 224274 370102
rect 224330 370046 224398 370102
rect 224454 370046 224522 370102
rect 224578 370046 224646 370102
rect 224702 370046 224798 370102
rect 224178 369978 224798 370046
rect 224178 369922 224274 369978
rect 224330 369922 224398 369978
rect 224454 369922 224522 369978
rect 224578 369922 224646 369978
rect 224702 369922 224798 369978
rect 224178 352350 224798 369922
rect 224178 352294 224274 352350
rect 224330 352294 224398 352350
rect 224454 352294 224522 352350
rect 224578 352294 224646 352350
rect 224702 352294 224798 352350
rect 224178 352226 224798 352294
rect 224178 352170 224274 352226
rect 224330 352170 224398 352226
rect 224454 352170 224522 352226
rect 224578 352170 224646 352226
rect 224702 352170 224798 352226
rect 224178 352102 224798 352170
rect 224178 352046 224274 352102
rect 224330 352046 224398 352102
rect 224454 352046 224522 352102
rect 224578 352046 224646 352102
rect 224702 352046 224798 352102
rect 224178 351978 224798 352046
rect 224178 351922 224274 351978
rect 224330 351922 224398 351978
rect 224454 351922 224522 351978
rect 224578 351922 224646 351978
rect 224702 351922 224798 351978
rect 224178 334350 224798 351922
rect 224178 334294 224274 334350
rect 224330 334294 224398 334350
rect 224454 334294 224522 334350
rect 224578 334294 224646 334350
rect 224702 334294 224798 334350
rect 224178 334226 224798 334294
rect 224178 334170 224274 334226
rect 224330 334170 224398 334226
rect 224454 334170 224522 334226
rect 224578 334170 224646 334226
rect 224702 334170 224798 334226
rect 224178 334102 224798 334170
rect 224178 334046 224274 334102
rect 224330 334046 224398 334102
rect 224454 334046 224522 334102
rect 224578 334046 224646 334102
rect 224702 334046 224798 334102
rect 224178 333978 224798 334046
rect 224178 333922 224274 333978
rect 224330 333922 224398 333978
rect 224454 333922 224522 333978
rect 224578 333922 224646 333978
rect 224702 333922 224798 333978
rect 224178 316350 224798 333922
rect 224178 316294 224274 316350
rect 224330 316294 224398 316350
rect 224454 316294 224522 316350
rect 224578 316294 224646 316350
rect 224702 316294 224798 316350
rect 224178 316226 224798 316294
rect 224178 316170 224274 316226
rect 224330 316170 224398 316226
rect 224454 316170 224522 316226
rect 224578 316170 224646 316226
rect 224702 316170 224798 316226
rect 224178 316102 224798 316170
rect 224178 316046 224274 316102
rect 224330 316046 224398 316102
rect 224454 316046 224522 316102
rect 224578 316046 224646 316102
rect 224702 316046 224798 316102
rect 224178 315978 224798 316046
rect 224178 315922 224274 315978
rect 224330 315922 224398 315978
rect 224454 315922 224522 315978
rect 224578 315922 224646 315978
rect 224702 315922 224798 315978
rect 224178 298350 224798 315922
rect 224178 298294 224274 298350
rect 224330 298294 224398 298350
rect 224454 298294 224522 298350
rect 224578 298294 224646 298350
rect 224702 298294 224798 298350
rect 224178 298226 224798 298294
rect 224178 298170 224274 298226
rect 224330 298170 224398 298226
rect 224454 298170 224522 298226
rect 224578 298170 224646 298226
rect 224702 298170 224798 298226
rect 224178 298102 224798 298170
rect 224178 298046 224274 298102
rect 224330 298046 224398 298102
rect 224454 298046 224522 298102
rect 224578 298046 224646 298102
rect 224702 298046 224798 298102
rect 224178 297978 224798 298046
rect 224178 297922 224274 297978
rect 224330 297922 224398 297978
rect 224454 297922 224522 297978
rect 224578 297922 224646 297978
rect 224702 297922 224798 297978
rect 224178 280350 224798 297922
rect 224178 280294 224274 280350
rect 224330 280294 224398 280350
rect 224454 280294 224522 280350
rect 224578 280294 224646 280350
rect 224702 280294 224798 280350
rect 224178 280226 224798 280294
rect 224178 280170 224274 280226
rect 224330 280170 224398 280226
rect 224454 280170 224522 280226
rect 224578 280170 224646 280226
rect 224702 280170 224798 280226
rect 224178 280102 224798 280170
rect 224178 280046 224274 280102
rect 224330 280046 224398 280102
rect 224454 280046 224522 280102
rect 224578 280046 224646 280102
rect 224702 280046 224798 280102
rect 224178 279978 224798 280046
rect 224178 279922 224274 279978
rect 224330 279922 224398 279978
rect 224454 279922 224522 279978
rect 224578 279922 224646 279978
rect 224702 279922 224798 279978
rect 224178 262350 224798 279922
rect 224178 262294 224274 262350
rect 224330 262294 224398 262350
rect 224454 262294 224522 262350
rect 224578 262294 224646 262350
rect 224702 262294 224798 262350
rect 224178 262226 224798 262294
rect 224178 262170 224274 262226
rect 224330 262170 224398 262226
rect 224454 262170 224522 262226
rect 224578 262170 224646 262226
rect 224702 262170 224798 262226
rect 224178 262102 224798 262170
rect 224178 262046 224274 262102
rect 224330 262046 224398 262102
rect 224454 262046 224522 262102
rect 224578 262046 224646 262102
rect 224702 262046 224798 262102
rect 224178 261978 224798 262046
rect 224178 261922 224274 261978
rect 224330 261922 224398 261978
rect 224454 261922 224522 261978
rect 224578 261922 224646 261978
rect 224702 261922 224798 261978
rect 224178 244350 224798 261922
rect 224178 244294 224274 244350
rect 224330 244294 224398 244350
rect 224454 244294 224522 244350
rect 224578 244294 224646 244350
rect 224702 244294 224798 244350
rect 224178 244226 224798 244294
rect 224178 244170 224274 244226
rect 224330 244170 224398 244226
rect 224454 244170 224522 244226
rect 224578 244170 224646 244226
rect 224702 244170 224798 244226
rect 224178 244102 224798 244170
rect 224178 244046 224274 244102
rect 224330 244046 224398 244102
rect 224454 244046 224522 244102
rect 224578 244046 224646 244102
rect 224702 244046 224798 244102
rect 224178 243978 224798 244046
rect 224178 243922 224274 243978
rect 224330 243922 224398 243978
rect 224454 243922 224522 243978
rect 224578 243922 224646 243978
rect 224702 243922 224798 243978
rect 224178 226350 224798 243922
rect 224178 226294 224274 226350
rect 224330 226294 224398 226350
rect 224454 226294 224522 226350
rect 224578 226294 224646 226350
rect 224702 226294 224798 226350
rect 224178 226226 224798 226294
rect 224178 226170 224274 226226
rect 224330 226170 224398 226226
rect 224454 226170 224522 226226
rect 224578 226170 224646 226226
rect 224702 226170 224798 226226
rect 224178 226102 224798 226170
rect 224178 226046 224274 226102
rect 224330 226046 224398 226102
rect 224454 226046 224522 226102
rect 224578 226046 224646 226102
rect 224702 226046 224798 226102
rect 224178 225978 224798 226046
rect 224178 225922 224274 225978
rect 224330 225922 224398 225978
rect 224454 225922 224522 225978
rect 224578 225922 224646 225978
rect 224702 225922 224798 225978
rect 224178 208350 224798 225922
rect 224178 208294 224274 208350
rect 224330 208294 224398 208350
rect 224454 208294 224522 208350
rect 224578 208294 224646 208350
rect 224702 208294 224798 208350
rect 224178 208226 224798 208294
rect 224178 208170 224274 208226
rect 224330 208170 224398 208226
rect 224454 208170 224522 208226
rect 224578 208170 224646 208226
rect 224702 208170 224798 208226
rect 224178 208102 224798 208170
rect 224178 208046 224274 208102
rect 224330 208046 224398 208102
rect 224454 208046 224522 208102
rect 224578 208046 224646 208102
rect 224702 208046 224798 208102
rect 224178 207978 224798 208046
rect 224178 207922 224274 207978
rect 224330 207922 224398 207978
rect 224454 207922 224522 207978
rect 224578 207922 224646 207978
rect 224702 207922 224798 207978
rect 224178 190350 224798 207922
rect 224178 190294 224274 190350
rect 224330 190294 224398 190350
rect 224454 190294 224522 190350
rect 224578 190294 224646 190350
rect 224702 190294 224798 190350
rect 224178 190226 224798 190294
rect 224178 190170 224274 190226
rect 224330 190170 224398 190226
rect 224454 190170 224522 190226
rect 224578 190170 224646 190226
rect 224702 190170 224798 190226
rect 224178 190102 224798 190170
rect 224178 190046 224274 190102
rect 224330 190046 224398 190102
rect 224454 190046 224522 190102
rect 224578 190046 224646 190102
rect 224702 190046 224798 190102
rect 224178 189978 224798 190046
rect 224178 189922 224274 189978
rect 224330 189922 224398 189978
rect 224454 189922 224522 189978
rect 224578 189922 224646 189978
rect 224702 189922 224798 189978
rect 224178 172350 224798 189922
rect 224178 172294 224274 172350
rect 224330 172294 224398 172350
rect 224454 172294 224522 172350
rect 224578 172294 224646 172350
rect 224702 172294 224798 172350
rect 224178 172226 224798 172294
rect 224178 172170 224274 172226
rect 224330 172170 224398 172226
rect 224454 172170 224522 172226
rect 224578 172170 224646 172226
rect 224702 172170 224798 172226
rect 224178 172102 224798 172170
rect 224178 172046 224274 172102
rect 224330 172046 224398 172102
rect 224454 172046 224522 172102
rect 224578 172046 224646 172102
rect 224702 172046 224798 172102
rect 224178 171978 224798 172046
rect 224178 171922 224274 171978
rect 224330 171922 224398 171978
rect 224454 171922 224522 171978
rect 224578 171922 224646 171978
rect 224702 171922 224798 171978
rect 224178 154350 224798 171922
rect 224178 154294 224274 154350
rect 224330 154294 224398 154350
rect 224454 154294 224522 154350
rect 224578 154294 224646 154350
rect 224702 154294 224798 154350
rect 224178 154226 224798 154294
rect 224178 154170 224274 154226
rect 224330 154170 224398 154226
rect 224454 154170 224522 154226
rect 224578 154170 224646 154226
rect 224702 154170 224798 154226
rect 224178 154102 224798 154170
rect 224178 154046 224274 154102
rect 224330 154046 224398 154102
rect 224454 154046 224522 154102
rect 224578 154046 224646 154102
rect 224702 154046 224798 154102
rect 224178 153978 224798 154046
rect 224178 153922 224274 153978
rect 224330 153922 224398 153978
rect 224454 153922 224522 153978
rect 224578 153922 224646 153978
rect 224702 153922 224798 153978
rect 224178 136350 224798 153922
rect 224178 136294 224274 136350
rect 224330 136294 224398 136350
rect 224454 136294 224522 136350
rect 224578 136294 224646 136350
rect 224702 136294 224798 136350
rect 224178 136226 224798 136294
rect 224178 136170 224274 136226
rect 224330 136170 224398 136226
rect 224454 136170 224522 136226
rect 224578 136170 224646 136226
rect 224702 136170 224798 136226
rect 224178 136102 224798 136170
rect 224178 136046 224274 136102
rect 224330 136046 224398 136102
rect 224454 136046 224522 136102
rect 224578 136046 224646 136102
rect 224702 136046 224798 136102
rect 224178 135978 224798 136046
rect 224178 135922 224274 135978
rect 224330 135922 224398 135978
rect 224454 135922 224522 135978
rect 224578 135922 224646 135978
rect 224702 135922 224798 135978
rect 224178 118350 224798 135922
rect 224178 118294 224274 118350
rect 224330 118294 224398 118350
rect 224454 118294 224522 118350
rect 224578 118294 224646 118350
rect 224702 118294 224798 118350
rect 224178 118226 224798 118294
rect 224178 118170 224274 118226
rect 224330 118170 224398 118226
rect 224454 118170 224522 118226
rect 224578 118170 224646 118226
rect 224702 118170 224798 118226
rect 224178 118102 224798 118170
rect 224178 118046 224274 118102
rect 224330 118046 224398 118102
rect 224454 118046 224522 118102
rect 224578 118046 224646 118102
rect 224702 118046 224798 118102
rect 224178 117978 224798 118046
rect 224178 117922 224274 117978
rect 224330 117922 224398 117978
rect 224454 117922 224522 117978
rect 224578 117922 224646 117978
rect 224702 117922 224798 117978
rect 224178 100350 224798 117922
rect 224178 100294 224274 100350
rect 224330 100294 224398 100350
rect 224454 100294 224522 100350
rect 224578 100294 224646 100350
rect 224702 100294 224798 100350
rect 224178 100226 224798 100294
rect 224178 100170 224274 100226
rect 224330 100170 224398 100226
rect 224454 100170 224522 100226
rect 224578 100170 224646 100226
rect 224702 100170 224798 100226
rect 224178 100102 224798 100170
rect 224178 100046 224274 100102
rect 224330 100046 224398 100102
rect 224454 100046 224522 100102
rect 224578 100046 224646 100102
rect 224702 100046 224798 100102
rect 224178 99978 224798 100046
rect 224178 99922 224274 99978
rect 224330 99922 224398 99978
rect 224454 99922 224522 99978
rect 224578 99922 224646 99978
rect 224702 99922 224798 99978
rect 224178 82350 224798 99922
rect 224178 82294 224274 82350
rect 224330 82294 224398 82350
rect 224454 82294 224522 82350
rect 224578 82294 224646 82350
rect 224702 82294 224798 82350
rect 224178 82226 224798 82294
rect 224178 82170 224274 82226
rect 224330 82170 224398 82226
rect 224454 82170 224522 82226
rect 224578 82170 224646 82226
rect 224702 82170 224798 82226
rect 224178 82102 224798 82170
rect 224178 82046 224274 82102
rect 224330 82046 224398 82102
rect 224454 82046 224522 82102
rect 224578 82046 224646 82102
rect 224702 82046 224798 82102
rect 224178 81978 224798 82046
rect 224178 81922 224274 81978
rect 224330 81922 224398 81978
rect 224454 81922 224522 81978
rect 224578 81922 224646 81978
rect 224702 81922 224798 81978
rect 220458 58294 220554 58350
rect 220610 58294 220678 58350
rect 220734 58294 220802 58350
rect 220858 58294 220926 58350
rect 220982 58294 221078 58350
rect 220458 58226 221078 58294
rect 220458 58170 220554 58226
rect 220610 58170 220678 58226
rect 220734 58170 220802 58226
rect 220858 58170 220926 58226
rect 220982 58170 221078 58226
rect 220458 58102 221078 58170
rect 220458 58046 220554 58102
rect 220610 58046 220678 58102
rect 220734 58046 220802 58102
rect 220858 58046 220926 58102
rect 220982 58046 221078 58102
rect 220458 57978 221078 58046
rect 220458 57922 220554 57978
rect 220610 57922 220678 57978
rect 220734 57922 220802 57978
rect 220858 57922 220926 57978
rect 220982 57922 221078 57978
rect 220108 40978 220164 40988
rect 216748 20132 217028 20188
rect 215068 4162 215124 4172
rect 216972 4228 217028 20132
rect 216972 4162 217028 4172
rect 220108 4228 220164 40922
rect 220108 4162 220164 4172
rect 220458 40350 221078 57922
rect 223468 67978 223524 67988
rect 220458 40294 220554 40350
rect 220610 40294 220678 40350
rect 220734 40294 220802 40350
rect 220858 40294 220926 40350
rect 220982 40294 221078 40350
rect 220458 40226 221078 40294
rect 220458 40170 220554 40226
rect 220610 40170 220678 40226
rect 220734 40170 220802 40226
rect 220858 40170 220926 40226
rect 220982 40170 221078 40226
rect 220458 40102 221078 40170
rect 220458 40046 220554 40102
rect 220610 40046 220678 40102
rect 220734 40046 220802 40102
rect 220858 40046 220926 40102
rect 220982 40046 221078 40102
rect 220458 39978 221078 40046
rect 220458 39922 220554 39978
rect 220610 39922 220678 39978
rect 220734 39922 220802 39978
rect 220858 39922 220926 39978
rect 220982 39922 221078 39978
rect 220458 22350 221078 39922
rect 220458 22294 220554 22350
rect 220610 22294 220678 22350
rect 220734 22294 220802 22350
rect 220858 22294 220926 22350
rect 220982 22294 221078 22350
rect 220458 22226 221078 22294
rect 220458 22170 220554 22226
rect 220610 22170 220678 22226
rect 220734 22170 220802 22226
rect 220858 22170 220926 22226
rect 220982 22170 221078 22226
rect 220458 22102 221078 22170
rect 220458 22046 220554 22102
rect 220610 22046 220678 22102
rect 220734 22046 220802 22102
rect 220858 22046 220926 22102
rect 220982 22046 221078 22102
rect 220458 21978 221078 22046
rect 220458 21922 220554 21978
rect 220610 21922 220678 21978
rect 220734 21922 220802 21978
rect 220858 21922 220926 21978
rect 220982 21922 221078 21978
rect 220458 4350 221078 21922
rect 220458 4294 220554 4350
rect 220610 4294 220678 4350
rect 220734 4294 220802 4350
rect 220858 4294 220926 4350
rect 220982 4294 221078 4350
rect 220458 4226 221078 4294
rect 220458 4170 220554 4226
rect 220610 4170 220678 4226
rect 220734 4170 220802 4226
rect 220858 4170 220926 4226
rect 220982 4170 221078 4226
rect 209356 3602 209412 3612
rect 220458 4102 221078 4170
rect 221788 47638 221844 47648
rect 221788 4228 221844 47582
rect 221788 4162 221844 4172
rect 223468 4228 223524 67922
rect 223468 4162 223524 4172
rect 224178 64350 224798 81922
rect 251178 597212 251798 598268
rect 251178 597156 251274 597212
rect 251330 597156 251398 597212
rect 251454 597156 251522 597212
rect 251578 597156 251646 597212
rect 251702 597156 251798 597212
rect 251178 597088 251798 597156
rect 251178 597032 251274 597088
rect 251330 597032 251398 597088
rect 251454 597032 251522 597088
rect 251578 597032 251646 597088
rect 251702 597032 251798 597088
rect 251178 596964 251798 597032
rect 251178 596908 251274 596964
rect 251330 596908 251398 596964
rect 251454 596908 251522 596964
rect 251578 596908 251646 596964
rect 251702 596908 251798 596964
rect 251178 596840 251798 596908
rect 251178 596784 251274 596840
rect 251330 596784 251398 596840
rect 251454 596784 251522 596840
rect 251578 596784 251646 596840
rect 251702 596784 251798 596840
rect 251178 580350 251798 596784
rect 251178 580294 251274 580350
rect 251330 580294 251398 580350
rect 251454 580294 251522 580350
rect 251578 580294 251646 580350
rect 251702 580294 251798 580350
rect 251178 580226 251798 580294
rect 251178 580170 251274 580226
rect 251330 580170 251398 580226
rect 251454 580170 251522 580226
rect 251578 580170 251646 580226
rect 251702 580170 251798 580226
rect 251178 580102 251798 580170
rect 251178 580046 251274 580102
rect 251330 580046 251398 580102
rect 251454 580046 251522 580102
rect 251578 580046 251646 580102
rect 251702 580046 251798 580102
rect 251178 579978 251798 580046
rect 251178 579922 251274 579978
rect 251330 579922 251398 579978
rect 251454 579922 251522 579978
rect 251578 579922 251646 579978
rect 251702 579922 251798 579978
rect 251178 562350 251798 579922
rect 251178 562294 251274 562350
rect 251330 562294 251398 562350
rect 251454 562294 251522 562350
rect 251578 562294 251646 562350
rect 251702 562294 251798 562350
rect 251178 562226 251798 562294
rect 251178 562170 251274 562226
rect 251330 562170 251398 562226
rect 251454 562170 251522 562226
rect 251578 562170 251646 562226
rect 251702 562170 251798 562226
rect 251178 562102 251798 562170
rect 251178 562046 251274 562102
rect 251330 562046 251398 562102
rect 251454 562046 251522 562102
rect 251578 562046 251646 562102
rect 251702 562046 251798 562102
rect 251178 561978 251798 562046
rect 251178 561922 251274 561978
rect 251330 561922 251398 561978
rect 251454 561922 251522 561978
rect 251578 561922 251646 561978
rect 251702 561922 251798 561978
rect 251178 544350 251798 561922
rect 251178 544294 251274 544350
rect 251330 544294 251398 544350
rect 251454 544294 251522 544350
rect 251578 544294 251646 544350
rect 251702 544294 251798 544350
rect 251178 544226 251798 544294
rect 251178 544170 251274 544226
rect 251330 544170 251398 544226
rect 251454 544170 251522 544226
rect 251578 544170 251646 544226
rect 251702 544170 251798 544226
rect 251178 544102 251798 544170
rect 251178 544046 251274 544102
rect 251330 544046 251398 544102
rect 251454 544046 251522 544102
rect 251578 544046 251646 544102
rect 251702 544046 251798 544102
rect 251178 543978 251798 544046
rect 251178 543922 251274 543978
rect 251330 543922 251398 543978
rect 251454 543922 251522 543978
rect 251578 543922 251646 543978
rect 251702 543922 251798 543978
rect 251178 526350 251798 543922
rect 251178 526294 251274 526350
rect 251330 526294 251398 526350
rect 251454 526294 251522 526350
rect 251578 526294 251646 526350
rect 251702 526294 251798 526350
rect 251178 526226 251798 526294
rect 251178 526170 251274 526226
rect 251330 526170 251398 526226
rect 251454 526170 251522 526226
rect 251578 526170 251646 526226
rect 251702 526170 251798 526226
rect 251178 526102 251798 526170
rect 251178 526046 251274 526102
rect 251330 526046 251398 526102
rect 251454 526046 251522 526102
rect 251578 526046 251646 526102
rect 251702 526046 251798 526102
rect 251178 525978 251798 526046
rect 251178 525922 251274 525978
rect 251330 525922 251398 525978
rect 251454 525922 251522 525978
rect 251578 525922 251646 525978
rect 251702 525922 251798 525978
rect 251178 508350 251798 525922
rect 251178 508294 251274 508350
rect 251330 508294 251398 508350
rect 251454 508294 251522 508350
rect 251578 508294 251646 508350
rect 251702 508294 251798 508350
rect 251178 508226 251798 508294
rect 251178 508170 251274 508226
rect 251330 508170 251398 508226
rect 251454 508170 251522 508226
rect 251578 508170 251646 508226
rect 251702 508170 251798 508226
rect 251178 508102 251798 508170
rect 251178 508046 251274 508102
rect 251330 508046 251398 508102
rect 251454 508046 251522 508102
rect 251578 508046 251646 508102
rect 251702 508046 251798 508102
rect 251178 507978 251798 508046
rect 251178 507922 251274 507978
rect 251330 507922 251398 507978
rect 251454 507922 251522 507978
rect 251578 507922 251646 507978
rect 251702 507922 251798 507978
rect 251178 490350 251798 507922
rect 251178 490294 251274 490350
rect 251330 490294 251398 490350
rect 251454 490294 251522 490350
rect 251578 490294 251646 490350
rect 251702 490294 251798 490350
rect 251178 490226 251798 490294
rect 251178 490170 251274 490226
rect 251330 490170 251398 490226
rect 251454 490170 251522 490226
rect 251578 490170 251646 490226
rect 251702 490170 251798 490226
rect 251178 490102 251798 490170
rect 251178 490046 251274 490102
rect 251330 490046 251398 490102
rect 251454 490046 251522 490102
rect 251578 490046 251646 490102
rect 251702 490046 251798 490102
rect 251178 489978 251798 490046
rect 251178 489922 251274 489978
rect 251330 489922 251398 489978
rect 251454 489922 251522 489978
rect 251578 489922 251646 489978
rect 251702 489922 251798 489978
rect 251178 472350 251798 489922
rect 251178 472294 251274 472350
rect 251330 472294 251398 472350
rect 251454 472294 251522 472350
rect 251578 472294 251646 472350
rect 251702 472294 251798 472350
rect 251178 472226 251798 472294
rect 251178 472170 251274 472226
rect 251330 472170 251398 472226
rect 251454 472170 251522 472226
rect 251578 472170 251646 472226
rect 251702 472170 251798 472226
rect 251178 472102 251798 472170
rect 251178 472046 251274 472102
rect 251330 472046 251398 472102
rect 251454 472046 251522 472102
rect 251578 472046 251646 472102
rect 251702 472046 251798 472102
rect 251178 471978 251798 472046
rect 251178 471922 251274 471978
rect 251330 471922 251398 471978
rect 251454 471922 251522 471978
rect 251578 471922 251646 471978
rect 251702 471922 251798 471978
rect 251178 454350 251798 471922
rect 251178 454294 251274 454350
rect 251330 454294 251398 454350
rect 251454 454294 251522 454350
rect 251578 454294 251646 454350
rect 251702 454294 251798 454350
rect 251178 454226 251798 454294
rect 251178 454170 251274 454226
rect 251330 454170 251398 454226
rect 251454 454170 251522 454226
rect 251578 454170 251646 454226
rect 251702 454170 251798 454226
rect 251178 454102 251798 454170
rect 251178 454046 251274 454102
rect 251330 454046 251398 454102
rect 251454 454046 251522 454102
rect 251578 454046 251646 454102
rect 251702 454046 251798 454102
rect 251178 453978 251798 454046
rect 251178 453922 251274 453978
rect 251330 453922 251398 453978
rect 251454 453922 251522 453978
rect 251578 453922 251646 453978
rect 251702 453922 251798 453978
rect 251178 436350 251798 453922
rect 251178 436294 251274 436350
rect 251330 436294 251398 436350
rect 251454 436294 251522 436350
rect 251578 436294 251646 436350
rect 251702 436294 251798 436350
rect 251178 436226 251798 436294
rect 251178 436170 251274 436226
rect 251330 436170 251398 436226
rect 251454 436170 251522 436226
rect 251578 436170 251646 436226
rect 251702 436170 251798 436226
rect 251178 436102 251798 436170
rect 251178 436046 251274 436102
rect 251330 436046 251398 436102
rect 251454 436046 251522 436102
rect 251578 436046 251646 436102
rect 251702 436046 251798 436102
rect 251178 435978 251798 436046
rect 251178 435922 251274 435978
rect 251330 435922 251398 435978
rect 251454 435922 251522 435978
rect 251578 435922 251646 435978
rect 251702 435922 251798 435978
rect 251178 418350 251798 435922
rect 251178 418294 251274 418350
rect 251330 418294 251398 418350
rect 251454 418294 251522 418350
rect 251578 418294 251646 418350
rect 251702 418294 251798 418350
rect 251178 418226 251798 418294
rect 251178 418170 251274 418226
rect 251330 418170 251398 418226
rect 251454 418170 251522 418226
rect 251578 418170 251646 418226
rect 251702 418170 251798 418226
rect 251178 418102 251798 418170
rect 251178 418046 251274 418102
rect 251330 418046 251398 418102
rect 251454 418046 251522 418102
rect 251578 418046 251646 418102
rect 251702 418046 251798 418102
rect 251178 417978 251798 418046
rect 251178 417922 251274 417978
rect 251330 417922 251398 417978
rect 251454 417922 251522 417978
rect 251578 417922 251646 417978
rect 251702 417922 251798 417978
rect 251178 400350 251798 417922
rect 251178 400294 251274 400350
rect 251330 400294 251398 400350
rect 251454 400294 251522 400350
rect 251578 400294 251646 400350
rect 251702 400294 251798 400350
rect 251178 400226 251798 400294
rect 251178 400170 251274 400226
rect 251330 400170 251398 400226
rect 251454 400170 251522 400226
rect 251578 400170 251646 400226
rect 251702 400170 251798 400226
rect 251178 400102 251798 400170
rect 251178 400046 251274 400102
rect 251330 400046 251398 400102
rect 251454 400046 251522 400102
rect 251578 400046 251646 400102
rect 251702 400046 251798 400102
rect 251178 399978 251798 400046
rect 251178 399922 251274 399978
rect 251330 399922 251398 399978
rect 251454 399922 251522 399978
rect 251578 399922 251646 399978
rect 251702 399922 251798 399978
rect 251178 382350 251798 399922
rect 251178 382294 251274 382350
rect 251330 382294 251398 382350
rect 251454 382294 251522 382350
rect 251578 382294 251646 382350
rect 251702 382294 251798 382350
rect 251178 382226 251798 382294
rect 251178 382170 251274 382226
rect 251330 382170 251398 382226
rect 251454 382170 251522 382226
rect 251578 382170 251646 382226
rect 251702 382170 251798 382226
rect 251178 382102 251798 382170
rect 251178 382046 251274 382102
rect 251330 382046 251398 382102
rect 251454 382046 251522 382102
rect 251578 382046 251646 382102
rect 251702 382046 251798 382102
rect 251178 381978 251798 382046
rect 251178 381922 251274 381978
rect 251330 381922 251398 381978
rect 251454 381922 251522 381978
rect 251578 381922 251646 381978
rect 251702 381922 251798 381978
rect 251178 364350 251798 381922
rect 251178 364294 251274 364350
rect 251330 364294 251398 364350
rect 251454 364294 251522 364350
rect 251578 364294 251646 364350
rect 251702 364294 251798 364350
rect 251178 364226 251798 364294
rect 251178 364170 251274 364226
rect 251330 364170 251398 364226
rect 251454 364170 251522 364226
rect 251578 364170 251646 364226
rect 251702 364170 251798 364226
rect 251178 364102 251798 364170
rect 251178 364046 251274 364102
rect 251330 364046 251398 364102
rect 251454 364046 251522 364102
rect 251578 364046 251646 364102
rect 251702 364046 251798 364102
rect 251178 363978 251798 364046
rect 251178 363922 251274 363978
rect 251330 363922 251398 363978
rect 251454 363922 251522 363978
rect 251578 363922 251646 363978
rect 251702 363922 251798 363978
rect 251178 346350 251798 363922
rect 251178 346294 251274 346350
rect 251330 346294 251398 346350
rect 251454 346294 251522 346350
rect 251578 346294 251646 346350
rect 251702 346294 251798 346350
rect 251178 346226 251798 346294
rect 251178 346170 251274 346226
rect 251330 346170 251398 346226
rect 251454 346170 251522 346226
rect 251578 346170 251646 346226
rect 251702 346170 251798 346226
rect 251178 346102 251798 346170
rect 251178 346046 251274 346102
rect 251330 346046 251398 346102
rect 251454 346046 251522 346102
rect 251578 346046 251646 346102
rect 251702 346046 251798 346102
rect 251178 345978 251798 346046
rect 251178 345922 251274 345978
rect 251330 345922 251398 345978
rect 251454 345922 251522 345978
rect 251578 345922 251646 345978
rect 251702 345922 251798 345978
rect 251178 328350 251798 345922
rect 251178 328294 251274 328350
rect 251330 328294 251398 328350
rect 251454 328294 251522 328350
rect 251578 328294 251646 328350
rect 251702 328294 251798 328350
rect 251178 328226 251798 328294
rect 251178 328170 251274 328226
rect 251330 328170 251398 328226
rect 251454 328170 251522 328226
rect 251578 328170 251646 328226
rect 251702 328170 251798 328226
rect 251178 328102 251798 328170
rect 251178 328046 251274 328102
rect 251330 328046 251398 328102
rect 251454 328046 251522 328102
rect 251578 328046 251646 328102
rect 251702 328046 251798 328102
rect 251178 327978 251798 328046
rect 251178 327922 251274 327978
rect 251330 327922 251398 327978
rect 251454 327922 251522 327978
rect 251578 327922 251646 327978
rect 251702 327922 251798 327978
rect 251178 310350 251798 327922
rect 251178 310294 251274 310350
rect 251330 310294 251398 310350
rect 251454 310294 251522 310350
rect 251578 310294 251646 310350
rect 251702 310294 251798 310350
rect 251178 310226 251798 310294
rect 251178 310170 251274 310226
rect 251330 310170 251398 310226
rect 251454 310170 251522 310226
rect 251578 310170 251646 310226
rect 251702 310170 251798 310226
rect 251178 310102 251798 310170
rect 251178 310046 251274 310102
rect 251330 310046 251398 310102
rect 251454 310046 251522 310102
rect 251578 310046 251646 310102
rect 251702 310046 251798 310102
rect 251178 309978 251798 310046
rect 251178 309922 251274 309978
rect 251330 309922 251398 309978
rect 251454 309922 251522 309978
rect 251578 309922 251646 309978
rect 251702 309922 251798 309978
rect 251178 292350 251798 309922
rect 251178 292294 251274 292350
rect 251330 292294 251398 292350
rect 251454 292294 251522 292350
rect 251578 292294 251646 292350
rect 251702 292294 251798 292350
rect 251178 292226 251798 292294
rect 251178 292170 251274 292226
rect 251330 292170 251398 292226
rect 251454 292170 251522 292226
rect 251578 292170 251646 292226
rect 251702 292170 251798 292226
rect 251178 292102 251798 292170
rect 251178 292046 251274 292102
rect 251330 292046 251398 292102
rect 251454 292046 251522 292102
rect 251578 292046 251646 292102
rect 251702 292046 251798 292102
rect 251178 291978 251798 292046
rect 251178 291922 251274 291978
rect 251330 291922 251398 291978
rect 251454 291922 251522 291978
rect 251578 291922 251646 291978
rect 251702 291922 251798 291978
rect 251178 274350 251798 291922
rect 251178 274294 251274 274350
rect 251330 274294 251398 274350
rect 251454 274294 251522 274350
rect 251578 274294 251646 274350
rect 251702 274294 251798 274350
rect 251178 274226 251798 274294
rect 251178 274170 251274 274226
rect 251330 274170 251398 274226
rect 251454 274170 251522 274226
rect 251578 274170 251646 274226
rect 251702 274170 251798 274226
rect 251178 274102 251798 274170
rect 251178 274046 251274 274102
rect 251330 274046 251398 274102
rect 251454 274046 251522 274102
rect 251578 274046 251646 274102
rect 251702 274046 251798 274102
rect 251178 273978 251798 274046
rect 251178 273922 251274 273978
rect 251330 273922 251398 273978
rect 251454 273922 251522 273978
rect 251578 273922 251646 273978
rect 251702 273922 251798 273978
rect 251178 256350 251798 273922
rect 251178 256294 251274 256350
rect 251330 256294 251398 256350
rect 251454 256294 251522 256350
rect 251578 256294 251646 256350
rect 251702 256294 251798 256350
rect 251178 256226 251798 256294
rect 251178 256170 251274 256226
rect 251330 256170 251398 256226
rect 251454 256170 251522 256226
rect 251578 256170 251646 256226
rect 251702 256170 251798 256226
rect 251178 256102 251798 256170
rect 251178 256046 251274 256102
rect 251330 256046 251398 256102
rect 251454 256046 251522 256102
rect 251578 256046 251646 256102
rect 251702 256046 251798 256102
rect 251178 255978 251798 256046
rect 251178 255922 251274 255978
rect 251330 255922 251398 255978
rect 251454 255922 251522 255978
rect 251578 255922 251646 255978
rect 251702 255922 251798 255978
rect 251178 238350 251798 255922
rect 251178 238294 251274 238350
rect 251330 238294 251398 238350
rect 251454 238294 251522 238350
rect 251578 238294 251646 238350
rect 251702 238294 251798 238350
rect 251178 238226 251798 238294
rect 251178 238170 251274 238226
rect 251330 238170 251398 238226
rect 251454 238170 251522 238226
rect 251578 238170 251646 238226
rect 251702 238170 251798 238226
rect 251178 238102 251798 238170
rect 251178 238046 251274 238102
rect 251330 238046 251398 238102
rect 251454 238046 251522 238102
rect 251578 238046 251646 238102
rect 251702 238046 251798 238102
rect 251178 237978 251798 238046
rect 251178 237922 251274 237978
rect 251330 237922 251398 237978
rect 251454 237922 251522 237978
rect 251578 237922 251646 237978
rect 251702 237922 251798 237978
rect 251178 220350 251798 237922
rect 251178 220294 251274 220350
rect 251330 220294 251398 220350
rect 251454 220294 251522 220350
rect 251578 220294 251646 220350
rect 251702 220294 251798 220350
rect 251178 220226 251798 220294
rect 251178 220170 251274 220226
rect 251330 220170 251398 220226
rect 251454 220170 251522 220226
rect 251578 220170 251646 220226
rect 251702 220170 251798 220226
rect 251178 220102 251798 220170
rect 251178 220046 251274 220102
rect 251330 220046 251398 220102
rect 251454 220046 251522 220102
rect 251578 220046 251646 220102
rect 251702 220046 251798 220102
rect 251178 219978 251798 220046
rect 251178 219922 251274 219978
rect 251330 219922 251398 219978
rect 251454 219922 251522 219978
rect 251578 219922 251646 219978
rect 251702 219922 251798 219978
rect 251178 202350 251798 219922
rect 251178 202294 251274 202350
rect 251330 202294 251398 202350
rect 251454 202294 251522 202350
rect 251578 202294 251646 202350
rect 251702 202294 251798 202350
rect 251178 202226 251798 202294
rect 251178 202170 251274 202226
rect 251330 202170 251398 202226
rect 251454 202170 251522 202226
rect 251578 202170 251646 202226
rect 251702 202170 251798 202226
rect 251178 202102 251798 202170
rect 251178 202046 251274 202102
rect 251330 202046 251398 202102
rect 251454 202046 251522 202102
rect 251578 202046 251646 202102
rect 251702 202046 251798 202102
rect 251178 201978 251798 202046
rect 251178 201922 251274 201978
rect 251330 201922 251398 201978
rect 251454 201922 251522 201978
rect 251578 201922 251646 201978
rect 251702 201922 251798 201978
rect 251178 184350 251798 201922
rect 251178 184294 251274 184350
rect 251330 184294 251398 184350
rect 251454 184294 251522 184350
rect 251578 184294 251646 184350
rect 251702 184294 251798 184350
rect 251178 184226 251798 184294
rect 251178 184170 251274 184226
rect 251330 184170 251398 184226
rect 251454 184170 251522 184226
rect 251578 184170 251646 184226
rect 251702 184170 251798 184226
rect 251178 184102 251798 184170
rect 251178 184046 251274 184102
rect 251330 184046 251398 184102
rect 251454 184046 251522 184102
rect 251578 184046 251646 184102
rect 251702 184046 251798 184102
rect 251178 183978 251798 184046
rect 251178 183922 251274 183978
rect 251330 183922 251398 183978
rect 251454 183922 251522 183978
rect 251578 183922 251646 183978
rect 251702 183922 251798 183978
rect 251178 166350 251798 183922
rect 251178 166294 251274 166350
rect 251330 166294 251398 166350
rect 251454 166294 251522 166350
rect 251578 166294 251646 166350
rect 251702 166294 251798 166350
rect 251178 166226 251798 166294
rect 251178 166170 251274 166226
rect 251330 166170 251398 166226
rect 251454 166170 251522 166226
rect 251578 166170 251646 166226
rect 251702 166170 251798 166226
rect 251178 166102 251798 166170
rect 251178 166046 251274 166102
rect 251330 166046 251398 166102
rect 251454 166046 251522 166102
rect 251578 166046 251646 166102
rect 251702 166046 251798 166102
rect 251178 165978 251798 166046
rect 251178 165922 251274 165978
rect 251330 165922 251398 165978
rect 251454 165922 251522 165978
rect 251578 165922 251646 165978
rect 251702 165922 251798 165978
rect 251178 148350 251798 165922
rect 251178 148294 251274 148350
rect 251330 148294 251398 148350
rect 251454 148294 251522 148350
rect 251578 148294 251646 148350
rect 251702 148294 251798 148350
rect 251178 148226 251798 148294
rect 251178 148170 251274 148226
rect 251330 148170 251398 148226
rect 251454 148170 251522 148226
rect 251578 148170 251646 148226
rect 251702 148170 251798 148226
rect 251178 148102 251798 148170
rect 251178 148046 251274 148102
rect 251330 148046 251398 148102
rect 251454 148046 251522 148102
rect 251578 148046 251646 148102
rect 251702 148046 251798 148102
rect 251178 147978 251798 148046
rect 251178 147922 251274 147978
rect 251330 147922 251398 147978
rect 251454 147922 251522 147978
rect 251578 147922 251646 147978
rect 251702 147922 251798 147978
rect 251178 130350 251798 147922
rect 251178 130294 251274 130350
rect 251330 130294 251398 130350
rect 251454 130294 251522 130350
rect 251578 130294 251646 130350
rect 251702 130294 251798 130350
rect 251178 130226 251798 130294
rect 251178 130170 251274 130226
rect 251330 130170 251398 130226
rect 251454 130170 251522 130226
rect 251578 130170 251646 130226
rect 251702 130170 251798 130226
rect 251178 130102 251798 130170
rect 251178 130046 251274 130102
rect 251330 130046 251398 130102
rect 251454 130046 251522 130102
rect 251578 130046 251646 130102
rect 251702 130046 251798 130102
rect 251178 129978 251798 130046
rect 251178 129922 251274 129978
rect 251330 129922 251398 129978
rect 251454 129922 251522 129978
rect 251578 129922 251646 129978
rect 251702 129922 251798 129978
rect 251178 112350 251798 129922
rect 251178 112294 251274 112350
rect 251330 112294 251398 112350
rect 251454 112294 251522 112350
rect 251578 112294 251646 112350
rect 251702 112294 251798 112350
rect 251178 112226 251798 112294
rect 251178 112170 251274 112226
rect 251330 112170 251398 112226
rect 251454 112170 251522 112226
rect 251578 112170 251646 112226
rect 251702 112170 251798 112226
rect 251178 112102 251798 112170
rect 251178 112046 251274 112102
rect 251330 112046 251398 112102
rect 251454 112046 251522 112102
rect 251578 112046 251646 112102
rect 251702 112046 251798 112102
rect 251178 111978 251798 112046
rect 251178 111922 251274 111978
rect 251330 111922 251398 111978
rect 251454 111922 251522 111978
rect 251578 111922 251646 111978
rect 251702 111922 251798 111978
rect 251178 94350 251798 111922
rect 251178 94294 251274 94350
rect 251330 94294 251398 94350
rect 251454 94294 251522 94350
rect 251578 94294 251646 94350
rect 251702 94294 251798 94350
rect 251178 94226 251798 94294
rect 251178 94170 251274 94226
rect 251330 94170 251398 94226
rect 251454 94170 251522 94226
rect 251578 94170 251646 94226
rect 251702 94170 251798 94226
rect 251178 94102 251798 94170
rect 251178 94046 251274 94102
rect 251330 94046 251398 94102
rect 251454 94046 251522 94102
rect 251578 94046 251646 94102
rect 251702 94046 251798 94102
rect 251178 93978 251798 94046
rect 251178 93922 251274 93978
rect 251330 93922 251398 93978
rect 251454 93922 251522 93978
rect 251578 93922 251646 93978
rect 251702 93922 251798 93978
rect 251178 76350 251798 93922
rect 251178 76294 251274 76350
rect 251330 76294 251398 76350
rect 251454 76294 251522 76350
rect 251578 76294 251646 76350
rect 251702 76294 251798 76350
rect 251178 76226 251798 76294
rect 251178 76170 251274 76226
rect 251330 76170 251398 76226
rect 251454 76170 251522 76226
rect 251578 76170 251646 76226
rect 251702 76170 251798 76226
rect 251178 76102 251798 76170
rect 251178 76046 251274 76102
rect 251330 76046 251398 76102
rect 251454 76046 251522 76102
rect 251578 76046 251646 76102
rect 251702 76046 251798 76102
rect 251178 75978 251798 76046
rect 251178 75922 251274 75978
rect 251330 75922 251398 75978
rect 251454 75922 251522 75978
rect 251578 75922 251646 75978
rect 251702 75922 251798 75978
rect 248668 71218 248724 71228
rect 238588 69418 238644 69428
rect 224178 64294 224274 64350
rect 224330 64294 224398 64350
rect 224454 64294 224522 64350
rect 224578 64294 224646 64350
rect 224702 64294 224798 64350
rect 224178 64226 224798 64294
rect 224178 64170 224274 64226
rect 224330 64170 224398 64226
rect 224454 64170 224522 64226
rect 224578 64170 224646 64226
rect 224702 64170 224798 64226
rect 224178 64102 224798 64170
rect 224178 64046 224274 64102
rect 224330 64046 224398 64102
rect 224454 64046 224522 64102
rect 224578 64046 224646 64102
rect 224702 64046 224798 64102
rect 224178 63978 224798 64046
rect 224178 63922 224274 63978
rect 224330 63922 224398 63978
rect 224454 63922 224522 63978
rect 224578 63922 224646 63978
rect 224702 63922 224798 63978
rect 224178 46350 224798 63922
rect 224178 46294 224274 46350
rect 224330 46294 224398 46350
rect 224454 46294 224522 46350
rect 224578 46294 224646 46350
rect 224702 46294 224798 46350
rect 224178 46226 224798 46294
rect 224178 46170 224274 46226
rect 224330 46170 224398 46226
rect 224454 46170 224522 46226
rect 224578 46170 224646 46226
rect 224702 46170 224798 46226
rect 224178 46102 224798 46170
rect 224178 46046 224274 46102
rect 224330 46046 224398 46102
rect 224454 46046 224522 46102
rect 224578 46046 224646 46102
rect 224702 46046 224798 46102
rect 224178 45978 224798 46046
rect 224178 45922 224274 45978
rect 224330 45922 224398 45978
rect 224454 45922 224522 45978
rect 224578 45922 224646 45978
rect 224702 45922 224798 45978
rect 224178 28350 224798 45922
rect 235228 66358 235284 66368
rect 231868 37378 231924 37388
rect 224178 28294 224274 28350
rect 224330 28294 224398 28350
rect 224454 28294 224522 28350
rect 224578 28294 224646 28350
rect 224702 28294 224798 28350
rect 224178 28226 224798 28294
rect 224178 28170 224274 28226
rect 224330 28170 224398 28226
rect 224454 28170 224522 28226
rect 224578 28170 224646 28226
rect 224702 28170 224798 28226
rect 224178 28102 224798 28170
rect 224178 28046 224274 28102
rect 224330 28046 224398 28102
rect 224454 28046 224522 28102
rect 224578 28046 224646 28102
rect 224702 28046 224798 28102
rect 224178 27978 224798 28046
rect 224178 27922 224274 27978
rect 224330 27922 224398 27978
rect 224454 27922 224522 27978
rect 224578 27922 224646 27978
rect 224702 27922 224798 27978
rect 224178 10350 224798 27922
rect 224178 10294 224274 10350
rect 224330 10294 224398 10350
rect 224454 10294 224522 10350
rect 224578 10294 224646 10350
rect 224702 10294 224798 10350
rect 224178 10226 224798 10294
rect 224178 10170 224274 10226
rect 224330 10170 224398 10226
rect 224454 10170 224522 10226
rect 224578 10170 224646 10226
rect 224702 10170 224798 10226
rect 224178 10102 224798 10170
rect 224178 10046 224274 10102
rect 224330 10046 224398 10102
rect 224454 10046 224522 10102
rect 224578 10046 224646 10102
rect 224702 10046 224798 10102
rect 224178 9978 224798 10046
rect 224178 9922 224274 9978
rect 224330 9922 224398 9978
rect 224454 9922 224522 9978
rect 224578 9922 224646 9978
rect 224702 9922 224798 9978
rect 220458 4046 220554 4102
rect 220610 4046 220678 4102
rect 220734 4046 220802 4102
rect 220858 4046 220926 4102
rect 220982 4046 221078 4102
rect 220458 3978 221078 4046
rect 220458 3922 220554 3978
rect 220610 3922 220678 3978
rect 220734 3922 220802 3978
rect 220858 3922 220926 3978
rect 220982 3922 221078 3978
rect 197932 2998 197988 3008
rect 197932 1988 197988 2942
rect 197932 1922 197988 1932
rect 211260 644 211316 654
rect 211260 118 211316 588
rect 211260 52 211316 62
rect 193458 -1176 193554 -1120
rect 193610 -1176 193678 -1120
rect 193734 -1176 193802 -1120
rect 193858 -1176 193926 -1120
rect 193982 -1176 194078 -1120
rect 193458 -1244 194078 -1176
rect 193458 -1300 193554 -1244
rect 193610 -1300 193678 -1244
rect 193734 -1300 193802 -1244
rect 193858 -1300 193926 -1244
rect 193982 -1300 194078 -1244
rect 193458 -1368 194078 -1300
rect 193458 -1424 193554 -1368
rect 193610 -1424 193678 -1368
rect 193734 -1424 193802 -1368
rect 193858 -1424 193926 -1368
rect 193982 -1424 194078 -1368
rect 193458 -1492 194078 -1424
rect 193458 -1548 193554 -1492
rect 193610 -1548 193678 -1492
rect 193734 -1548 193802 -1492
rect 193858 -1548 193926 -1492
rect 193982 -1548 194078 -1492
rect 193458 -1644 194078 -1548
rect 220458 -160 221078 3922
rect 220458 -216 220554 -160
rect 220610 -216 220678 -160
rect 220734 -216 220802 -160
rect 220858 -216 220926 -160
rect 220982 -216 221078 -160
rect 220458 -284 221078 -216
rect 220458 -340 220554 -284
rect 220610 -340 220678 -284
rect 220734 -340 220802 -284
rect 220858 -340 220926 -284
rect 220982 -340 221078 -284
rect 220458 -408 221078 -340
rect 220458 -464 220554 -408
rect 220610 -464 220678 -408
rect 220734 -464 220802 -408
rect 220858 -464 220926 -408
rect 220982 -464 221078 -408
rect 220458 -532 221078 -464
rect 220458 -588 220554 -532
rect 220610 -588 220678 -532
rect 220734 -588 220802 -532
rect 220858 -588 220926 -532
rect 220982 -588 221078 -532
rect 220458 -1644 221078 -588
rect 224178 -1120 224798 9922
rect 228508 36118 228564 36128
rect 228508 4228 228564 36062
rect 228508 4162 228564 4172
rect 231868 4228 231924 37322
rect 231868 4162 231924 4172
rect 233548 32338 233604 32348
rect 233548 4228 233604 32282
rect 233548 4162 233604 4172
rect 235228 4228 235284 66302
rect 235228 4162 235284 4172
rect 236908 25858 236964 25868
rect 236908 4228 236964 25802
rect 236908 4162 236964 4172
rect 238588 4228 238644 69362
rect 238588 4162 238644 4172
rect 243628 35938 243684 35948
rect 243628 4228 243684 35882
rect 243628 4162 243684 4172
rect 245532 18658 245588 18668
rect 245532 4228 245588 18602
rect 245532 4162 245588 4172
rect 248668 4228 248724 71162
rect 251178 58350 251798 75922
rect 254898 598172 255518 598268
rect 254898 598116 254994 598172
rect 255050 598116 255118 598172
rect 255174 598116 255242 598172
rect 255298 598116 255366 598172
rect 255422 598116 255518 598172
rect 254898 598048 255518 598116
rect 254898 597992 254994 598048
rect 255050 597992 255118 598048
rect 255174 597992 255242 598048
rect 255298 597992 255366 598048
rect 255422 597992 255518 598048
rect 254898 597924 255518 597992
rect 254898 597868 254994 597924
rect 255050 597868 255118 597924
rect 255174 597868 255242 597924
rect 255298 597868 255366 597924
rect 255422 597868 255518 597924
rect 254898 597800 255518 597868
rect 254898 597744 254994 597800
rect 255050 597744 255118 597800
rect 255174 597744 255242 597800
rect 255298 597744 255366 597800
rect 255422 597744 255518 597800
rect 254898 586350 255518 597744
rect 254898 586294 254994 586350
rect 255050 586294 255118 586350
rect 255174 586294 255242 586350
rect 255298 586294 255366 586350
rect 255422 586294 255518 586350
rect 254898 586226 255518 586294
rect 254898 586170 254994 586226
rect 255050 586170 255118 586226
rect 255174 586170 255242 586226
rect 255298 586170 255366 586226
rect 255422 586170 255518 586226
rect 254898 586102 255518 586170
rect 254898 586046 254994 586102
rect 255050 586046 255118 586102
rect 255174 586046 255242 586102
rect 255298 586046 255366 586102
rect 255422 586046 255518 586102
rect 254898 585978 255518 586046
rect 254898 585922 254994 585978
rect 255050 585922 255118 585978
rect 255174 585922 255242 585978
rect 255298 585922 255366 585978
rect 255422 585922 255518 585978
rect 254898 568350 255518 585922
rect 254898 568294 254994 568350
rect 255050 568294 255118 568350
rect 255174 568294 255242 568350
rect 255298 568294 255366 568350
rect 255422 568294 255518 568350
rect 254898 568226 255518 568294
rect 254898 568170 254994 568226
rect 255050 568170 255118 568226
rect 255174 568170 255242 568226
rect 255298 568170 255366 568226
rect 255422 568170 255518 568226
rect 254898 568102 255518 568170
rect 254898 568046 254994 568102
rect 255050 568046 255118 568102
rect 255174 568046 255242 568102
rect 255298 568046 255366 568102
rect 255422 568046 255518 568102
rect 254898 567978 255518 568046
rect 254898 567922 254994 567978
rect 255050 567922 255118 567978
rect 255174 567922 255242 567978
rect 255298 567922 255366 567978
rect 255422 567922 255518 567978
rect 254898 550350 255518 567922
rect 254898 550294 254994 550350
rect 255050 550294 255118 550350
rect 255174 550294 255242 550350
rect 255298 550294 255366 550350
rect 255422 550294 255518 550350
rect 254898 550226 255518 550294
rect 254898 550170 254994 550226
rect 255050 550170 255118 550226
rect 255174 550170 255242 550226
rect 255298 550170 255366 550226
rect 255422 550170 255518 550226
rect 254898 550102 255518 550170
rect 254898 550046 254994 550102
rect 255050 550046 255118 550102
rect 255174 550046 255242 550102
rect 255298 550046 255366 550102
rect 255422 550046 255518 550102
rect 254898 549978 255518 550046
rect 254898 549922 254994 549978
rect 255050 549922 255118 549978
rect 255174 549922 255242 549978
rect 255298 549922 255366 549978
rect 255422 549922 255518 549978
rect 254898 532350 255518 549922
rect 254898 532294 254994 532350
rect 255050 532294 255118 532350
rect 255174 532294 255242 532350
rect 255298 532294 255366 532350
rect 255422 532294 255518 532350
rect 254898 532226 255518 532294
rect 254898 532170 254994 532226
rect 255050 532170 255118 532226
rect 255174 532170 255242 532226
rect 255298 532170 255366 532226
rect 255422 532170 255518 532226
rect 254898 532102 255518 532170
rect 254898 532046 254994 532102
rect 255050 532046 255118 532102
rect 255174 532046 255242 532102
rect 255298 532046 255366 532102
rect 255422 532046 255518 532102
rect 254898 531978 255518 532046
rect 254898 531922 254994 531978
rect 255050 531922 255118 531978
rect 255174 531922 255242 531978
rect 255298 531922 255366 531978
rect 255422 531922 255518 531978
rect 254898 514350 255518 531922
rect 254898 514294 254994 514350
rect 255050 514294 255118 514350
rect 255174 514294 255242 514350
rect 255298 514294 255366 514350
rect 255422 514294 255518 514350
rect 254898 514226 255518 514294
rect 254898 514170 254994 514226
rect 255050 514170 255118 514226
rect 255174 514170 255242 514226
rect 255298 514170 255366 514226
rect 255422 514170 255518 514226
rect 254898 514102 255518 514170
rect 254898 514046 254994 514102
rect 255050 514046 255118 514102
rect 255174 514046 255242 514102
rect 255298 514046 255366 514102
rect 255422 514046 255518 514102
rect 254898 513978 255518 514046
rect 254898 513922 254994 513978
rect 255050 513922 255118 513978
rect 255174 513922 255242 513978
rect 255298 513922 255366 513978
rect 255422 513922 255518 513978
rect 254898 496350 255518 513922
rect 254898 496294 254994 496350
rect 255050 496294 255118 496350
rect 255174 496294 255242 496350
rect 255298 496294 255366 496350
rect 255422 496294 255518 496350
rect 254898 496226 255518 496294
rect 254898 496170 254994 496226
rect 255050 496170 255118 496226
rect 255174 496170 255242 496226
rect 255298 496170 255366 496226
rect 255422 496170 255518 496226
rect 254898 496102 255518 496170
rect 254898 496046 254994 496102
rect 255050 496046 255118 496102
rect 255174 496046 255242 496102
rect 255298 496046 255366 496102
rect 255422 496046 255518 496102
rect 254898 495978 255518 496046
rect 254898 495922 254994 495978
rect 255050 495922 255118 495978
rect 255174 495922 255242 495978
rect 255298 495922 255366 495978
rect 255422 495922 255518 495978
rect 254898 478350 255518 495922
rect 254898 478294 254994 478350
rect 255050 478294 255118 478350
rect 255174 478294 255242 478350
rect 255298 478294 255366 478350
rect 255422 478294 255518 478350
rect 254898 478226 255518 478294
rect 254898 478170 254994 478226
rect 255050 478170 255118 478226
rect 255174 478170 255242 478226
rect 255298 478170 255366 478226
rect 255422 478170 255518 478226
rect 254898 478102 255518 478170
rect 254898 478046 254994 478102
rect 255050 478046 255118 478102
rect 255174 478046 255242 478102
rect 255298 478046 255366 478102
rect 255422 478046 255518 478102
rect 254898 477978 255518 478046
rect 254898 477922 254994 477978
rect 255050 477922 255118 477978
rect 255174 477922 255242 477978
rect 255298 477922 255366 477978
rect 255422 477922 255518 477978
rect 254898 460350 255518 477922
rect 254898 460294 254994 460350
rect 255050 460294 255118 460350
rect 255174 460294 255242 460350
rect 255298 460294 255366 460350
rect 255422 460294 255518 460350
rect 254898 460226 255518 460294
rect 254898 460170 254994 460226
rect 255050 460170 255118 460226
rect 255174 460170 255242 460226
rect 255298 460170 255366 460226
rect 255422 460170 255518 460226
rect 254898 460102 255518 460170
rect 254898 460046 254994 460102
rect 255050 460046 255118 460102
rect 255174 460046 255242 460102
rect 255298 460046 255366 460102
rect 255422 460046 255518 460102
rect 254898 459978 255518 460046
rect 254898 459922 254994 459978
rect 255050 459922 255118 459978
rect 255174 459922 255242 459978
rect 255298 459922 255366 459978
rect 255422 459922 255518 459978
rect 254898 442350 255518 459922
rect 254898 442294 254994 442350
rect 255050 442294 255118 442350
rect 255174 442294 255242 442350
rect 255298 442294 255366 442350
rect 255422 442294 255518 442350
rect 254898 442226 255518 442294
rect 254898 442170 254994 442226
rect 255050 442170 255118 442226
rect 255174 442170 255242 442226
rect 255298 442170 255366 442226
rect 255422 442170 255518 442226
rect 254898 442102 255518 442170
rect 254898 442046 254994 442102
rect 255050 442046 255118 442102
rect 255174 442046 255242 442102
rect 255298 442046 255366 442102
rect 255422 442046 255518 442102
rect 254898 441978 255518 442046
rect 254898 441922 254994 441978
rect 255050 441922 255118 441978
rect 255174 441922 255242 441978
rect 255298 441922 255366 441978
rect 255422 441922 255518 441978
rect 254898 424350 255518 441922
rect 254898 424294 254994 424350
rect 255050 424294 255118 424350
rect 255174 424294 255242 424350
rect 255298 424294 255366 424350
rect 255422 424294 255518 424350
rect 254898 424226 255518 424294
rect 254898 424170 254994 424226
rect 255050 424170 255118 424226
rect 255174 424170 255242 424226
rect 255298 424170 255366 424226
rect 255422 424170 255518 424226
rect 254898 424102 255518 424170
rect 254898 424046 254994 424102
rect 255050 424046 255118 424102
rect 255174 424046 255242 424102
rect 255298 424046 255366 424102
rect 255422 424046 255518 424102
rect 254898 423978 255518 424046
rect 254898 423922 254994 423978
rect 255050 423922 255118 423978
rect 255174 423922 255242 423978
rect 255298 423922 255366 423978
rect 255422 423922 255518 423978
rect 254898 406350 255518 423922
rect 254898 406294 254994 406350
rect 255050 406294 255118 406350
rect 255174 406294 255242 406350
rect 255298 406294 255366 406350
rect 255422 406294 255518 406350
rect 254898 406226 255518 406294
rect 254898 406170 254994 406226
rect 255050 406170 255118 406226
rect 255174 406170 255242 406226
rect 255298 406170 255366 406226
rect 255422 406170 255518 406226
rect 254898 406102 255518 406170
rect 254898 406046 254994 406102
rect 255050 406046 255118 406102
rect 255174 406046 255242 406102
rect 255298 406046 255366 406102
rect 255422 406046 255518 406102
rect 254898 405978 255518 406046
rect 254898 405922 254994 405978
rect 255050 405922 255118 405978
rect 255174 405922 255242 405978
rect 255298 405922 255366 405978
rect 255422 405922 255518 405978
rect 254898 388350 255518 405922
rect 254898 388294 254994 388350
rect 255050 388294 255118 388350
rect 255174 388294 255242 388350
rect 255298 388294 255366 388350
rect 255422 388294 255518 388350
rect 254898 388226 255518 388294
rect 254898 388170 254994 388226
rect 255050 388170 255118 388226
rect 255174 388170 255242 388226
rect 255298 388170 255366 388226
rect 255422 388170 255518 388226
rect 254898 388102 255518 388170
rect 254898 388046 254994 388102
rect 255050 388046 255118 388102
rect 255174 388046 255242 388102
rect 255298 388046 255366 388102
rect 255422 388046 255518 388102
rect 254898 387978 255518 388046
rect 254898 387922 254994 387978
rect 255050 387922 255118 387978
rect 255174 387922 255242 387978
rect 255298 387922 255366 387978
rect 255422 387922 255518 387978
rect 254898 370350 255518 387922
rect 254898 370294 254994 370350
rect 255050 370294 255118 370350
rect 255174 370294 255242 370350
rect 255298 370294 255366 370350
rect 255422 370294 255518 370350
rect 254898 370226 255518 370294
rect 254898 370170 254994 370226
rect 255050 370170 255118 370226
rect 255174 370170 255242 370226
rect 255298 370170 255366 370226
rect 255422 370170 255518 370226
rect 254898 370102 255518 370170
rect 254898 370046 254994 370102
rect 255050 370046 255118 370102
rect 255174 370046 255242 370102
rect 255298 370046 255366 370102
rect 255422 370046 255518 370102
rect 254898 369978 255518 370046
rect 254898 369922 254994 369978
rect 255050 369922 255118 369978
rect 255174 369922 255242 369978
rect 255298 369922 255366 369978
rect 255422 369922 255518 369978
rect 254898 352350 255518 369922
rect 254898 352294 254994 352350
rect 255050 352294 255118 352350
rect 255174 352294 255242 352350
rect 255298 352294 255366 352350
rect 255422 352294 255518 352350
rect 254898 352226 255518 352294
rect 254898 352170 254994 352226
rect 255050 352170 255118 352226
rect 255174 352170 255242 352226
rect 255298 352170 255366 352226
rect 255422 352170 255518 352226
rect 254898 352102 255518 352170
rect 254898 352046 254994 352102
rect 255050 352046 255118 352102
rect 255174 352046 255242 352102
rect 255298 352046 255366 352102
rect 255422 352046 255518 352102
rect 254898 351978 255518 352046
rect 254898 351922 254994 351978
rect 255050 351922 255118 351978
rect 255174 351922 255242 351978
rect 255298 351922 255366 351978
rect 255422 351922 255518 351978
rect 254898 334350 255518 351922
rect 254898 334294 254994 334350
rect 255050 334294 255118 334350
rect 255174 334294 255242 334350
rect 255298 334294 255366 334350
rect 255422 334294 255518 334350
rect 254898 334226 255518 334294
rect 254898 334170 254994 334226
rect 255050 334170 255118 334226
rect 255174 334170 255242 334226
rect 255298 334170 255366 334226
rect 255422 334170 255518 334226
rect 254898 334102 255518 334170
rect 254898 334046 254994 334102
rect 255050 334046 255118 334102
rect 255174 334046 255242 334102
rect 255298 334046 255366 334102
rect 255422 334046 255518 334102
rect 254898 333978 255518 334046
rect 254898 333922 254994 333978
rect 255050 333922 255118 333978
rect 255174 333922 255242 333978
rect 255298 333922 255366 333978
rect 255422 333922 255518 333978
rect 254898 316350 255518 333922
rect 254898 316294 254994 316350
rect 255050 316294 255118 316350
rect 255174 316294 255242 316350
rect 255298 316294 255366 316350
rect 255422 316294 255518 316350
rect 254898 316226 255518 316294
rect 254898 316170 254994 316226
rect 255050 316170 255118 316226
rect 255174 316170 255242 316226
rect 255298 316170 255366 316226
rect 255422 316170 255518 316226
rect 254898 316102 255518 316170
rect 254898 316046 254994 316102
rect 255050 316046 255118 316102
rect 255174 316046 255242 316102
rect 255298 316046 255366 316102
rect 255422 316046 255518 316102
rect 254898 315978 255518 316046
rect 254898 315922 254994 315978
rect 255050 315922 255118 315978
rect 255174 315922 255242 315978
rect 255298 315922 255366 315978
rect 255422 315922 255518 315978
rect 254898 298350 255518 315922
rect 254898 298294 254994 298350
rect 255050 298294 255118 298350
rect 255174 298294 255242 298350
rect 255298 298294 255366 298350
rect 255422 298294 255518 298350
rect 254898 298226 255518 298294
rect 254898 298170 254994 298226
rect 255050 298170 255118 298226
rect 255174 298170 255242 298226
rect 255298 298170 255366 298226
rect 255422 298170 255518 298226
rect 254898 298102 255518 298170
rect 254898 298046 254994 298102
rect 255050 298046 255118 298102
rect 255174 298046 255242 298102
rect 255298 298046 255366 298102
rect 255422 298046 255518 298102
rect 254898 297978 255518 298046
rect 254898 297922 254994 297978
rect 255050 297922 255118 297978
rect 255174 297922 255242 297978
rect 255298 297922 255366 297978
rect 255422 297922 255518 297978
rect 254898 280350 255518 297922
rect 254898 280294 254994 280350
rect 255050 280294 255118 280350
rect 255174 280294 255242 280350
rect 255298 280294 255366 280350
rect 255422 280294 255518 280350
rect 254898 280226 255518 280294
rect 254898 280170 254994 280226
rect 255050 280170 255118 280226
rect 255174 280170 255242 280226
rect 255298 280170 255366 280226
rect 255422 280170 255518 280226
rect 254898 280102 255518 280170
rect 254898 280046 254994 280102
rect 255050 280046 255118 280102
rect 255174 280046 255242 280102
rect 255298 280046 255366 280102
rect 255422 280046 255518 280102
rect 254898 279978 255518 280046
rect 254898 279922 254994 279978
rect 255050 279922 255118 279978
rect 255174 279922 255242 279978
rect 255298 279922 255366 279978
rect 255422 279922 255518 279978
rect 254898 262350 255518 279922
rect 254898 262294 254994 262350
rect 255050 262294 255118 262350
rect 255174 262294 255242 262350
rect 255298 262294 255366 262350
rect 255422 262294 255518 262350
rect 254898 262226 255518 262294
rect 254898 262170 254994 262226
rect 255050 262170 255118 262226
rect 255174 262170 255242 262226
rect 255298 262170 255366 262226
rect 255422 262170 255518 262226
rect 254898 262102 255518 262170
rect 254898 262046 254994 262102
rect 255050 262046 255118 262102
rect 255174 262046 255242 262102
rect 255298 262046 255366 262102
rect 255422 262046 255518 262102
rect 254898 261978 255518 262046
rect 254898 261922 254994 261978
rect 255050 261922 255118 261978
rect 255174 261922 255242 261978
rect 255298 261922 255366 261978
rect 255422 261922 255518 261978
rect 254898 244350 255518 261922
rect 254898 244294 254994 244350
rect 255050 244294 255118 244350
rect 255174 244294 255242 244350
rect 255298 244294 255366 244350
rect 255422 244294 255518 244350
rect 254898 244226 255518 244294
rect 254898 244170 254994 244226
rect 255050 244170 255118 244226
rect 255174 244170 255242 244226
rect 255298 244170 255366 244226
rect 255422 244170 255518 244226
rect 254898 244102 255518 244170
rect 254898 244046 254994 244102
rect 255050 244046 255118 244102
rect 255174 244046 255242 244102
rect 255298 244046 255366 244102
rect 255422 244046 255518 244102
rect 254898 243978 255518 244046
rect 254898 243922 254994 243978
rect 255050 243922 255118 243978
rect 255174 243922 255242 243978
rect 255298 243922 255366 243978
rect 255422 243922 255518 243978
rect 254898 226350 255518 243922
rect 254898 226294 254994 226350
rect 255050 226294 255118 226350
rect 255174 226294 255242 226350
rect 255298 226294 255366 226350
rect 255422 226294 255518 226350
rect 254898 226226 255518 226294
rect 254898 226170 254994 226226
rect 255050 226170 255118 226226
rect 255174 226170 255242 226226
rect 255298 226170 255366 226226
rect 255422 226170 255518 226226
rect 254898 226102 255518 226170
rect 254898 226046 254994 226102
rect 255050 226046 255118 226102
rect 255174 226046 255242 226102
rect 255298 226046 255366 226102
rect 255422 226046 255518 226102
rect 254898 225978 255518 226046
rect 254898 225922 254994 225978
rect 255050 225922 255118 225978
rect 255174 225922 255242 225978
rect 255298 225922 255366 225978
rect 255422 225922 255518 225978
rect 254898 208350 255518 225922
rect 254898 208294 254994 208350
rect 255050 208294 255118 208350
rect 255174 208294 255242 208350
rect 255298 208294 255366 208350
rect 255422 208294 255518 208350
rect 254898 208226 255518 208294
rect 254898 208170 254994 208226
rect 255050 208170 255118 208226
rect 255174 208170 255242 208226
rect 255298 208170 255366 208226
rect 255422 208170 255518 208226
rect 254898 208102 255518 208170
rect 254898 208046 254994 208102
rect 255050 208046 255118 208102
rect 255174 208046 255242 208102
rect 255298 208046 255366 208102
rect 255422 208046 255518 208102
rect 254898 207978 255518 208046
rect 254898 207922 254994 207978
rect 255050 207922 255118 207978
rect 255174 207922 255242 207978
rect 255298 207922 255366 207978
rect 255422 207922 255518 207978
rect 254898 190350 255518 207922
rect 254898 190294 254994 190350
rect 255050 190294 255118 190350
rect 255174 190294 255242 190350
rect 255298 190294 255366 190350
rect 255422 190294 255518 190350
rect 254898 190226 255518 190294
rect 254898 190170 254994 190226
rect 255050 190170 255118 190226
rect 255174 190170 255242 190226
rect 255298 190170 255366 190226
rect 255422 190170 255518 190226
rect 254898 190102 255518 190170
rect 254898 190046 254994 190102
rect 255050 190046 255118 190102
rect 255174 190046 255242 190102
rect 255298 190046 255366 190102
rect 255422 190046 255518 190102
rect 254898 189978 255518 190046
rect 254898 189922 254994 189978
rect 255050 189922 255118 189978
rect 255174 189922 255242 189978
rect 255298 189922 255366 189978
rect 255422 189922 255518 189978
rect 254898 172350 255518 189922
rect 254898 172294 254994 172350
rect 255050 172294 255118 172350
rect 255174 172294 255242 172350
rect 255298 172294 255366 172350
rect 255422 172294 255518 172350
rect 254898 172226 255518 172294
rect 254898 172170 254994 172226
rect 255050 172170 255118 172226
rect 255174 172170 255242 172226
rect 255298 172170 255366 172226
rect 255422 172170 255518 172226
rect 254898 172102 255518 172170
rect 254898 172046 254994 172102
rect 255050 172046 255118 172102
rect 255174 172046 255242 172102
rect 255298 172046 255366 172102
rect 255422 172046 255518 172102
rect 254898 171978 255518 172046
rect 254898 171922 254994 171978
rect 255050 171922 255118 171978
rect 255174 171922 255242 171978
rect 255298 171922 255366 171978
rect 255422 171922 255518 171978
rect 254898 154350 255518 171922
rect 254898 154294 254994 154350
rect 255050 154294 255118 154350
rect 255174 154294 255242 154350
rect 255298 154294 255366 154350
rect 255422 154294 255518 154350
rect 254898 154226 255518 154294
rect 254898 154170 254994 154226
rect 255050 154170 255118 154226
rect 255174 154170 255242 154226
rect 255298 154170 255366 154226
rect 255422 154170 255518 154226
rect 254898 154102 255518 154170
rect 254898 154046 254994 154102
rect 255050 154046 255118 154102
rect 255174 154046 255242 154102
rect 255298 154046 255366 154102
rect 255422 154046 255518 154102
rect 254898 153978 255518 154046
rect 254898 153922 254994 153978
rect 255050 153922 255118 153978
rect 255174 153922 255242 153978
rect 255298 153922 255366 153978
rect 255422 153922 255518 153978
rect 254898 136350 255518 153922
rect 254898 136294 254994 136350
rect 255050 136294 255118 136350
rect 255174 136294 255242 136350
rect 255298 136294 255366 136350
rect 255422 136294 255518 136350
rect 254898 136226 255518 136294
rect 254898 136170 254994 136226
rect 255050 136170 255118 136226
rect 255174 136170 255242 136226
rect 255298 136170 255366 136226
rect 255422 136170 255518 136226
rect 254898 136102 255518 136170
rect 254898 136046 254994 136102
rect 255050 136046 255118 136102
rect 255174 136046 255242 136102
rect 255298 136046 255366 136102
rect 255422 136046 255518 136102
rect 254898 135978 255518 136046
rect 254898 135922 254994 135978
rect 255050 135922 255118 135978
rect 255174 135922 255242 135978
rect 255298 135922 255366 135978
rect 255422 135922 255518 135978
rect 254898 118350 255518 135922
rect 254898 118294 254994 118350
rect 255050 118294 255118 118350
rect 255174 118294 255242 118350
rect 255298 118294 255366 118350
rect 255422 118294 255518 118350
rect 254898 118226 255518 118294
rect 254898 118170 254994 118226
rect 255050 118170 255118 118226
rect 255174 118170 255242 118226
rect 255298 118170 255366 118226
rect 255422 118170 255518 118226
rect 254898 118102 255518 118170
rect 254898 118046 254994 118102
rect 255050 118046 255118 118102
rect 255174 118046 255242 118102
rect 255298 118046 255366 118102
rect 255422 118046 255518 118102
rect 254898 117978 255518 118046
rect 254898 117922 254994 117978
rect 255050 117922 255118 117978
rect 255174 117922 255242 117978
rect 255298 117922 255366 117978
rect 255422 117922 255518 117978
rect 254898 100350 255518 117922
rect 254898 100294 254994 100350
rect 255050 100294 255118 100350
rect 255174 100294 255242 100350
rect 255298 100294 255366 100350
rect 255422 100294 255518 100350
rect 254898 100226 255518 100294
rect 254898 100170 254994 100226
rect 255050 100170 255118 100226
rect 255174 100170 255242 100226
rect 255298 100170 255366 100226
rect 255422 100170 255518 100226
rect 254898 100102 255518 100170
rect 254898 100046 254994 100102
rect 255050 100046 255118 100102
rect 255174 100046 255242 100102
rect 255298 100046 255366 100102
rect 255422 100046 255518 100102
rect 254898 99978 255518 100046
rect 254898 99922 254994 99978
rect 255050 99922 255118 99978
rect 255174 99922 255242 99978
rect 255298 99922 255366 99978
rect 255422 99922 255518 99978
rect 254898 82350 255518 99922
rect 254898 82294 254994 82350
rect 255050 82294 255118 82350
rect 255174 82294 255242 82350
rect 255298 82294 255366 82350
rect 255422 82294 255518 82350
rect 254898 82226 255518 82294
rect 254898 82170 254994 82226
rect 255050 82170 255118 82226
rect 255174 82170 255242 82226
rect 255298 82170 255366 82226
rect 255422 82170 255518 82226
rect 254898 82102 255518 82170
rect 254898 82046 254994 82102
rect 255050 82046 255118 82102
rect 255174 82046 255242 82102
rect 255298 82046 255366 82102
rect 255422 82046 255518 82102
rect 254898 81978 255518 82046
rect 254898 81922 254994 81978
rect 255050 81922 255118 81978
rect 255174 81922 255242 81978
rect 255298 81922 255366 81978
rect 255422 81922 255518 81978
rect 251178 58294 251274 58350
rect 251330 58294 251398 58350
rect 251454 58294 251522 58350
rect 251578 58294 251646 58350
rect 251702 58294 251798 58350
rect 251178 58226 251798 58294
rect 251178 58170 251274 58226
rect 251330 58170 251398 58226
rect 251454 58170 251522 58226
rect 251578 58170 251646 58226
rect 251702 58170 251798 58226
rect 251178 58102 251798 58170
rect 251178 58046 251274 58102
rect 251330 58046 251398 58102
rect 251454 58046 251522 58102
rect 251578 58046 251646 58102
rect 251702 58046 251798 58102
rect 251178 57978 251798 58046
rect 251178 57922 251274 57978
rect 251330 57922 251398 57978
rect 251454 57922 251522 57978
rect 251578 57922 251646 57978
rect 251702 57922 251798 57978
rect 251178 40350 251798 57922
rect 251178 40294 251274 40350
rect 251330 40294 251398 40350
rect 251454 40294 251522 40350
rect 251578 40294 251646 40350
rect 251702 40294 251798 40350
rect 251178 40226 251798 40294
rect 251178 40170 251274 40226
rect 251330 40170 251398 40226
rect 251454 40170 251522 40226
rect 251578 40170 251646 40226
rect 251702 40170 251798 40226
rect 251178 40102 251798 40170
rect 251178 40046 251274 40102
rect 251330 40046 251398 40102
rect 251454 40046 251522 40102
rect 251578 40046 251646 40102
rect 251702 40046 251798 40102
rect 251178 39978 251798 40046
rect 251178 39922 251274 39978
rect 251330 39922 251398 39978
rect 251454 39922 251522 39978
rect 251578 39922 251646 39978
rect 251702 39922 251798 39978
rect 251178 22350 251798 39922
rect 251178 22294 251274 22350
rect 251330 22294 251398 22350
rect 251454 22294 251522 22350
rect 251578 22294 251646 22350
rect 251702 22294 251798 22350
rect 251178 22226 251798 22294
rect 251178 22170 251274 22226
rect 251330 22170 251398 22226
rect 251454 22170 251522 22226
rect 251578 22170 251646 22226
rect 251702 22170 251798 22226
rect 251178 22102 251798 22170
rect 251178 22046 251274 22102
rect 251330 22046 251398 22102
rect 251454 22046 251522 22102
rect 251578 22046 251646 22102
rect 251702 22046 251798 22102
rect 251178 21978 251798 22046
rect 251178 21922 251274 21978
rect 251330 21922 251398 21978
rect 251454 21922 251522 21978
rect 251578 21922 251646 21978
rect 251702 21922 251798 21978
rect 248668 4162 248724 4172
rect 250348 13798 250404 13808
rect 250348 4228 250404 13742
rect 250348 4162 250404 4172
rect 251178 4350 251798 21922
rect 251178 4294 251274 4350
rect 251330 4294 251398 4350
rect 251454 4294 251522 4350
rect 251578 4294 251646 4350
rect 251702 4294 251798 4350
rect 251178 4226 251798 4294
rect 251178 4170 251274 4226
rect 251330 4170 251398 4226
rect 251454 4170 251522 4226
rect 251578 4170 251646 4226
rect 251702 4170 251798 4226
rect 224178 -1176 224274 -1120
rect 224330 -1176 224398 -1120
rect 224454 -1176 224522 -1120
rect 224578 -1176 224646 -1120
rect 224702 -1176 224798 -1120
rect 224178 -1244 224798 -1176
rect 224178 -1300 224274 -1244
rect 224330 -1300 224398 -1244
rect 224454 -1300 224522 -1244
rect 224578 -1300 224646 -1244
rect 224702 -1300 224798 -1244
rect 224178 -1368 224798 -1300
rect 224178 -1424 224274 -1368
rect 224330 -1424 224398 -1368
rect 224454 -1424 224522 -1368
rect 224578 -1424 224646 -1368
rect 224702 -1424 224798 -1368
rect 224178 -1492 224798 -1424
rect 224178 -1548 224274 -1492
rect 224330 -1548 224398 -1492
rect 224454 -1548 224522 -1492
rect 224578 -1548 224646 -1492
rect 224702 -1548 224798 -1492
rect 224178 -1644 224798 -1548
rect 251178 4102 251798 4170
rect 252028 64918 252084 64928
rect 252028 4228 252084 64862
rect 252028 4162 252084 4172
rect 253708 64738 253764 64748
rect 253708 4228 253764 64682
rect 253708 4162 253764 4172
rect 254898 64350 255518 81922
rect 281898 597212 282518 598268
rect 281898 597156 281994 597212
rect 282050 597156 282118 597212
rect 282174 597156 282242 597212
rect 282298 597156 282366 597212
rect 282422 597156 282518 597212
rect 281898 597088 282518 597156
rect 281898 597032 281994 597088
rect 282050 597032 282118 597088
rect 282174 597032 282242 597088
rect 282298 597032 282366 597088
rect 282422 597032 282518 597088
rect 281898 596964 282518 597032
rect 281898 596908 281994 596964
rect 282050 596908 282118 596964
rect 282174 596908 282242 596964
rect 282298 596908 282366 596964
rect 282422 596908 282518 596964
rect 281898 596840 282518 596908
rect 281898 596784 281994 596840
rect 282050 596784 282118 596840
rect 282174 596784 282242 596840
rect 282298 596784 282366 596840
rect 282422 596784 282518 596840
rect 281898 580350 282518 596784
rect 281898 580294 281994 580350
rect 282050 580294 282118 580350
rect 282174 580294 282242 580350
rect 282298 580294 282366 580350
rect 282422 580294 282518 580350
rect 281898 580226 282518 580294
rect 281898 580170 281994 580226
rect 282050 580170 282118 580226
rect 282174 580170 282242 580226
rect 282298 580170 282366 580226
rect 282422 580170 282518 580226
rect 281898 580102 282518 580170
rect 281898 580046 281994 580102
rect 282050 580046 282118 580102
rect 282174 580046 282242 580102
rect 282298 580046 282366 580102
rect 282422 580046 282518 580102
rect 281898 579978 282518 580046
rect 281898 579922 281994 579978
rect 282050 579922 282118 579978
rect 282174 579922 282242 579978
rect 282298 579922 282366 579978
rect 282422 579922 282518 579978
rect 281898 562350 282518 579922
rect 281898 562294 281994 562350
rect 282050 562294 282118 562350
rect 282174 562294 282242 562350
rect 282298 562294 282366 562350
rect 282422 562294 282518 562350
rect 281898 562226 282518 562294
rect 281898 562170 281994 562226
rect 282050 562170 282118 562226
rect 282174 562170 282242 562226
rect 282298 562170 282366 562226
rect 282422 562170 282518 562226
rect 281898 562102 282518 562170
rect 281898 562046 281994 562102
rect 282050 562046 282118 562102
rect 282174 562046 282242 562102
rect 282298 562046 282366 562102
rect 282422 562046 282518 562102
rect 281898 561978 282518 562046
rect 281898 561922 281994 561978
rect 282050 561922 282118 561978
rect 282174 561922 282242 561978
rect 282298 561922 282366 561978
rect 282422 561922 282518 561978
rect 281898 544350 282518 561922
rect 281898 544294 281994 544350
rect 282050 544294 282118 544350
rect 282174 544294 282242 544350
rect 282298 544294 282366 544350
rect 282422 544294 282518 544350
rect 281898 544226 282518 544294
rect 281898 544170 281994 544226
rect 282050 544170 282118 544226
rect 282174 544170 282242 544226
rect 282298 544170 282366 544226
rect 282422 544170 282518 544226
rect 281898 544102 282518 544170
rect 281898 544046 281994 544102
rect 282050 544046 282118 544102
rect 282174 544046 282242 544102
rect 282298 544046 282366 544102
rect 282422 544046 282518 544102
rect 281898 543978 282518 544046
rect 281898 543922 281994 543978
rect 282050 543922 282118 543978
rect 282174 543922 282242 543978
rect 282298 543922 282366 543978
rect 282422 543922 282518 543978
rect 281898 526350 282518 543922
rect 281898 526294 281994 526350
rect 282050 526294 282118 526350
rect 282174 526294 282242 526350
rect 282298 526294 282366 526350
rect 282422 526294 282518 526350
rect 281898 526226 282518 526294
rect 281898 526170 281994 526226
rect 282050 526170 282118 526226
rect 282174 526170 282242 526226
rect 282298 526170 282366 526226
rect 282422 526170 282518 526226
rect 281898 526102 282518 526170
rect 281898 526046 281994 526102
rect 282050 526046 282118 526102
rect 282174 526046 282242 526102
rect 282298 526046 282366 526102
rect 282422 526046 282518 526102
rect 281898 525978 282518 526046
rect 281898 525922 281994 525978
rect 282050 525922 282118 525978
rect 282174 525922 282242 525978
rect 282298 525922 282366 525978
rect 282422 525922 282518 525978
rect 281898 508350 282518 525922
rect 281898 508294 281994 508350
rect 282050 508294 282118 508350
rect 282174 508294 282242 508350
rect 282298 508294 282366 508350
rect 282422 508294 282518 508350
rect 281898 508226 282518 508294
rect 281898 508170 281994 508226
rect 282050 508170 282118 508226
rect 282174 508170 282242 508226
rect 282298 508170 282366 508226
rect 282422 508170 282518 508226
rect 281898 508102 282518 508170
rect 281898 508046 281994 508102
rect 282050 508046 282118 508102
rect 282174 508046 282242 508102
rect 282298 508046 282366 508102
rect 282422 508046 282518 508102
rect 281898 507978 282518 508046
rect 281898 507922 281994 507978
rect 282050 507922 282118 507978
rect 282174 507922 282242 507978
rect 282298 507922 282366 507978
rect 282422 507922 282518 507978
rect 281898 490350 282518 507922
rect 281898 490294 281994 490350
rect 282050 490294 282118 490350
rect 282174 490294 282242 490350
rect 282298 490294 282366 490350
rect 282422 490294 282518 490350
rect 281898 490226 282518 490294
rect 281898 490170 281994 490226
rect 282050 490170 282118 490226
rect 282174 490170 282242 490226
rect 282298 490170 282366 490226
rect 282422 490170 282518 490226
rect 281898 490102 282518 490170
rect 281898 490046 281994 490102
rect 282050 490046 282118 490102
rect 282174 490046 282242 490102
rect 282298 490046 282366 490102
rect 282422 490046 282518 490102
rect 281898 489978 282518 490046
rect 281898 489922 281994 489978
rect 282050 489922 282118 489978
rect 282174 489922 282242 489978
rect 282298 489922 282366 489978
rect 282422 489922 282518 489978
rect 281898 472350 282518 489922
rect 281898 472294 281994 472350
rect 282050 472294 282118 472350
rect 282174 472294 282242 472350
rect 282298 472294 282366 472350
rect 282422 472294 282518 472350
rect 281898 472226 282518 472294
rect 281898 472170 281994 472226
rect 282050 472170 282118 472226
rect 282174 472170 282242 472226
rect 282298 472170 282366 472226
rect 282422 472170 282518 472226
rect 281898 472102 282518 472170
rect 281898 472046 281994 472102
rect 282050 472046 282118 472102
rect 282174 472046 282242 472102
rect 282298 472046 282366 472102
rect 282422 472046 282518 472102
rect 281898 471978 282518 472046
rect 281898 471922 281994 471978
rect 282050 471922 282118 471978
rect 282174 471922 282242 471978
rect 282298 471922 282366 471978
rect 282422 471922 282518 471978
rect 281898 454350 282518 471922
rect 281898 454294 281994 454350
rect 282050 454294 282118 454350
rect 282174 454294 282242 454350
rect 282298 454294 282366 454350
rect 282422 454294 282518 454350
rect 281898 454226 282518 454294
rect 281898 454170 281994 454226
rect 282050 454170 282118 454226
rect 282174 454170 282242 454226
rect 282298 454170 282366 454226
rect 282422 454170 282518 454226
rect 281898 454102 282518 454170
rect 281898 454046 281994 454102
rect 282050 454046 282118 454102
rect 282174 454046 282242 454102
rect 282298 454046 282366 454102
rect 282422 454046 282518 454102
rect 281898 453978 282518 454046
rect 281898 453922 281994 453978
rect 282050 453922 282118 453978
rect 282174 453922 282242 453978
rect 282298 453922 282366 453978
rect 282422 453922 282518 453978
rect 281898 436350 282518 453922
rect 281898 436294 281994 436350
rect 282050 436294 282118 436350
rect 282174 436294 282242 436350
rect 282298 436294 282366 436350
rect 282422 436294 282518 436350
rect 281898 436226 282518 436294
rect 281898 436170 281994 436226
rect 282050 436170 282118 436226
rect 282174 436170 282242 436226
rect 282298 436170 282366 436226
rect 282422 436170 282518 436226
rect 281898 436102 282518 436170
rect 281898 436046 281994 436102
rect 282050 436046 282118 436102
rect 282174 436046 282242 436102
rect 282298 436046 282366 436102
rect 282422 436046 282518 436102
rect 281898 435978 282518 436046
rect 281898 435922 281994 435978
rect 282050 435922 282118 435978
rect 282174 435922 282242 435978
rect 282298 435922 282366 435978
rect 282422 435922 282518 435978
rect 281898 418350 282518 435922
rect 281898 418294 281994 418350
rect 282050 418294 282118 418350
rect 282174 418294 282242 418350
rect 282298 418294 282366 418350
rect 282422 418294 282518 418350
rect 281898 418226 282518 418294
rect 281898 418170 281994 418226
rect 282050 418170 282118 418226
rect 282174 418170 282242 418226
rect 282298 418170 282366 418226
rect 282422 418170 282518 418226
rect 281898 418102 282518 418170
rect 281898 418046 281994 418102
rect 282050 418046 282118 418102
rect 282174 418046 282242 418102
rect 282298 418046 282366 418102
rect 282422 418046 282518 418102
rect 281898 417978 282518 418046
rect 281898 417922 281994 417978
rect 282050 417922 282118 417978
rect 282174 417922 282242 417978
rect 282298 417922 282366 417978
rect 282422 417922 282518 417978
rect 281898 400350 282518 417922
rect 281898 400294 281994 400350
rect 282050 400294 282118 400350
rect 282174 400294 282242 400350
rect 282298 400294 282366 400350
rect 282422 400294 282518 400350
rect 281898 400226 282518 400294
rect 281898 400170 281994 400226
rect 282050 400170 282118 400226
rect 282174 400170 282242 400226
rect 282298 400170 282366 400226
rect 282422 400170 282518 400226
rect 281898 400102 282518 400170
rect 281898 400046 281994 400102
rect 282050 400046 282118 400102
rect 282174 400046 282242 400102
rect 282298 400046 282366 400102
rect 282422 400046 282518 400102
rect 281898 399978 282518 400046
rect 281898 399922 281994 399978
rect 282050 399922 282118 399978
rect 282174 399922 282242 399978
rect 282298 399922 282366 399978
rect 282422 399922 282518 399978
rect 281898 382350 282518 399922
rect 281898 382294 281994 382350
rect 282050 382294 282118 382350
rect 282174 382294 282242 382350
rect 282298 382294 282366 382350
rect 282422 382294 282518 382350
rect 281898 382226 282518 382294
rect 281898 382170 281994 382226
rect 282050 382170 282118 382226
rect 282174 382170 282242 382226
rect 282298 382170 282366 382226
rect 282422 382170 282518 382226
rect 281898 382102 282518 382170
rect 281898 382046 281994 382102
rect 282050 382046 282118 382102
rect 282174 382046 282242 382102
rect 282298 382046 282366 382102
rect 282422 382046 282518 382102
rect 281898 381978 282518 382046
rect 281898 381922 281994 381978
rect 282050 381922 282118 381978
rect 282174 381922 282242 381978
rect 282298 381922 282366 381978
rect 282422 381922 282518 381978
rect 281898 364350 282518 381922
rect 281898 364294 281994 364350
rect 282050 364294 282118 364350
rect 282174 364294 282242 364350
rect 282298 364294 282366 364350
rect 282422 364294 282518 364350
rect 281898 364226 282518 364294
rect 281898 364170 281994 364226
rect 282050 364170 282118 364226
rect 282174 364170 282242 364226
rect 282298 364170 282366 364226
rect 282422 364170 282518 364226
rect 281898 364102 282518 364170
rect 281898 364046 281994 364102
rect 282050 364046 282118 364102
rect 282174 364046 282242 364102
rect 282298 364046 282366 364102
rect 282422 364046 282518 364102
rect 281898 363978 282518 364046
rect 281898 363922 281994 363978
rect 282050 363922 282118 363978
rect 282174 363922 282242 363978
rect 282298 363922 282366 363978
rect 282422 363922 282518 363978
rect 281898 346350 282518 363922
rect 281898 346294 281994 346350
rect 282050 346294 282118 346350
rect 282174 346294 282242 346350
rect 282298 346294 282366 346350
rect 282422 346294 282518 346350
rect 281898 346226 282518 346294
rect 281898 346170 281994 346226
rect 282050 346170 282118 346226
rect 282174 346170 282242 346226
rect 282298 346170 282366 346226
rect 282422 346170 282518 346226
rect 281898 346102 282518 346170
rect 281898 346046 281994 346102
rect 282050 346046 282118 346102
rect 282174 346046 282242 346102
rect 282298 346046 282366 346102
rect 282422 346046 282518 346102
rect 281898 345978 282518 346046
rect 281898 345922 281994 345978
rect 282050 345922 282118 345978
rect 282174 345922 282242 345978
rect 282298 345922 282366 345978
rect 282422 345922 282518 345978
rect 281898 328350 282518 345922
rect 281898 328294 281994 328350
rect 282050 328294 282118 328350
rect 282174 328294 282242 328350
rect 282298 328294 282366 328350
rect 282422 328294 282518 328350
rect 281898 328226 282518 328294
rect 281898 328170 281994 328226
rect 282050 328170 282118 328226
rect 282174 328170 282242 328226
rect 282298 328170 282366 328226
rect 282422 328170 282518 328226
rect 281898 328102 282518 328170
rect 281898 328046 281994 328102
rect 282050 328046 282118 328102
rect 282174 328046 282242 328102
rect 282298 328046 282366 328102
rect 282422 328046 282518 328102
rect 281898 327978 282518 328046
rect 281898 327922 281994 327978
rect 282050 327922 282118 327978
rect 282174 327922 282242 327978
rect 282298 327922 282366 327978
rect 282422 327922 282518 327978
rect 281898 310350 282518 327922
rect 281898 310294 281994 310350
rect 282050 310294 282118 310350
rect 282174 310294 282242 310350
rect 282298 310294 282366 310350
rect 282422 310294 282518 310350
rect 281898 310226 282518 310294
rect 281898 310170 281994 310226
rect 282050 310170 282118 310226
rect 282174 310170 282242 310226
rect 282298 310170 282366 310226
rect 282422 310170 282518 310226
rect 281898 310102 282518 310170
rect 281898 310046 281994 310102
rect 282050 310046 282118 310102
rect 282174 310046 282242 310102
rect 282298 310046 282366 310102
rect 282422 310046 282518 310102
rect 281898 309978 282518 310046
rect 281898 309922 281994 309978
rect 282050 309922 282118 309978
rect 282174 309922 282242 309978
rect 282298 309922 282366 309978
rect 282422 309922 282518 309978
rect 281898 292350 282518 309922
rect 281898 292294 281994 292350
rect 282050 292294 282118 292350
rect 282174 292294 282242 292350
rect 282298 292294 282366 292350
rect 282422 292294 282518 292350
rect 281898 292226 282518 292294
rect 281898 292170 281994 292226
rect 282050 292170 282118 292226
rect 282174 292170 282242 292226
rect 282298 292170 282366 292226
rect 282422 292170 282518 292226
rect 281898 292102 282518 292170
rect 281898 292046 281994 292102
rect 282050 292046 282118 292102
rect 282174 292046 282242 292102
rect 282298 292046 282366 292102
rect 282422 292046 282518 292102
rect 281898 291978 282518 292046
rect 281898 291922 281994 291978
rect 282050 291922 282118 291978
rect 282174 291922 282242 291978
rect 282298 291922 282366 291978
rect 282422 291922 282518 291978
rect 281898 274350 282518 291922
rect 281898 274294 281994 274350
rect 282050 274294 282118 274350
rect 282174 274294 282242 274350
rect 282298 274294 282366 274350
rect 282422 274294 282518 274350
rect 281898 274226 282518 274294
rect 281898 274170 281994 274226
rect 282050 274170 282118 274226
rect 282174 274170 282242 274226
rect 282298 274170 282366 274226
rect 282422 274170 282518 274226
rect 281898 274102 282518 274170
rect 281898 274046 281994 274102
rect 282050 274046 282118 274102
rect 282174 274046 282242 274102
rect 282298 274046 282366 274102
rect 282422 274046 282518 274102
rect 281898 273978 282518 274046
rect 281898 273922 281994 273978
rect 282050 273922 282118 273978
rect 282174 273922 282242 273978
rect 282298 273922 282366 273978
rect 282422 273922 282518 273978
rect 281898 256350 282518 273922
rect 281898 256294 281994 256350
rect 282050 256294 282118 256350
rect 282174 256294 282242 256350
rect 282298 256294 282366 256350
rect 282422 256294 282518 256350
rect 281898 256226 282518 256294
rect 281898 256170 281994 256226
rect 282050 256170 282118 256226
rect 282174 256170 282242 256226
rect 282298 256170 282366 256226
rect 282422 256170 282518 256226
rect 281898 256102 282518 256170
rect 281898 256046 281994 256102
rect 282050 256046 282118 256102
rect 282174 256046 282242 256102
rect 282298 256046 282366 256102
rect 282422 256046 282518 256102
rect 281898 255978 282518 256046
rect 281898 255922 281994 255978
rect 282050 255922 282118 255978
rect 282174 255922 282242 255978
rect 282298 255922 282366 255978
rect 282422 255922 282518 255978
rect 281898 238350 282518 255922
rect 281898 238294 281994 238350
rect 282050 238294 282118 238350
rect 282174 238294 282242 238350
rect 282298 238294 282366 238350
rect 282422 238294 282518 238350
rect 281898 238226 282518 238294
rect 281898 238170 281994 238226
rect 282050 238170 282118 238226
rect 282174 238170 282242 238226
rect 282298 238170 282366 238226
rect 282422 238170 282518 238226
rect 281898 238102 282518 238170
rect 281898 238046 281994 238102
rect 282050 238046 282118 238102
rect 282174 238046 282242 238102
rect 282298 238046 282366 238102
rect 282422 238046 282518 238102
rect 281898 237978 282518 238046
rect 281898 237922 281994 237978
rect 282050 237922 282118 237978
rect 282174 237922 282242 237978
rect 282298 237922 282366 237978
rect 282422 237922 282518 237978
rect 281898 220350 282518 237922
rect 281898 220294 281994 220350
rect 282050 220294 282118 220350
rect 282174 220294 282242 220350
rect 282298 220294 282366 220350
rect 282422 220294 282518 220350
rect 281898 220226 282518 220294
rect 281898 220170 281994 220226
rect 282050 220170 282118 220226
rect 282174 220170 282242 220226
rect 282298 220170 282366 220226
rect 282422 220170 282518 220226
rect 281898 220102 282518 220170
rect 281898 220046 281994 220102
rect 282050 220046 282118 220102
rect 282174 220046 282242 220102
rect 282298 220046 282366 220102
rect 282422 220046 282518 220102
rect 281898 219978 282518 220046
rect 281898 219922 281994 219978
rect 282050 219922 282118 219978
rect 282174 219922 282242 219978
rect 282298 219922 282366 219978
rect 282422 219922 282518 219978
rect 281898 202350 282518 219922
rect 281898 202294 281994 202350
rect 282050 202294 282118 202350
rect 282174 202294 282242 202350
rect 282298 202294 282366 202350
rect 282422 202294 282518 202350
rect 281898 202226 282518 202294
rect 281898 202170 281994 202226
rect 282050 202170 282118 202226
rect 282174 202170 282242 202226
rect 282298 202170 282366 202226
rect 282422 202170 282518 202226
rect 281898 202102 282518 202170
rect 281898 202046 281994 202102
rect 282050 202046 282118 202102
rect 282174 202046 282242 202102
rect 282298 202046 282366 202102
rect 282422 202046 282518 202102
rect 281898 201978 282518 202046
rect 281898 201922 281994 201978
rect 282050 201922 282118 201978
rect 282174 201922 282242 201978
rect 282298 201922 282366 201978
rect 282422 201922 282518 201978
rect 281898 184350 282518 201922
rect 281898 184294 281994 184350
rect 282050 184294 282118 184350
rect 282174 184294 282242 184350
rect 282298 184294 282366 184350
rect 282422 184294 282518 184350
rect 281898 184226 282518 184294
rect 281898 184170 281994 184226
rect 282050 184170 282118 184226
rect 282174 184170 282242 184226
rect 282298 184170 282366 184226
rect 282422 184170 282518 184226
rect 281898 184102 282518 184170
rect 281898 184046 281994 184102
rect 282050 184046 282118 184102
rect 282174 184046 282242 184102
rect 282298 184046 282366 184102
rect 282422 184046 282518 184102
rect 281898 183978 282518 184046
rect 281898 183922 281994 183978
rect 282050 183922 282118 183978
rect 282174 183922 282242 183978
rect 282298 183922 282366 183978
rect 282422 183922 282518 183978
rect 281898 166350 282518 183922
rect 281898 166294 281994 166350
rect 282050 166294 282118 166350
rect 282174 166294 282242 166350
rect 282298 166294 282366 166350
rect 282422 166294 282518 166350
rect 281898 166226 282518 166294
rect 281898 166170 281994 166226
rect 282050 166170 282118 166226
rect 282174 166170 282242 166226
rect 282298 166170 282366 166226
rect 282422 166170 282518 166226
rect 281898 166102 282518 166170
rect 281898 166046 281994 166102
rect 282050 166046 282118 166102
rect 282174 166046 282242 166102
rect 282298 166046 282366 166102
rect 282422 166046 282518 166102
rect 281898 165978 282518 166046
rect 281898 165922 281994 165978
rect 282050 165922 282118 165978
rect 282174 165922 282242 165978
rect 282298 165922 282366 165978
rect 282422 165922 282518 165978
rect 281898 148350 282518 165922
rect 281898 148294 281994 148350
rect 282050 148294 282118 148350
rect 282174 148294 282242 148350
rect 282298 148294 282366 148350
rect 282422 148294 282518 148350
rect 281898 148226 282518 148294
rect 281898 148170 281994 148226
rect 282050 148170 282118 148226
rect 282174 148170 282242 148226
rect 282298 148170 282366 148226
rect 282422 148170 282518 148226
rect 281898 148102 282518 148170
rect 281898 148046 281994 148102
rect 282050 148046 282118 148102
rect 282174 148046 282242 148102
rect 282298 148046 282366 148102
rect 282422 148046 282518 148102
rect 281898 147978 282518 148046
rect 281898 147922 281994 147978
rect 282050 147922 282118 147978
rect 282174 147922 282242 147978
rect 282298 147922 282366 147978
rect 282422 147922 282518 147978
rect 281898 130350 282518 147922
rect 281898 130294 281994 130350
rect 282050 130294 282118 130350
rect 282174 130294 282242 130350
rect 282298 130294 282366 130350
rect 282422 130294 282518 130350
rect 281898 130226 282518 130294
rect 281898 130170 281994 130226
rect 282050 130170 282118 130226
rect 282174 130170 282242 130226
rect 282298 130170 282366 130226
rect 282422 130170 282518 130226
rect 281898 130102 282518 130170
rect 281898 130046 281994 130102
rect 282050 130046 282118 130102
rect 282174 130046 282242 130102
rect 282298 130046 282366 130102
rect 282422 130046 282518 130102
rect 281898 129978 282518 130046
rect 281898 129922 281994 129978
rect 282050 129922 282118 129978
rect 282174 129922 282242 129978
rect 282298 129922 282366 129978
rect 282422 129922 282518 129978
rect 281898 112350 282518 129922
rect 281898 112294 281994 112350
rect 282050 112294 282118 112350
rect 282174 112294 282242 112350
rect 282298 112294 282366 112350
rect 282422 112294 282518 112350
rect 281898 112226 282518 112294
rect 281898 112170 281994 112226
rect 282050 112170 282118 112226
rect 282174 112170 282242 112226
rect 282298 112170 282366 112226
rect 282422 112170 282518 112226
rect 281898 112102 282518 112170
rect 281898 112046 281994 112102
rect 282050 112046 282118 112102
rect 282174 112046 282242 112102
rect 282298 112046 282366 112102
rect 282422 112046 282518 112102
rect 281898 111978 282518 112046
rect 281898 111922 281994 111978
rect 282050 111922 282118 111978
rect 282174 111922 282242 111978
rect 282298 111922 282366 111978
rect 282422 111922 282518 111978
rect 281898 94350 282518 111922
rect 281898 94294 281994 94350
rect 282050 94294 282118 94350
rect 282174 94294 282242 94350
rect 282298 94294 282366 94350
rect 282422 94294 282518 94350
rect 281898 94226 282518 94294
rect 281898 94170 281994 94226
rect 282050 94170 282118 94226
rect 282174 94170 282242 94226
rect 282298 94170 282366 94226
rect 282422 94170 282518 94226
rect 281898 94102 282518 94170
rect 281898 94046 281994 94102
rect 282050 94046 282118 94102
rect 282174 94046 282242 94102
rect 282298 94046 282366 94102
rect 282422 94046 282518 94102
rect 281898 93978 282518 94046
rect 281898 93922 281994 93978
rect 282050 93922 282118 93978
rect 282174 93922 282242 93978
rect 282298 93922 282366 93978
rect 282422 93922 282518 93978
rect 281898 76350 282518 93922
rect 281898 76294 281994 76350
rect 282050 76294 282118 76350
rect 282174 76294 282242 76350
rect 282298 76294 282366 76350
rect 282422 76294 282518 76350
rect 281898 76226 282518 76294
rect 281898 76170 281994 76226
rect 282050 76170 282118 76226
rect 282174 76170 282242 76226
rect 282298 76170 282366 76226
rect 282422 76170 282518 76226
rect 281898 76102 282518 76170
rect 281898 76046 281994 76102
rect 282050 76046 282118 76102
rect 282174 76046 282242 76102
rect 282298 76046 282366 76102
rect 282422 76046 282518 76102
rect 281898 75978 282518 76046
rect 281898 75922 281994 75978
rect 282050 75922 282118 75978
rect 282174 75922 282242 75978
rect 282298 75922 282366 75978
rect 282422 75922 282518 75978
rect 263788 71038 263844 71048
rect 254898 64294 254994 64350
rect 255050 64294 255118 64350
rect 255174 64294 255242 64350
rect 255298 64294 255366 64350
rect 255422 64294 255518 64350
rect 254898 64226 255518 64294
rect 254898 64170 254994 64226
rect 255050 64170 255118 64226
rect 255174 64170 255242 64226
rect 255298 64170 255366 64226
rect 255422 64170 255518 64226
rect 254898 64102 255518 64170
rect 254898 64046 254994 64102
rect 255050 64046 255118 64102
rect 255174 64046 255242 64102
rect 255298 64046 255366 64102
rect 255422 64046 255518 64102
rect 254898 63978 255518 64046
rect 254898 63922 254994 63978
rect 255050 63922 255118 63978
rect 255174 63922 255242 63978
rect 255298 63922 255366 63978
rect 255422 63922 255518 63978
rect 254898 46350 255518 63922
rect 254898 46294 254994 46350
rect 255050 46294 255118 46350
rect 255174 46294 255242 46350
rect 255298 46294 255366 46350
rect 255422 46294 255518 46350
rect 254898 46226 255518 46294
rect 254898 46170 254994 46226
rect 255050 46170 255118 46226
rect 255174 46170 255242 46226
rect 255298 46170 255366 46226
rect 255422 46170 255518 46226
rect 254898 46102 255518 46170
rect 254898 46046 254994 46102
rect 255050 46046 255118 46102
rect 255174 46046 255242 46102
rect 255298 46046 255366 46102
rect 255422 46046 255518 46102
rect 254898 45978 255518 46046
rect 254898 45922 254994 45978
rect 255050 45922 255118 45978
rect 255174 45922 255242 45978
rect 255298 45922 255366 45978
rect 255422 45922 255518 45978
rect 254898 28350 255518 45922
rect 254898 28294 254994 28350
rect 255050 28294 255118 28350
rect 255174 28294 255242 28350
rect 255298 28294 255366 28350
rect 255422 28294 255518 28350
rect 254898 28226 255518 28294
rect 254898 28170 254994 28226
rect 255050 28170 255118 28226
rect 255174 28170 255242 28226
rect 255298 28170 255366 28226
rect 255422 28170 255518 28226
rect 254898 28102 255518 28170
rect 254898 28046 254994 28102
rect 255050 28046 255118 28102
rect 255174 28046 255242 28102
rect 255298 28046 255366 28102
rect 255422 28046 255518 28102
rect 254898 27978 255518 28046
rect 254898 27922 254994 27978
rect 255050 27922 255118 27978
rect 255174 27922 255242 27978
rect 255298 27922 255366 27978
rect 255422 27922 255518 27978
rect 254898 10350 255518 27922
rect 258748 66178 258804 66188
rect 258748 20188 258804 66122
rect 260428 42418 260484 42428
rect 258748 20132 258916 20188
rect 254898 10294 254994 10350
rect 255050 10294 255118 10350
rect 255174 10294 255242 10350
rect 255298 10294 255366 10350
rect 255422 10294 255518 10350
rect 254898 10226 255518 10294
rect 254898 10170 254994 10226
rect 255050 10170 255118 10226
rect 255174 10170 255242 10226
rect 255298 10170 255366 10226
rect 255422 10170 255518 10226
rect 254898 10102 255518 10170
rect 254898 10046 254994 10102
rect 255050 10046 255118 10102
rect 255174 10046 255242 10102
rect 255298 10046 255366 10102
rect 255422 10046 255518 10102
rect 254898 9978 255518 10046
rect 254898 9922 254994 9978
rect 255050 9922 255118 9978
rect 255174 9922 255242 9978
rect 255298 9922 255366 9978
rect 255422 9922 255518 9978
rect 251178 4046 251274 4102
rect 251330 4046 251398 4102
rect 251454 4046 251522 4102
rect 251578 4046 251646 4102
rect 251702 4046 251798 4102
rect 251178 3978 251798 4046
rect 251178 3922 251274 3978
rect 251330 3922 251398 3978
rect 251454 3922 251522 3978
rect 251578 3922 251646 3978
rect 251702 3922 251798 3978
rect 251178 -160 251798 3922
rect 251178 -216 251274 -160
rect 251330 -216 251398 -160
rect 251454 -216 251522 -160
rect 251578 -216 251646 -160
rect 251702 -216 251798 -160
rect 251178 -284 251798 -216
rect 251178 -340 251274 -284
rect 251330 -340 251398 -284
rect 251454 -340 251522 -284
rect 251578 -340 251646 -284
rect 251702 -340 251798 -284
rect 251178 -408 251798 -340
rect 251178 -464 251274 -408
rect 251330 -464 251398 -408
rect 251454 -464 251522 -408
rect 251578 -464 251646 -408
rect 251702 -464 251798 -408
rect 251178 -532 251798 -464
rect 251178 -588 251274 -532
rect 251330 -588 251398 -532
rect 251454 -588 251522 -532
rect 251578 -588 251646 -532
rect 251702 -588 251798 -532
rect 251178 -1644 251798 -588
rect 254898 -1120 255518 9922
rect 257068 7138 257124 7148
rect 257068 3556 257124 7082
rect 258860 4228 258916 20132
rect 258860 4162 258916 4172
rect 260428 4228 260484 42362
rect 260428 4162 260484 4172
rect 262108 15598 262164 15608
rect 262108 4228 262164 15542
rect 262108 4162 262164 4172
rect 263788 4228 263844 70982
rect 273868 59698 273924 59708
rect 263788 4162 263844 4172
rect 265468 56098 265524 56108
rect 265468 4228 265524 56042
rect 273868 20188 273924 59642
rect 281898 58350 282518 75922
rect 281898 58294 281994 58350
rect 282050 58294 282118 58350
rect 282174 58294 282242 58350
rect 282298 58294 282366 58350
rect 282422 58294 282518 58350
rect 281898 58226 282518 58294
rect 281898 58170 281994 58226
rect 282050 58170 282118 58226
rect 282174 58170 282242 58226
rect 282298 58170 282366 58226
rect 282422 58170 282518 58226
rect 281898 58102 282518 58170
rect 281898 58046 281994 58102
rect 282050 58046 282118 58102
rect 282174 58046 282242 58102
rect 282298 58046 282366 58102
rect 282422 58046 282518 58102
rect 281898 57978 282518 58046
rect 281898 57922 281994 57978
rect 282050 57922 282118 57978
rect 282174 57922 282242 57978
rect 282298 57922 282366 57978
rect 282422 57922 282518 57978
rect 281898 40350 282518 57922
rect 285618 598172 286238 598268
rect 285618 598116 285714 598172
rect 285770 598116 285838 598172
rect 285894 598116 285962 598172
rect 286018 598116 286086 598172
rect 286142 598116 286238 598172
rect 285618 598048 286238 598116
rect 285618 597992 285714 598048
rect 285770 597992 285838 598048
rect 285894 597992 285962 598048
rect 286018 597992 286086 598048
rect 286142 597992 286238 598048
rect 285618 597924 286238 597992
rect 285618 597868 285714 597924
rect 285770 597868 285838 597924
rect 285894 597868 285962 597924
rect 286018 597868 286086 597924
rect 286142 597868 286238 597924
rect 285618 597800 286238 597868
rect 285618 597744 285714 597800
rect 285770 597744 285838 597800
rect 285894 597744 285962 597800
rect 286018 597744 286086 597800
rect 286142 597744 286238 597800
rect 285618 586350 286238 597744
rect 312618 597212 313238 598268
rect 312618 597156 312714 597212
rect 312770 597156 312838 597212
rect 312894 597156 312962 597212
rect 313018 597156 313086 597212
rect 313142 597156 313238 597212
rect 312618 597088 313238 597156
rect 312618 597032 312714 597088
rect 312770 597032 312838 597088
rect 312894 597032 312962 597088
rect 313018 597032 313086 597088
rect 313142 597032 313238 597088
rect 312618 596964 313238 597032
rect 312618 596908 312714 596964
rect 312770 596908 312838 596964
rect 312894 596908 312962 596964
rect 313018 596908 313086 596964
rect 313142 596908 313238 596964
rect 312618 596840 313238 596908
rect 312618 596784 312714 596840
rect 312770 596784 312838 596840
rect 312894 596784 312962 596840
rect 313018 596784 313086 596840
rect 313142 596784 313238 596840
rect 285618 586294 285714 586350
rect 285770 586294 285838 586350
rect 285894 586294 285962 586350
rect 286018 586294 286086 586350
rect 286142 586294 286238 586350
rect 285618 586226 286238 586294
rect 285618 586170 285714 586226
rect 285770 586170 285838 586226
rect 285894 586170 285962 586226
rect 286018 586170 286086 586226
rect 286142 586170 286238 586226
rect 285618 586102 286238 586170
rect 285618 586046 285714 586102
rect 285770 586046 285838 586102
rect 285894 586046 285962 586102
rect 286018 586046 286086 586102
rect 286142 586046 286238 586102
rect 285618 585978 286238 586046
rect 285618 585922 285714 585978
rect 285770 585922 285838 585978
rect 285894 585922 285962 585978
rect 286018 585922 286086 585978
rect 286142 585922 286238 585978
rect 285618 568350 286238 585922
rect 285618 568294 285714 568350
rect 285770 568294 285838 568350
rect 285894 568294 285962 568350
rect 286018 568294 286086 568350
rect 286142 568294 286238 568350
rect 285618 568226 286238 568294
rect 285618 568170 285714 568226
rect 285770 568170 285838 568226
rect 285894 568170 285962 568226
rect 286018 568170 286086 568226
rect 286142 568170 286238 568226
rect 285618 568102 286238 568170
rect 285618 568046 285714 568102
rect 285770 568046 285838 568102
rect 285894 568046 285962 568102
rect 286018 568046 286086 568102
rect 286142 568046 286238 568102
rect 285618 567978 286238 568046
rect 285618 567922 285714 567978
rect 285770 567922 285838 567978
rect 285894 567922 285962 567978
rect 286018 567922 286086 567978
rect 286142 567922 286238 567978
rect 285618 550350 286238 567922
rect 285618 550294 285714 550350
rect 285770 550294 285838 550350
rect 285894 550294 285962 550350
rect 286018 550294 286086 550350
rect 286142 550294 286238 550350
rect 285618 550226 286238 550294
rect 285618 550170 285714 550226
rect 285770 550170 285838 550226
rect 285894 550170 285962 550226
rect 286018 550170 286086 550226
rect 286142 550170 286238 550226
rect 285618 550102 286238 550170
rect 285618 550046 285714 550102
rect 285770 550046 285838 550102
rect 285894 550046 285962 550102
rect 286018 550046 286086 550102
rect 286142 550046 286238 550102
rect 285618 549978 286238 550046
rect 285618 549922 285714 549978
rect 285770 549922 285838 549978
rect 285894 549922 285962 549978
rect 286018 549922 286086 549978
rect 286142 549922 286238 549978
rect 285618 532350 286238 549922
rect 285618 532294 285714 532350
rect 285770 532294 285838 532350
rect 285894 532294 285962 532350
rect 286018 532294 286086 532350
rect 286142 532294 286238 532350
rect 285618 532226 286238 532294
rect 285618 532170 285714 532226
rect 285770 532170 285838 532226
rect 285894 532170 285962 532226
rect 286018 532170 286086 532226
rect 286142 532170 286238 532226
rect 285618 532102 286238 532170
rect 285618 532046 285714 532102
rect 285770 532046 285838 532102
rect 285894 532046 285962 532102
rect 286018 532046 286086 532102
rect 286142 532046 286238 532102
rect 285618 531978 286238 532046
rect 285618 531922 285714 531978
rect 285770 531922 285838 531978
rect 285894 531922 285962 531978
rect 286018 531922 286086 531978
rect 286142 531922 286238 531978
rect 285618 514350 286238 531922
rect 285618 514294 285714 514350
rect 285770 514294 285838 514350
rect 285894 514294 285962 514350
rect 286018 514294 286086 514350
rect 286142 514294 286238 514350
rect 285618 514226 286238 514294
rect 285618 514170 285714 514226
rect 285770 514170 285838 514226
rect 285894 514170 285962 514226
rect 286018 514170 286086 514226
rect 286142 514170 286238 514226
rect 285618 514102 286238 514170
rect 285618 514046 285714 514102
rect 285770 514046 285838 514102
rect 285894 514046 285962 514102
rect 286018 514046 286086 514102
rect 286142 514046 286238 514102
rect 285618 513978 286238 514046
rect 285618 513922 285714 513978
rect 285770 513922 285838 513978
rect 285894 513922 285962 513978
rect 286018 513922 286086 513978
rect 286142 513922 286238 513978
rect 285618 496350 286238 513922
rect 285618 496294 285714 496350
rect 285770 496294 285838 496350
rect 285894 496294 285962 496350
rect 286018 496294 286086 496350
rect 286142 496294 286238 496350
rect 285618 496226 286238 496294
rect 285618 496170 285714 496226
rect 285770 496170 285838 496226
rect 285894 496170 285962 496226
rect 286018 496170 286086 496226
rect 286142 496170 286238 496226
rect 285618 496102 286238 496170
rect 285618 496046 285714 496102
rect 285770 496046 285838 496102
rect 285894 496046 285962 496102
rect 286018 496046 286086 496102
rect 286142 496046 286238 496102
rect 285618 495978 286238 496046
rect 285618 495922 285714 495978
rect 285770 495922 285838 495978
rect 285894 495922 285962 495978
rect 286018 495922 286086 495978
rect 286142 495922 286238 495978
rect 285618 478350 286238 495922
rect 285618 478294 285714 478350
rect 285770 478294 285838 478350
rect 285894 478294 285962 478350
rect 286018 478294 286086 478350
rect 286142 478294 286238 478350
rect 285618 478226 286238 478294
rect 285618 478170 285714 478226
rect 285770 478170 285838 478226
rect 285894 478170 285962 478226
rect 286018 478170 286086 478226
rect 286142 478170 286238 478226
rect 285618 478102 286238 478170
rect 285618 478046 285714 478102
rect 285770 478046 285838 478102
rect 285894 478046 285962 478102
rect 286018 478046 286086 478102
rect 286142 478046 286238 478102
rect 285618 477978 286238 478046
rect 285618 477922 285714 477978
rect 285770 477922 285838 477978
rect 285894 477922 285962 477978
rect 286018 477922 286086 477978
rect 286142 477922 286238 477978
rect 285618 460350 286238 477922
rect 285618 460294 285714 460350
rect 285770 460294 285838 460350
rect 285894 460294 285962 460350
rect 286018 460294 286086 460350
rect 286142 460294 286238 460350
rect 285618 460226 286238 460294
rect 285618 460170 285714 460226
rect 285770 460170 285838 460226
rect 285894 460170 285962 460226
rect 286018 460170 286086 460226
rect 286142 460170 286238 460226
rect 285618 460102 286238 460170
rect 285618 460046 285714 460102
rect 285770 460046 285838 460102
rect 285894 460046 285962 460102
rect 286018 460046 286086 460102
rect 286142 460046 286238 460102
rect 285618 459978 286238 460046
rect 285618 459922 285714 459978
rect 285770 459922 285838 459978
rect 285894 459922 285962 459978
rect 286018 459922 286086 459978
rect 286142 459922 286238 459978
rect 285618 442350 286238 459922
rect 285618 442294 285714 442350
rect 285770 442294 285838 442350
rect 285894 442294 285962 442350
rect 286018 442294 286086 442350
rect 286142 442294 286238 442350
rect 285618 442226 286238 442294
rect 285618 442170 285714 442226
rect 285770 442170 285838 442226
rect 285894 442170 285962 442226
rect 286018 442170 286086 442226
rect 286142 442170 286238 442226
rect 285618 442102 286238 442170
rect 285618 442046 285714 442102
rect 285770 442046 285838 442102
rect 285894 442046 285962 442102
rect 286018 442046 286086 442102
rect 286142 442046 286238 442102
rect 285618 441978 286238 442046
rect 285618 441922 285714 441978
rect 285770 441922 285838 441978
rect 285894 441922 285962 441978
rect 286018 441922 286086 441978
rect 286142 441922 286238 441978
rect 285618 424350 286238 441922
rect 285618 424294 285714 424350
rect 285770 424294 285838 424350
rect 285894 424294 285962 424350
rect 286018 424294 286086 424350
rect 286142 424294 286238 424350
rect 285618 424226 286238 424294
rect 285618 424170 285714 424226
rect 285770 424170 285838 424226
rect 285894 424170 285962 424226
rect 286018 424170 286086 424226
rect 286142 424170 286238 424226
rect 285618 424102 286238 424170
rect 285618 424046 285714 424102
rect 285770 424046 285838 424102
rect 285894 424046 285962 424102
rect 286018 424046 286086 424102
rect 286142 424046 286238 424102
rect 285618 423978 286238 424046
rect 285618 423922 285714 423978
rect 285770 423922 285838 423978
rect 285894 423922 285962 423978
rect 286018 423922 286086 423978
rect 286142 423922 286238 423978
rect 285618 406350 286238 423922
rect 285618 406294 285714 406350
rect 285770 406294 285838 406350
rect 285894 406294 285962 406350
rect 286018 406294 286086 406350
rect 286142 406294 286238 406350
rect 285618 406226 286238 406294
rect 285618 406170 285714 406226
rect 285770 406170 285838 406226
rect 285894 406170 285962 406226
rect 286018 406170 286086 406226
rect 286142 406170 286238 406226
rect 285618 406102 286238 406170
rect 285618 406046 285714 406102
rect 285770 406046 285838 406102
rect 285894 406046 285962 406102
rect 286018 406046 286086 406102
rect 286142 406046 286238 406102
rect 285618 405978 286238 406046
rect 285618 405922 285714 405978
rect 285770 405922 285838 405978
rect 285894 405922 285962 405978
rect 286018 405922 286086 405978
rect 286142 405922 286238 405978
rect 285618 388350 286238 405922
rect 285618 388294 285714 388350
rect 285770 388294 285838 388350
rect 285894 388294 285962 388350
rect 286018 388294 286086 388350
rect 286142 388294 286238 388350
rect 285618 388226 286238 388294
rect 285618 388170 285714 388226
rect 285770 388170 285838 388226
rect 285894 388170 285962 388226
rect 286018 388170 286086 388226
rect 286142 388170 286238 388226
rect 285618 388102 286238 388170
rect 285618 388046 285714 388102
rect 285770 388046 285838 388102
rect 285894 388046 285962 388102
rect 286018 388046 286086 388102
rect 286142 388046 286238 388102
rect 285618 387978 286238 388046
rect 285618 387922 285714 387978
rect 285770 387922 285838 387978
rect 285894 387922 285962 387978
rect 286018 387922 286086 387978
rect 286142 387922 286238 387978
rect 285618 370350 286238 387922
rect 285618 370294 285714 370350
rect 285770 370294 285838 370350
rect 285894 370294 285962 370350
rect 286018 370294 286086 370350
rect 286142 370294 286238 370350
rect 285618 370226 286238 370294
rect 285618 370170 285714 370226
rect 285770 370170 285838 370226
rect 285894 370170 285962 370226
rect 286018 370170 286086 370226
rect 286142 370170 286238 370226
rect 285618 370102 286238 370170
rect 285618 370046 285714 370102
rect 285770 370046 285838 370102
rect 285894 370046 285962 370102
rect 286018 370046 286086 370102
rect 286142 370046 286238 370102
rect 285618 369978 286238 370046
rect 285618 369922 285714 369978
rect 285770 369922 285838 369978
rect 285894 369922 285962 369978
rect 286018 369922 286086 369978
rect 286142 369922 286238 369978
rect 285618 352350 286238 369922
rect 285618 352294 285714 352350
rect 285770 352294 285838 352350
rect 285894 352294 285962 352350
rect 286018 352294 286086 352350
rect 286142 352294 286238 352350
rect 285618 352226 286238 352294
rect 285618 352170 285714 352226
rect 285770 352170 285838 352226
rect 285894 352170 285962 352226
rect 286018 352170 286086 352226
rect 286142 352170 286238 352226
rect 285618 352102 286238 352170
rect 285618 352046 285714 352102
rect 285770 352046 285838 352102
rect 285894 352046 285962 352102
rect 286018 352046 286086 352102
rect 286142 352046 286238 352102
rect 285618 351978 286238 352046
rect 285618 351922 285714 351978
rect 285770 351922 285838 351978
rect 285894 351922 285962 351978
rect 286018 351922 286086 351978
rect 286142 351922 286238 351978
rect 285618 334350 286238 351922
rect 285618 334294 285714 334350
rect 285770 334294 285838 334350
rect 285894 334294 285962 334350
rect 286018 334294 286086 334350
rect 286142 334294 286238 334350
rect 285618 334226 286238 334294
rect 285618 334170 285714 334226
rect 285770 334170 285838 334226
rect 285894 334170 285962 334226
rect 286018 334170 286086 334226
rect 286142 334170 286238 334226
rect 285618 334102 286238 334170
rect 285618 334046 285714 334102
rect 285770 334046 285838 334102
rect 285894 334046 285962 334102
rect 286018 334046 286086 334102
rect 286142 334046 286238 334102
rect 285618 333978 286238 334046
rect 285618 333922 285714 333978
rect 285770 333922 285838 333978
rect 285894 333922 285962 333978
rect 286018 333922 286086 333978
rect 286142 333922 286238 333978
rect 285618 316350 286238 333922
rect 285618 316294 285714 316350
rect 285770 316294 285838 316350
rect 285894 316294 285962 316350
rect 286018 316294 286086 316350
rect 286142 316294 286238 316350
rect 285618 316226 286238 316294
rect 285618 316170 285714 316226
rect 285770 316170 285838 316226
rect 285894 316170 285962 316226
rect 286018 316170 286086 316226
rect 286142 316170 286238 316226
rect 285618 316102 286238 316170
rect 285618 316046 285714 316102
rect 285770 316046 285838 316102
rect 285894 316046 285962 316102
rect 286018 316046 286086 316102
rect 286142 316046 286238 316102
rect 285618 315978 286238 316046
rect 285618 315922 285714 315978
rect 285770 315922 285838 315978
rect 285894 315922 285962 315978
rect 286018 315922 286086 315978
rect 286142 315922 286238 315978
rect 285618 298350 286238 315922
rect 285618 298294 285714 298350
rect 285770 298294 285838 298350
rect 285894 298294 285962 298350
rect 286018 298294 286086 298350
rect 286142 298294 286238 298350
rect 285618 298226 286238 298294
rect 285618 298170 285714 298226
rect 285770 298170 285838 298226
rect 285894 298170 285962 298226
rect 286018 298170 286086 298226
rect 286142 298170 286238 298226
rect 285618 298102 286238 298170
rect 285618 298046 285714 298102
rect 285770 298046 285838 298102
rect 285894 298046 285962 298102
rect 286018 298046 286086 298102
rect 286142 298046 286238 298102
rect 285618 297978 286238 298046
rect 285618 297922 285714 297978
rect 285770 297922 285838 297978
rect 285894 297922 285962 297978
rect 286018 297922 286086 297978
rect 286142 297922 286238 297978
rect 285618 280350 286238 297922
rect 285618 280294 285714 280350
rect 285770 280294 285838 280350
rect 285894 280294 285962 280350
rect 286018 280294 286086 280350
rect 286142 280294 286238 280350
rect 285618 280226 286238 280294
rect 285618 280170 285714 280226
rect 285770 280170 285838 280226
rect 285894 280170 285962 280226
rect 286018 280170 286086 280226
rect 286142 280170 286238 280226
rect 285618 280102 286238 280170
rect 285618 280046 285714 280102
rect 285770 280046 285838 280102
rect 285894 280046 285962 280102
rect 286018 280046 286086 280102
rect 286142 280046 286238 280102
rect 285618 279978 286238 280046
rect 285618 279922 285714 279978
rect 285770 279922 285838 279978
rect 285894 279922 285962 279978
rect 286018 279922 286086 279978
rect 286142 279922 286238 279978
rect 285618 262350 286238 279922
rect 285618 262294 285714 262350
rect 285770 262294 285838 262350
rect 285894 262294 285962 262350
rect 286018 262294 286086 262350
rect 286142 262294 286238 262350
rect 285618 262226 286238 262294
rect 285618 262170 285714 262226
rect 285770 262170 285838 262226
rect 285894 262170 285962 262226
rect 286018 262170 286086 262226
rect 286142 262170 286238 262226
rect 285618 262102 286238 262170
rect 285618 262046 285714 262102
rect 285770 262046 285838 262102
rect 285894 262046 285962 262102
rect 286018 262046 286086 262102
rect 286142 262046 286238 262102
rect 285618 261978 286238 262046
rect 285618 261922 285714 261978
rect 285770 261922 285838 261978
rect 285894 261922 285962 261978
rect 286018 261922 286086 261978
rect 286142 261922 286238 261978
rect 285618 244350 286238 261922
rect 285618 244294 285714 244350
rect 285770 244294 285838 244350
rect 285894 244294 285962 244350
rect 286018 244294 286086 244350
rect 286142 244294 286238 244350
rect 285618 244226 286238 244294
rect 285618 244170 285714 244226
rect 285770 244170 285838 244226
rect 285894 244170 285962 244226
rect 286018 244170 286086 244226
rect 286142 244170 286238 244226
rect 285618 244102 286238 244170
rect 285618 244046 285714 244102
rect 285770 244046 285838 244102
rect 285894 244046 285962 244102
rect 286018 244046 286086 244102
rect 286142 244046 286238 244102
rect 285618 243978 286238 244046
rect 285618 243922 285714 243978
rect 285770 243922 285838 243978
rect 285894 243922 285962 243978
rect 286018 243922 286086 243978
rect 286142 243922 286238 243978
rect 285618 226350 286238 243922
rect 285618 226294 285714 226350
rect 285770 226294 285838 226350
rect 285894 226294 285962 226350
rect 286018 226294 286086 226350
rect 286142 226294 286238 226350
rect 285618 226226 286238 226294
rect 285618 226170 285714 226226
rect 285770 226170 285838 226226
rect 285894 226170 285962 226226
rect 286018 226170 286086 226226
rect 286142 226170 286238 226226
rect 285618 226102 286238 226170
rect 285618 226046 285714 226102
rect 285770 226046 285838 226102
rect 285894 226046 285962 226102
rect 286018 226046 286086 226102
rect 286142 226046 286238 226102
rect 285618 225978 286238 226046
rect 285618 225922 285714 225978
rect 285770 225922 285838 225978
rect 285894 225922 285962 225978
rect 286018 225922 286086 225978
rect 286142 225922 286238 225978
rect 285618 208350 286238 225922
rect 285618 208294 285714 208350
rect 285770 208294 285838 208350
rect 285894 208294 285962 208350
rect 286018 208294 286086 208350
rect 286142 208294 286238 208350
rect 285618 208226 286238 208294
rect 285618 208170 285714 208226
rect 285770 208170 285838 208226
rect 285894 208170 285962 208226
rect 286018 208170 286086 208226
rect 286142 208170 286238 208226
rect 285618 208102 286238 208170
rect 285618 208046 285714 208102
rect 285770 208046 285838 208102
rect 285894 208046 285962 208102
rect 286018 208046 286086 208102
rect 286142 208046 286238 208102
rect 285618 207978 286238 208046
rect 285618 207922 285714 207978
rect 285770 207922 285838 207978
rect 285894 207922 285962 207978
rect 286018 207922 286086 207978
rect 286142 207922 286238 207978
rect 285618 190350 286238 207922
rect 285618 190294 285714 190350
rect 285770 190294 285838 190350
rect 285894 190294 285962 190350
rect 286018 190294 286086 190350
rect 286142 190294 286238 190350
rect 285618 190226 286238 190294
rect 285618 190170 285714 190226
rect 285770 190170 285838 190226
rect 285894 190170 285962 190226
rect 286018 190170 286086 190226
rect 286142 190170 286238 190226
rect 285618 190102 286238 190170
rect 285618 190046 285714 190102
rect 285770 190046 285838 190102
rect 285894 190046 285962 190102
rect 286018 190046 286086 190102
rect 286142 190046 286238 190102
rect 285618 189978 286238 190046
rect 285618 189922 285714 189978
rect 285770 189922 285838 189978
rect 285894 189922 285962 189978
rect 286018 189922 286086 189978
rect 286142 189922 286238 189978
rect 285618 172350 286238 189922
rect 285618 172294 285714 172350
rect 285770 172294 285838 172350
rect 285894 172294 285962 172350
rect 286018 172294 286086 172350
rect 286142 172294 286238 172350
rect 285618 172226 286238 172294
rect 285618 172170 285714 172226
rect 285770 172170 285838 172226
rect 285894 172170 285962 172226
rect 286018 172170 286086 172226
rect 286142 172170 286238 172226
rect 285618 172102 286238 172170
rect 285618 172046 285714 172102
rect 285770 172046 285838 172102
rect 285894 172046 285962 172102
rect 286018 172046 286086 172102
rect 286142 172046 286238 172102
rect 285618 171978 286238 172046
rect 285618 171922 285714 171978
rect 285770 171922 285838 171978
rect 285894 171922 285962 171978
rect 286018 171922 286086 171978
rect 286142 171922 286238 171978
rect 285618 154350 286238 171922
rect 285618 154294 285714 154350
rect 285770 154294 285838 154350
rect 285894 154294 285962 154350
rect 286018 154294 286086 154350
rect 286142 154294 286238 154350
rect 285618 154226 286238 154294
rect 285618 154170 285714 154226
rect 285770 154170 285838 154226
rect 285894 154170 285962 154226
rect 286018 154170 286086 154226
rect 286142 154170 286238 154226
rect 285618 154102 286238 154170
rect 285618 154046 285714 154102
rect 285770 154046 285838 154102
rect 285894 154046 285962 154102
rect 286018 154046 286086 154102
rect 286142 154046 286238 154102
rect 285618 153978 286238 154046
rect 285618 153922 285714 153978
rect 285770 153922 285838 153978
rect 285894 153922 285962 153978
rect 286018 153922 286086 153978
rect 286142 153922 286238 153978
rect 285618 136350 286238 153922
rect 285618 136294 285714 136350
rect 285770 136294 285838 136350
rect 285894 136294 285962 136350
rect 286018 136294 286086 136350
rect 286142 136294 286238 136350
rect 285618 136226 286238 136294
rect 285618 136170 285714 136226
rect 285770 136170 285838 136226
rect 285894 136170 285962 136226
rect 286018 136170 286086 136226
rect 286142 136170 286238 136226
rect 285618 136102 286238 136170
rect 285618 136046 285714 136102
rect 285770 136046 285838 136102
rect 285894 136046 285962 136102
rect 286018 136046 286086 136102
rect 286142 136046 286238 136102
rect 285618 135978 286238 136046
rect 285618 135922 285714 135978
rect 285770 135922 285838 135978
rect 285894 135922 285962 135978
rect 286018 135922 286086 135978
rect 286142 135922 286238 135978
rect 285618 118350 286238 135922
rect 285618 118294 285714 118350
rect 285770 118294 285838 118350
rect 285894 118294 285962 118350
rect 286018 118294 286086 118350
rect 286142 118294 286238 118350
rect 285618 118226 286238 118294
rect 285618 118170 285714 118226
rect 285770 118170 285838 118226
rect 285894 118170 285962 118226
rect 286018 118170 286086 118226
rect 286142 118170 286238 118226
rect 285618 118102 286238 118170
rect 285618 118046 285714 118102
rect 285770 118046 285838 118102
rect 285894 118046 285962 118102
rect 286018 118046 286086 118102
rect 286142 118046 286238 118102
rect 285618 117978 286238 118046
rect 285618 117922 285714 117978
rect 285770 117922 285838 117978
rect 285894 117922 285962 117978
rect 286018 117922 286086 117978
rect 286142 117922 286238 117978
rect 285618 100350 286238 117922
rect 285618 100294 285714 100350
rect 285770 100294 285838 100350
rect 285894 100294 285962 100350
rect 286018 100294 286086 100350
rect 286142 100294 286238 100350
rect 285618 100226 286238 100294
rect 285618 100170 285714 100226
rect 285770 100170 285838 100226
rect 285894 100170 285962 100226
rect 286018 100170 286086 100226
rect 286142 100170 286238 100226
rect 285618 100102 286238 100170
rect 285618 100046 285714 100102
rect 285770 100046 285838 100102
rect 285894 100046 285962 100102
rect 286018 100046 286086 100102
rect 286142 100046 286238 100102
rect 285618 99978 286238 100046
rect 285618 99922 285714 99978
rect 285770 99922 285838 99978
rect 285894 99922 285962 99978
rect 286018 99922 286086 99978
rect 286142 99922 286238 99978
rect 285618 82350 286238 99922
rect 285618 82294 285714 82350
rect 285770 82294 285838 82350
rect 285894 82294 285962 82350
rect 286018 82294 286086 82350
rect 286142 82294 286238 82350
rect 285618 82226 286238 82294
rect 285618 82170 285714 82226
rect 285770 82170 285838 82226
rect 285894 82170 285962 82226
rect 286018 82170 286086 82226
rect 286142 82170 286238 82226
rect 285618 82102 286238 82170
rect 285618 82046 285714 82102
rect 285770 82046 285838 82102
rect 285894 82046 285962 82102
rect 286018 82046 286086 82102
rect 286142 82046 286238 82102
rect 285618 81978 286238 82046
rect 285618 81922 285714 81978
rect 285770 81922 285838 81978
rect 285894 81922 285962 81978
rect 286018 81922 286086 81978
rect 286142 81922 286238 81978
rect 285618 64350 286238 81922
rect 297388 590212 297444 590222
rect 297388 78238 297444 590156
rect 297388 78172 297444 78182
rect 312618 580350 313238 596784
rect 312618 580294 312714 580350
rect 312770 580294 312838 580350
rect 312894 580294 312962 580350
rect 313018 580294 313086 580350
rect 313142 580294 313238 580350
rect 312618 580226 313238 580294
rect 312618 580170 312714 580226
rect 312770 580170 312838 580226
rect 312894 580170 312962 580226
rect 313018 580170 313086 580226
rect 313142 580170 313238 580226
rect 312618 580102 313238 580170
rect 312618 580046 312714 580102
rect 312770 580046 312838 580102
rect 312894 580046 312962 580102
rect 313018 580046 313086 580102
rect 313142 580046 313238 580102
rect 312618 579978 313238 580046
rect 312618 579922 312714 579978
rect 312770 579922 312838 579978
rect 312894 579922 312962 579978
rect 313018 579922 313086 579978
rect 313142 579922 313238 579978
rect 312618 562350 313238 579922
rect 312618 562294 312714 562350
rect 312770 562294 312838 562350
rect 312894 562294 312962 562350
rect 313018 562294 313086 562350
rect 313142 562294 313238 562350
rect 312618 562226 313238 562294
rect 312618 562170 312714 562226
rect 312770 562170 312838 562226
rect 312894 562170 312962 562226
rect 313018 562170 313086 562226
rect 313142 562170 313238 562226
rect 312618 562102 313238 562170
rect 312618 562046 312714 562102
rect 312770 562046 312838 562102
rect 312894 562046 312962 562102
rect 313018 562046 313086 562102
rect 313142 562046 313238 562102
rect 312618 561978 313238 562046
rect 312618 561922 312714 561978
rect 312770 561922 312838 561978
rect 312894 561922 312962 561978
rect 313018 561922 313086 561978
rect 313142 561922 313238 561978
rect 312618 544350 313238 561922
rect 312618 544294 312714 544350
rect 312770 544294 312838 544350
rect 312894 544294 312962 544350
rect 313018 544294 313086 544350
rect 313142 544294 313238 544350
rect 312618 544226 313238 544294
rect 312618 544170 312714 544226
rect 312770 544170 312838 544226
rect 312894 544170 312962 544226
rect 313018 544170 313086 544226
rect 313142 544170 313238 544226
rect 312618 544102 313238 544170
rect 312618 544046 312714 544102
rect 312770 544046 312838 544102
rect 312894 544046 312962 544102
rect 313018 544046 313086 544102
rect 313142 544046 313238 544102
rect 312618 543978 313238 544046
rect 312618 543922 312714 543978
rect 312770 543922 312838 543978
rect 312894 543922 312962 543978
rect 313018 543922 313086 543978
rect 313142 543922 313238 543978
rect 312618 526350 313238 543922
rect 312618 526294 312714 526350
rect 312770 526294 312838 526350
rect 312894 526294 312962 526350
rect 313018 526294 313086 526350
rect 313142 526294 313238 526350
rect 312618 526226 313238 526294
rect 312618 526170 312714 526226
rect 312770 526170 312838 526226
rect 312894 526170 312962 526226
rect 313018 526170 313086 526226
rect 313142 526170 313238 526226
rect 312618 526102 313238 526170
rect 312618 526046 312714 526102
rect 312770 526046 312838 526102
rect 312894 526046 312962 526102
rect 313018 526046 313086 526102
rect 313142 526046 313238 526102
rect 312618 525978 313238 526046
rect 312618 525922 312714 525978
rect 312770 525922 312838 525978
rect 312894 525922 312962 525978
rect 313018 525922 313086 525978
rect 313142 525922 313238 525978
rect 312618 508350 313238 525922
rect 312618 508294 312714 508350
rect 312770 508294 312838 508350
rect 312894 508294 312962 508350
rect 313018 508294 313086 508350
rect 313142 508294 313238 508350
rect 312618 508226 313238 508294
rect 312618 508170 312714 508226
rect 312770 508170 312838 508226
rect 312894 508170 312962 508226
rect 313018 508170 313086 508226
rect 313142 508170 313238 508226
rect 312618 508102 313238 508170
rect 312618 508046 312714 508102
rect 312770 508046 312838 508102
rect 312894 508046 312962 508102
rect 313018 508046 313086 508102
rect 313142 508046 313238 508102
rect 312618 507978 313238 508046
rect 312618 507922 312714 507978
rect 312770 507922 312838 507978
rect 312894 507922 312962 507978
rect 313018 507922 313086 507978
rect 313142 507922 313238 507978
rect 312618 490350 313238 507922
rect 312618 490294 312714 490350
rect 312770 490294 312838 490350
rect 312894 490294 312962 490350
rect 313018 490294 313086 490350
rect 313142 490294 313238 490350
rect 312618 490226 313238 490294
rect 312618 490170 312714 490226
rect 312770 490170 312838 490226
rect 312894 490170 312962 490226
rect 313018 490170 313086 490226
rect 313142 490170 313238 490226
rect 312618 490102 313238 490170
rect 312618 490046 312714 490102
rect 312770 490046 312838 490102
rect 312894 490046 312962 490102
rect 313018 490046 313086 490102
rect 313142 490046 313238 490102
rect 312618 489978 313238 490046
rect 312618 489922 312714 489978
rect 312770 489922 312838 489978
rect 312894 489922 312962 489978
rect 313018 489922 313086 489978
rect 313142 489922 313238 489978
rect 312618 472350 313238 489922
rect 312618 472294 312714 472350
rect 312770 472294 312838 472350
rect 312894 472294 312962 472350
rect 313018 472294 313086 472350
rect 313142 472294 313238 472350
rect 312618 472226 313238 472294
rect 312618 472170 312714 472226
rect 312770 472170 312838 472226
rect 312894 472170 312962 472226
rect 313018 472170 313086 472226
rect 313142 472170 313238 472226
rect 312618 472102 313238 472170
rect 312618 472046 312714 472102
rect 312770 472046 312838 472102
rect 312894 472046 312962 472102
rect 313018 472046 313086 472102
rect 313142 472046 313238 472102
rect 312618 471978 313238 472046
rect 312618 471922 312714 471978
rect 312770 471922 312838 471978
rect 312894 471922 312962 471978
rect 313018 471922 313086 471978
rect 313142 471922 313238 471978
rect 312618 454350 313238 471922
rect 312618 454294 312714 454350
rect 312770 454294 312838 454350
rect 312894 454294 312962 454350
rect 313018 454294 313086 454350
rect 313142 454294 313238 454350
rect 312618 454226 313238 454294
rect 312618 454170 312714 454226
rect 312770 454170 312838 454226
rect 312894 454170 312962 454226
rect 313018 454170 313086 454226
rect 313142 454170 313238 454226
rect 312618 454102 313238 454170
rect 312618 454046 312714 454102
rect 312770 454046 312838 454102
rect 312894 454046 312962 454102
rect 313018 454046 313086 454102
rect 313142 454046 313238 454102
rect 312618 453978 313238 454046
rect 312618 453922 312714 453978
rect 312770 453922 312838 453978
rect 312894 453922 312962 453978
rect 313018 453922 313086 453978
rect 313142 453922 313238 453978
rect 312618 436350 313238 453922
rect 312618 436294 312714 436350
rect 312770 436294 312838 436350
rect 312894 436294 312962 436350
rect 313018 436294 313086 436350
rect 313142 436294 313238 436350
rect 312618 436226 313238 436294
rect 312618 436170 312714 436226
rect 312770 436170 312838 436226
rect 312894 436170 312962 436226
rect 313018 436170 313086 436226
rect 313142 436170 313238 436226
rect 312618 436102 313238 436170
rect 312618 436046 312714 436102
rect 312770 436046 312838 436102
rect 312894 436046 312962 436102
rect 313018 436046 313086 436102
rect 313142 436046 313238 436102
rect 312618 435978 313238 436046
rect 312618 435922 312714 435978
rect 312770 435922 312838 435978
rect 312894 435922 312962 435978
rect 313018 435922 313086 435978
rect 313142 435922 313238 435978
rect 312618 418350 313238 435922
rect 312618 418294 312714 418350
rect 312770 418294 312838 418350
rect 312894 418294 312962 418350
rect 313018 418294 313086 418350
rect 313142 418294 313238 418350
rect 312618 418226 313238 418294
rect 312618 418170 312714 418226
rect 312770 418170 312838 418226
rect 312894 418170 312962 418226
rect 313018 418170 313086 418226
rect 313142 418170 313238 418226
rect 312618 418102 313238 418170
rect 312618 418046 312714 418102
rect 312770 418046 312838 418102
rect 312894 418046 312962 418102
rect 313018 418046 313086 418102
rect 313142 418046 313238 418102
rect 312618 417978 313238 418046
rect 312618 417922 312714 417978
rect 312770 417922 312838 417978
rect 312894 417922 312962 417978
rect 313018 417922 313086 417978
rect 313142 417922 313238 417978
rect 312618 400350 313238 417922
rect 312618 400294 312714 400350
rect 312770 400294 312838 400350
rect 312894 400294 312962 400350
rect 313018 400294 313086 400350
rect 313142 400294 313238 400350
rect 312618 400226 313238 400294
rect 312618 400170 312714 400226
rect 312770 400170 312838 400226
rect 312894 400170 312962 400226
rect 313018 400170 313086 400226
rect 313142 400170 313238 400226
rect 312618 400102 313238 400170
rect 312618 400046 312714 400102
rect 312770 400046 312838 400102
rect 312894 400046 312962 400102
rect 313018 400046 313086 400102
rect 313142 400046 313238 400102
rect 312618 399978 313238 400046
rect 312618 399922 312714 399978
rect 312770 399922 312838 399978
rect 312894 399922 312962 399978
rect 313018 399922 313086 399978
rect 313142 399922 313238 399978
rect 312618 382350 313238 399922
rect 312618 382294 312714 382350
rect 312770 382294 312838 382350
rect 312894 382294 312962 382350
rect 313018 382294 313086 382350
rect 313142 382294 313238 382350
rect 312618 382226 313238 382294
rect 312618 382170 312714 382226
rect 312770 382170 312838 382226
rect 312894 382170 312962 382226
rect 313018 382170 313086 382226
rect 313142 382170 313238 382226
rect 312618 382102 313238 382170
rect 312618 382046 312714 382102
rect 312770 382046 312838 382102
rect 312894 382046 312962 382102
rect 313018 382046 313086 382102
rect 313142 382046 313238 382102
rect 312618 381978 313238 382046
rect 312618 381922 312714 381978
rect 312770 381922 312838 381978
rect 312894 381922 312962 381978
rect 313018 381922 313086 381978
rect 313142 381922 313238 381978
rect 312618 364350 313238 381922
rect 312618 364294 312714 364350
rect 312770 364294 312838 364350
rect 312894 364294 312962 364350
rect 313018 364294 313086 364350
rect 313142 364294 313238 364350
rect 312618 364226 313238 364294
rect 312618 364170 312714 364226
rect 312770 364170 312838 364226
rect 312894 364170 312962 364226
rect 313018 364170 313086 364226
rect 313142 364170 313238 364226
rect 312618 364102 313238 364170
rect 312618 364046 312714 364102
rect 312770 364046 312838 364102
rect 312894 364046 312962 364102
rect 313018 364046 313086 364102
rect 313142 364046 313238 364102
rect 312618 363978 313238 364046
rect 312618 363922 312714 363978
rect 312770 363922 312838 363978
rect 312894 363922 312962 363978
rect 313018 363922 313086 363978
rect 313142 363922 313238 363978
rect 312618 346350 313238 363922
rect 312618 346294 312714 346350
rect 312770 346294 312838 346350
rect 312894 346294 312962 346350
rect 313018 346294 313086 346350
rect 313142 346294 313238 346350
rect 312618 346226 313238 346294
rect 312618 346170 312714 346226
rect 312770 346170 312838 346226
rect 312894 346170 312962 346226
rect 313018 346170 313086 346226
rect 313142 346170 313238 346226
rect 312618 346102 313238 346170
rect 312618 346046 312714 346102
rect 312770 346046 312838 346102
rect 312894 346046 312962 346102
rect 313018 346046 313086 346102
rect 313142 346046 313238 346102
rect 312618 345978 313238 346046
rect 312618 345922 312714 345978
rect 312770 345922 312838 345978
rect 312894 345922 312962 345978
rect 313018 345922 313086 345978
rect 313142 345922 313238 345978
rect 312618 328350 313238 345922
rect 312618 328294 312714 328350
rect 312770 328294 312838 328350
rect 312894 328294 312962 328350
rect 313018 328294 313086 328350
rect 313142 328294 313238 328350
rect 312618 328226 313238 328294
rect 312618 328170 312714 328226
rect 312770 328170 312838 328226
rect 312894 328170 312962 328226
rect 313018 328170 313086 328226
rect 313142 328170 313238 328226
rect 312618 328102 313238 328170
rect 312618 328046 312714 328102
rect 312770 328046 312838 328102
rect 312894 328046 312962 328102
rect 313018 328046 313086 328102
rect 313142 328046 313238 328102
rect 312618 327978 313238 328046
rect 312618 327922 312714 327978
rect 312770 327922 312838 327978
rect 312894 327922 312962 327978
rect 313018 327922 313086 327978
rect 313142 327922 313238 327978
rect 312618 310350 313238 327922
rect 312618 310294 312714 310350
rect 312770 310294 312838 310350
rect 312894 310294 312962 310350
rect 313018 310294 313086 310350
rect 313142 310294 313238 310350
rect 312618 310226 313238 310294
rect 312618 310170 312714 310226
rect 312770 310170 312838 310226
rect 312894 310170 312962 310226
rect 313018 310170 313086 310226
rect 313142 310170 313238 310226
rect 312618 310102 313238 310170
rect 312618 310046 312714 310102
rect 312770 310046 312838 310102
rect 312894 310046 312962 310102
rect 313018 310046 313086 310102
rect 313142 310046 313238 310102
rect 312618 309978 313238 310046
rect 312618 309922 312714 309978
rect 312770 309922 312838 309978
rect 312894 309922 312962 309978
rect 313018 309922 313086 309978
rect 313142 309922 313238 309978
rect 312618 292350 313238 309922
rect 312618 292294 312714 292350
rect 312770 292294 312838 292350
rect 312894 292294 312962 292350
rect 313018 292294 313086 292350
rect 313142 292294 313238 292350
rect 312618 292226 313238 292294
rect 312618 292170 312714 292226
rect 312770 292170 312838 292226
rect 312894 292170 312962 292226
rect 313018 292170 313086 292226
rect 313142 292170 313238 292226
rect 312618 292102 313238 292170
rect 312618 292046 312714 292102
rect 312770 292046 312838 292102
rect 312894 292046 312962 292102
rect 313018 292046 313086 292102
rect 313142 292046 313238 292102
rect 312618 291978 313238 292046
rect 312618 291922 312714 291978
rect 312770 291922 312838 291978
rect 312894 291922 312962 291978
rect 313018 291922 313086 291978
rect 313142 291922 313238 291978
rect 312618 274350 313238 291922
rect 312618 274294 312714 274350
rect 312770 274294 312838 274350
rect 312894 274294 312962 274350
rect 313018 274294 313086 274350
rect 313142 274294 313238 274350
rect 312618 274226 313238 274294
rect 312618 274170 312714 274226
rect 312770 274170 312838 274226
rect 312894 274170 312962 274226
rect 313018 274170 313086 274226
rect 313142 274170 313238 274226
rect 312618 274102 313238 274170
rect 312618 274046 312714 274102
rect 312770 274046 312838 274102
rect 312894 274046 312962 274102
rect 313018 274046 313086 274102
rect 313142 274046 313238 274102
rect 312618 273978 313238 274046
rect 312618 273922 312714 273978
rect 312770 273922 312838 273978
rect 312894 273922 312962 273978
rect 313018 273922 313086 273978
rect 313142 273922 313238 273978
rect 312618 256350 313238 273922
rect 312618 256294 312714 256350
rect 312770 256294 312838 256350
rect 312894 256294 312962 256350
rect 313018 256294 313086 256350
rect 313142 256294 313238 256350
rect 312618 256226 313238 256294
rect 312618 256170 312714 256226
rect 312770 256170 312838 256226
rect 312894 256170 312962 256226
rect 313018 256170 313086 256226
rect 313142 256170 313238 256226
rect 312618 256102 313238 256170
rect 312618 256046 312714 256102
rect 312770 256046 312838 256102
rect 312894 256046 312962 256102
rect 313018 256046 313086 256102
rect 313142 256046 313238 256102
rect 312618 255978 313238 256046
rect 312618 255922 312714 255978
rect 312770 255922 312838 255978
rect 312894 255922 312962 255978
rect 313018 255922 313086 255978
rect 313142 255922 313238 255978
rect 312618 238350 313238 255922
rect 312618 238294 312714 238350
rect 312770 238294 312838 238350
rect 312894 238294 312962 238350
rect 313018 238294 313086 238350
rect 313142 238294 313238 238350
rect 312618 238226 313238 238294
rect 312618 238170 312714 238226
rect 312770 238170 312838 238226
rect 312894 238170 312962 238226
rect 313018 238170 313086 238226
rect 313142 238170 313238 238226
rect 312618 238102 313238 238170
rect 312618 238046 312714 238102
rect 312770 238046 312838 238102
rect 312894 238046 312962 238102
rect 313018 238046 313086 238102
rect 313142 238046 313238 238102
rect 312618 237978 313238 238046
rect 312618 237922 312714 237978
rect 312770 237922 312838 237978
rect 312894 237922 312962 237978
rect 313018 237922 313086 237978
rect 313142 237922 313238 237978
rect 312618 220350 313238 237922
rect 312618 220294 312714 220350
rect 312770 220294 312838 220350
rect 312894 220294 312962 220350
rect 313018 220294 313086 220350
rect 313142 220294 313238 220350
rect 312618 220226 313238 220294
rect 312618 220170 312714 220226
rect 312770 220170 312838 220226
rect 312894 220170 312962 220226
rect 313018 220170 313086 220226
rect 313142 220170 313238 220226
rect 312618 220102 313238 220170
rect 312618 220046 312714 220102
rect 312770 220046 312838 220102
rect 312894 220046 312962 220102
rect 313018 220046 313086 220102
rect 313142 220046 313238 220102
rect 312618 219978 313238 220046
rect 312618 219922 312714 219978
rect 312770 219922 312838 219978
rect 312894 219922 312962 219978
rect 313018 219922 313086 219978
rect 313142 219922 313238 219978
rect 312618 202350 313238 219922
rect 312618 202294 312714 202350
rect 312770 202294 312838 202350
rect 312894 202294 312962 202350
rect 313018 202294 313086 202350
rect 313142 202294 313238 202350
rect 312618 202226 313238 202294
rect 312618 202170 312714 202226
rect 312770 202170 312838 202226
rect 312894 202170 312962 202226
rect 313018 202170 313086 202226
rect 313142 202170 313238 202226
rect 312618 202102 313238 202170
rect 312618 202046 312714 202102
rect 312770 202046 312838 202102
rect 312894 202046 312962 202102
rect 313018 202046 313086 202102
rect 313142 202046 313238 202102
rect 312618 201978 313238 202046
rect 312618 201922 312714 201978
rect 312770 201922 312838 201978
rect 312894 201922 312962 201978
rect 313018 201922 313086 201978
rect 313142 201922 313238 201978
rect 312618 184350 313238 201922
rect 312618 184294 312714 184350
rect 312770 184294 312838 184350
rect 312894 184294 312962 184350
rect 313018 184294 313086 184350
rect 313142 184294 313238 184350
rect 312618 184226 313238 184294
rect 312618 184170 312714 184226
rect 312770 184170 312838 184226
rect 312894 184170 312962 184226
rect 313018 184170 313086 184226
rect 313142 184170 313238 184226
rect 312618 184102 313238 184170
rect 312618 184046 312714 184102
rect 312770 184046 312838 184102
rect 312894 184046 312962 184102
rect 313018 184046 313086 184102
rect 313142 184046 313238 184102
rect 312618 183978 313238 184046
rect 312618 183922 312714 183978
rect 312770 183922 312838 183978
rect 312894 183922 312962 183978
rect 313018 183922 313086 183978
rect 313142 183922 313238 183978
rect 312618 166350 313238 183922
rect 312618 166294 312714 166350
rect 312770 166294 312838 166350
rect 312894 166294 312962 166350
rect 313018 166294 313086 166350
rect 313142 166294 313238 166350
rect 312618 166226 313238 166294
rect 312618 166170 312714 166226
rect 312770 166170 312838 166226
rect 312894 166170 312962 166226
rect 313018 166170 313086 166226
rect 313142 166170 313238 166226
rect 312618 166102 313238 166170
rect 312618 166046 312714 166102
rect 312770 166046 312838 166102
rect 312894 166046 312962 166102
rect 313018 166046 313086 166102
rect 313142 166046 313238 166102
rect 312618 165978 313238 166046
rect 312618 165922 312714 165978
rect 312770 165922 312838 165978
rect 312894 165922 312962 165978
rect 313018 165922 313086 165978
rect 313142 165922 313238 165978
rect 312618 148350 313238 165922
rect 312618 148294 312714 148350
rect 312770 148294 312838 148350
rect 312894 148294 312962 148350
rect 313018 148294 313086 148350
rect 313142 148294 313238 148350
rect 312618 148226 313238 148294
rect 312618 148170 312714 148226
rect 312770 148170 312838 148226
rect 312894 148170 312962 148226
rect 313018 148170 313086 148226
rect 313142 148170 313238 148226
rect 312618 148102 313238 148170
rect 312618 148046 312714 148102
rect 312770 148046 312838 148102
rect 312894 148046 312962 148102
rect 313018 148046 313086 148102
rect 313142 148046 313238 148102
rect 312618 147978 313238 148046
rect 312618 147922 312714 147978
rect 312770 147922 312838 147978
rect 312894 147922 312962 147978
rect 313018 147922 313086 147978
rect 313142 147922 313238 147978
rect 312618 130350 313238 147922
rect 312618 130294 312714 130350
rect 312770 130294 312838 130350
rect 312894 130294 312962 130350
rect 313018 130294 313086 130350
rect 313142 130294 313238 130350
rect 312618 130226 313238 130294
rect 312618 130170 312714 130226
rect 312770 130170 312838 130226
rect 312894 130170 312962 130226
rect 313018 130170 313086 130226
rect 313142 130170 313238 130226
rect 312618 130102 313238 130170
rect 312618 130046 312714 130102
rect 312770 130046 312838 130102
rect 312894 130046 312962 130102
rect 313018 130046 313086 130102
rect 313142 130046 313238 130102
rect 312618 129978 313238 130046
rect 312618 129922 312714 129978
rect 312770 129922 312838 129978
rect 312894 129922 312962 129978
rect 313018 129922 313086 129978
rect 313142 129922 313238 129978
rect 312618 112350 313238 129922
rect 312618 112294 312714 112350
rect 312770 112294 312838 112350
rect 312894 112294 312962 112350
rect 313018 112294 313086 112350
rect 313142 112294 313238 112350
rect 312618 112226 313238 112294
rect 312618 112170 312714 112226
rect 312770 112170 312838 112226
rect 312894 112170 312962 112226
rect 313018 112170 313086 112226
rect 313142 112170 313238 112226
rect 312618 112102 313238 112170
rect 312618 112046 312714 112102
rect 312770 112046 312838 112102
rect 312894 112046 312962 112102
rect 313018 112046 313086 112102
rect 313142 112046 313238 112102
rect 312618 111978 313238 112046
rect 312618 111922 312714 111978
rect 312770 111922 312838 111978
rect 312894 111922 312962 111978
rect 313018 111922 313086 111978
rect 313142 111922 313238 111978
rect 312618 94350 313238 111922
rect 312618 94294 312714 94350
rect 312770 94294 312838 94350
rect 312894 94294 312962 94350
rect 313018 94294 313086 94350
rect 313142 94294 313238 94350
rect 312618 94226 313238 94294
rect 312618 94170 312714 94226
rect 312770 94170 312838 94226
rect 312894 94170 312962 94226
rect 313018 94170 313086 94226
rect 313142 94170 313238 94226
rect 312618 94102 313238 94170
rect 312618 94046 312714 94102
rect 312770 94046 312838 94102
rect 312894 94046 312962 94102
rect 313018 94046 313086 94102
rect 313142 94046 313238 94102
rect 312618 93978 313238 94046
rect 312618 93922 312714 93978
rect 312770 93922 312838 93978
rect 312894 93922 312962 93978
rect 313018 93922 313086 93978
rect 313142 93922 313238 93978
rect 312618 76350 313238 93922
rect 312618 76294 312714 76350
rect 312770 76294 312838 76350
rect 312894 76294 312962 76350
rect 313018 76294 313086 76350
rect 313142 76294 313238 76350
rect 312618 76226 313238 76294
rect 312618 76170 312714 76226
rect 312770 76170 312838 76226
rect 312894 76170 312962 76226
rect 313018 76170 313086 76226
rect 313142 76170 313238 76226
rect 312618 76102 313238 76170
rect 312618 76046 312714 76102
rect 312770 76046 312838 76102
rect 312894 76046 312962 76102
rect 313018 76046 313086 76102
rect 313142 76046 313238 76102
rect 312618 75978 313238 76046
rect 312618 75922 312714 75978
rect 312770 75922 312838 75978
rect 312894 75922 312962 75978
rect 313018 75922 313086 75978
rect 313142 75922 313238 75978
rect 288988 70858 289044 70868
rect 285618 64294 285714 64350
rect 285770 64294 285838 64350
rect 285894 64294 285962 64350
rect 286018 64294 286086 64350
rect 286142 64294 286238 64350
rect 285618 64226 286238 64294
rect 285618 64170 285714 64226
rect 285770 64170 285838 64226
rect 285894 64170 285962 64226
rect 286018 64170 286086 64226
rect 286142 64170 286238 64226
rect 285618 64102 286238 64170
rect 285618 64046 285714 64102
rect 285770 64046 285838 64102
rect 285894 64046 285962 64102
rect 286018 64046 286086 64102
rect 286142 64046 286238 64102
rect 285618 63978 286238 64046
rect 285618 63922 285714 63978
rect 285770 63922 285838 63978
rect 285894 63922 285962 63978
rect 286018 63922 286086 63978
rect 286142 63922 286238 63978
rect 281898 40294 281994 40350
rect 282050 40294 282118 40350
rect 282174 40294 282242 40350
rect 282298 40294 282366 40350
rect 282422 40294 282518 40350
rect 281898 40226 282518 40294
rect 281898 40170 281994 40226
rect 282050 40170 282118 40226
rect 282174 40170 282242 40226
rect 282298 40170 282366 40226
rect 282422 40170 282518 40226
rect 281898 40102 282518 40170
rect 281898 40046 281994 40102
rect 282050 40046 282118 40102
rect 282174 40046 282242 40102
rect 282298 40046 282366 40102
rect 282422 40046 282518 40102
rect 281898 39978 282518 40046
rect 281898 39922 281994 39978
rect 282050 39922 282118 39978
rect 282174 39922 282242 39978
rect 282298 39922 282366 39978
rect 282422 39922 282518 39978
rect 278908 34318 278964 34328
rect 273868 20132 274148 20188
rect 265468 4162 265524 4172
rect 268380 5698 268436 5708
rect 257068 3490 257124 3500
rect 268380 3444 268436 5642
rect 274092 4228 274148 20132
rect 274092 4162 274148 4172
rect 278908 4228 278964 34262
rect 278908 4162 278964 4172
rect 281898 22350 282518 39922
rect 281898 22294 281994 22350
rect 282050 22294 282118 22350
rect 282174 22294 282242 22350
rect 282298 22294 282366 22350
rect 282422 22294 282518 22350
rect 281898 22226 282518 22294
rect 281898 22170 281994 22226
rect 282050 22170 282118 22226
rect 282174 22170 282242 22226
rect 282298 22170 282366 22226
rect 282422 22170 282518 22226
rect 281898 22102 282518 22170
rect 281898 22046 281994 22102
rect 282050 22046 282118 22102
rect 282174 22046 282242 22102
rect 282298 22046 282366 22102
rect 282422 22046 282518 22102
rect 281898 21978 282518 22046
rect 281898 21922 281994 21978
rect 282050 21922 282118 21978
rect 282174 21922 282242 21978
rect 282298 21922 282366 21978
rect 282422 21922 282518 21978
rect 281898 4350 282518 21922
rect 281898 4294 281994 4350
rect 282050 4294 282118 4350
rect 282174 4294 282242 4350
rect 282298 4294 282366 4350
rect 282422 4294 282518 4350
rect 281898 4226 282518 4294
rect 281898 4170 281994 4226
rect 282050 4170 282118 4226
rect 282174 4170 282242 4226
rect 282298 4170 282366 4226
rect 282422 4170 282518 4226
rect 268380 3378 268436 3388
rect 281898 4102 282518 4170
rect 282604 49618 282660 49628
rect 282604 4228 282660 49562
rect 282604 4162 282660 4172
rect 285618 46350 286238 63922
rect 285618 46294 285714 46350
rect 285770 46294 285838 46350
rect 285894 46294 285962 46350
rect 286018 46294 286086 46350
rect 286142 46294 286238 46350
rect 285618 46226 286238 46294
rect 285618 46170 285714 46226
rect 285770 46170 285838 46226
rect 285894 46170 285962 46226
rect 286018 46170 286086 46226
rect 286142 46170 286238 46226
rect 285618 46102 286238 46170
rect 285618 46046 285714 46102
rect 285770 46046 285838 46102
rect 285894 46046 285962 46102
rect 286018 46046 286086 46102
rect 286142 46046 286238 46102
rect 285618 45978 286238 46046
rect 285618 45922 285714 45978
rect 285770 45922 285838 45978
rect 285894 45922 285962 45978
rect 286018 45922 286086 45978
rect 286142 45922 286238 45978
rect 285618 28350 286238 45922
rect 285618 28294 285714 28350
rect 285770 28294 285838 28350
rect 285894 28294 285962 28350
rect 286018 28294 286086 28350
rect 286142 28294 286238 28350
rect 285618 28226 286238 28294
rect 285618 28170 285714 28226
rect 285770 28170 285838 28226
rect 285894 28170 285962 28226
rect 286018 28170 286086 28226
rect 286142 28170 286238 28226
rect 285618 28102 286238 28170
rect 285618 28046 285714 28102
rect 285770 28046 285838 28102
rect 285894 28046 285962 28102
rect 286018 28046 286086 28102
rect 286142 28046 286238 28102
rect 285618 27978 286238 28046
rect 285618 27922 285714 27978
rect 285770 27922 285838 27978
rect 285894 27922 285962 27978
rect 286018 27922 286086 27978
rect 286142 27922 286238 27978
rect 285618 10350 286238 27922
rect 285618 10294 285714 10350
rect 285770 10294 285838 10350
rect 285894 10294 285962 10350
rect 286018 10294 286086 10350
rect 286142 10294 286238 10350
rect 285618 10226 286238 10294
rect 285618 10170 285714 10226
rect 285770 10170 285838 10226
rect 285894 10170 285962 10226
rect 286018 10170 286086 10226
rect 286142 10170 286238 10226
rect 285618 10102 286238 10170
rect 285618 10046 285714 10102
rect 285770 10046 285838 10102
rect 285894 10046 285962 10102
rect 286018 10046 286086 10102
rect 286142 10046 286238 10102
rect 285618 9978 286238 10046
rect 285618 9922 285714 9978
rect 285770 9922 285838 9978
rect 285894 9922 285962 9978
rect 286018 9922 286086 9978
rect 286142 9922 286238 9978
rect 281898 4046 281994 4102
rect 282050 4046 282118 4102
rect 282174 4046 282242 4102
rect 282298 4046 282366 4102
rect 282422 4046 282518 4102
rect 281898 3978 282518 4046
rect 281898 3922 281994 3978
rect 282050 3922 282118 3978
rect 282174 3922 282242 3978
rect 282298 3922 282366 3978
rect 282422 3922 282518 3978
rect 254898 -1176 254994 -1120
rect 255050 -1176 255118 -1120
rect 255174 -1176 255242 -1120
rect 255298 -1176 255366 -1120
rect 255422 -1176 255518 -1120
rect 254898 -1244 255518 -1176
rect 254898 -1300 254994 -1244
rect 255050 -1300 255118 -1244
rect 255174 -1300 255242 -1244
rect 255298 -1300 255366 -1244
rect 255422 -1300 255518 -1244
rect 254898 -1368 255518 -1300
rect 254898 -1424 254994 -1368
rect 255050 -1424 255118 -1368
rect 255174 -1424 255242 -1368
rect 255298 -1424 255366 -1368
rect 255422 -1424 255518 -1368
rect 254898 -1492 255518 -1424
rect 254898 -1548 254994 -1492
rect 255050 -1548 255118 -1492
rect 255174 -1548 255242 -1492
rect 255298 -1548 255366 -1492
rect 255422 -1548 255518 -1492
rect 254898 -1644 255518 -1548
rect 281898 -160 282518 3922
rect 281898 -216 281994 -160
rect 282050 -216 282118 -160
rect 282174 -216 282242 -160
rect 282298 -216 282366 -160
rect 282422 -216 282518 -160
rect 281898 -284 282518 -216
rect 281898 -340 281994 -284
rect 282050 -340 282118 -284
rect 282174 -340 282242 -284
rect 282298 -340 282366 -284
rect 282422 -340 282518 -284
rect 281898 -408 282518 -340
rect 281898 -464 281994 -408
rect 282050 -464 282118 -408
rect 282174 -464 282242 -408
rect 282298 -464 282366 -408
rect 282422 -464 282518 -408
rect 281898 -532 282518 -464
rect 281898 -588 281994 -532
rect 282050 -588 282118 -532
rect 282174 -588 282242 -532
rect 282298 -588 282366 -532
rect 282422 -588 282518 -532
rect 281898 -1644 282518 -588
rect 285618 -1120 286238 9922
rect 286300 69238 286356 69248
rect 286300 4228 286356 69182
rect 286300 4162 286356 4172
rect 288988 4228 289044 70802
rect 295708 70678 295764 70688
rect 294028 67618 294084 67628
rect 288988 4162 289044 4172
rect 290668 52678 290724 52688
rect 290668 4228 290724 52622
rect 290668 4162 290724 4172
rect 294028 4228 294084 67562
rect 294028 4162 294084 4172
rect 295708 4228 295764 70622
rect 302428 69058 302484 69068
rect 295708 4162 295764 4172
rect 300748 32158 300804 32168
rect 300748 4228 300804 32102
rect 302428 20188 302484 69002
rect 305788 67798 305844 67808
rect 302428 20132 302708 20188
rect 300748 4162 300804 4172
rect 302652 4228 302708 20132
rect 302652 4162 302708 4172
rect 305788 4228 305844 67742
rect 312618 58350 313238 75922
rect 312618 58294 312714 58350
rect 312770 58294 312838 58350
rect 312894 58294 312962 58350
rect 313018 58294 313086 58350
rect 313142 58294 313238 58350
rect 312618 58226 313238 58294
rect 312618 58170 312714 58226
rect 312770 58170 312838 58226
rect 312894 58170 312962 58226
rect 313018 58170 313086 58226
rect 313142 58170 313238 58226
rect 312618 58102 313238 58170
rect 312618 58046 312714 58102
rect 312770 58046 312838 58102
rect 312894 58046 312962 58102
rect 313018 58046 313086 58102
rect 313142 58046 313238 58102
rect 312618 57978 313238 58046
rect 312618 57922 312714 57978
rect 312770 57922 312838 57978
rect 312894 57922 312962 57978
rect 313018 57922 313086 57978
rect 313142 57922 313238 57978
rect 312618 40350 313238 57922
rect 312618 40294 312714 40350
rect 312770 40294 312838 40350
rect 312894 40294 312962 40350
rect 313018 40294 313086 40350
rect 313142 40294 313238 40350
rect 312618 40226 313238 40294
rect 312618 40170 312714 40226
rect 312770 40170 312838 40226
rect 312894 40170 312962 40226
rect 313018 40170 313086 40226
rect 313142 40170 313238 40226
rect 312618 40102 313238 40170
rect 312618 40046 312714 40102
rect 312770 40046 312838 40102
rect 312894 40046 312962 40102
rect 313018 40046 313086 40102
rect 313142 40046 313238 40102
rect 312618 39978 313238 40046
rect 312618 39922 312714 39978
rect 312770 39922 312838 39978
rect 312894 39922 312962 39978
rect 313018 39922 313086 39978
rect 313142 39922 313238 39978
rect 310828 35758 310884 35768
rect 305788 4162 305844 4172
rect 308364 5518 308420 5528
rect 308364 3444 308420 5462
rect 310828 4228 310884 35702
rect 310828 4162 310884 4172
rect 312618 22350 313238 39922
rect 316338 598172 316958 598268
rect 316338 598116 316434 598172
rect 316490 598116 316558 598172
rect 316614 598116 316682 598172
rect 316738 598116 316806 598172
rect 316862 598116 316958 598172
rect 316338 598048 316958 598116
rect 316338 597992 316434 598048
rect 316490 597992 316558 598048
rect 316614 597992 316682 598048
rect 316738 597992 316806 598048
rect 316862 597992 316958 598048
rect 316338 597924 316958 597992
rect 316338 597868 316434 597924
rect 316490 597868 316558 597924
rect 316614 597868 316682 597924
rect 316738 597868 316806 597924
rect 316862 597868 316958 597924
rect 316338 597800 316958 597868
rect 316338 597744 316434 597800
rect 316490 597744 316558 597800
rect 316614 597744 316682 597800
rect 316738 597744 316806 597800
rect 316862 597744 316958 597800
rect 316338 586350 316958 597744
rect 343338 597212 343958 598268
rect 343338 597156 343434 597212
rect 343490 597156 343558 597212
rect 343614 597156 343682 597212
rect 343738 597156 343806 597212
rect 343862 597156 343958 597212
rect 343338 597088 343958 597156
rect 343338 597032 343434 597088
rect 343490 597032 343558 597088
rect 343614 597032 343682 597088
rect 343738 597032 343806 597088
rect 343862 597032 343958 597088
rect 343338 596964 343958 597032
rect 343338 596908 343434 596964
rect 343490 596908 343558 596964
rect 343614 596908 343682 596964
rect 343738 596908 343806 596964
rect 343862 596908 343958 596964
rect 343338 596840 343958 596908
rect 343338 596784 343434 596840
rect 343490 596784 343558 596840
rect 343614 596784 343682 596840
rect 343738 596784 343806 596840
rect 343862 596784 343958 596840
rect 316338 586294 316434 586350
rect 316490 586294 316558 586350
rect 316614 586294 316682 586350
rect 316738 586294 316806 586350
rect 316862 586294 316958 586350
rect 316338 586226 316958 586294
rect 316338 586170 316434 586226
rect 316490 586170 316558 586226
rect 316614 586170 316682 586226
rect 316738 586170 316806 586226
rect 316862 586170 316958 586226
rect 316338 586102 316958 586170
rect 316338 586046 316434 586102
rect 316490 586046 316558 586102
rect 316614 586046 316682 586102
rect 316738 586046 316806 586102
rect 316862 586046 316958 586102
rect 316338 585978 316958 586046
rect 316338 585922 316434 585978
rect 316490 585922 316558 585978
rect 316614 585922 316682 585978
rect 316738 585922 316806 585978
rect 316862 585922 316958 585978
rect 316338 568350 316958 585922
rect 316338 568294 316434 568350
rect 316490 568294 316558 568350
rect 316614 568294 316682 568350
rect 316738 568294 316806 568350
rect 316862 568294 316958 568350
rect 316338 568226 316958 568294
rect 316338 568170 316434 568226
rect 316490 568170 316558 568226
rect 316614 568170 316682 568226
rect 316738 568170 316806 568226
rect 316862 568170 316958 568226
rect 316338 568102 316958 568170
rect 316338 568046 316434 568102
rect 316490 568046 316558 568102
rect 316614 568046 316682 568102
rect 316738 568046 316806 568102
rect 316862 568046 316958 568102
rect 316338 567978 316958 568046
rect 316338 567922 316434 567978
rect 316490 567922 316558 567978
rect 316614 567922 316682 567978
rect 316738 567922 316806 567978
rect 316862 567922 316958 567978
rect 316338 550350 316958 567922
rect 316338 550294 316434 550350
rect 316490 550294 316558 550350
rect 316614 550294 316682 550350
rect 316738 550294 316806 550350
rect 316862 550294 316958 550350
rect 316338 550226 316958 550294
rect 316338 550170 316434 550226
rect 316490 550170 316558 550226
rect 316614 550170 316682 550226
rect 316738 550170 316806 550226
rect 316862 550170 316958 550226
rect 316338 550102 316958 550170
rect 316338 550046 316434 550102
rect 316490 550046 316558 550102
rect 316614 550046 316682 550102
rect 316738 550046 316806 550102
rect 316862 550046 316958 550102
rect 316338 549978 316958 550046
rect 316338 549922 316434 549978
rect 316490 549922 316558 549978
rect 316614 549922 316682 549978
rect 316738 549922 316806 549978
rect 316862 549922 316958 549978
rect 316338 532350 316958 549922
rect 316338 532294 316434 532350
rect 316490 532294 316558 532350
rect 316614 532294 316682 532350
rect 316738 532294 316806 532350
rect 316862 532294 316958 532350
rect 316338 532226 316958 532294
rect 316338 532170 316434 532226
rect 316490 532170 316558 532226
rect 316614 532170 316682 532226
rect 316738 532170 316806 532226
rect 316862 532170 316958 532226
rect 316338 532102 316958 532170
rect 316338 532046 316434 532102
rect 316490 532046 316558 532102
rect 316614 532046 316682 532102
rect 316738 532046 316806 532102
rect 316862 532046 316958 532102
rect 316338 531978 316958 532046
rect 316338 531922 316434 531978
rect 316490 531922 316558 531978
rect 316614 531922 316682 531978
rect 316738 531922 316806 531978
rect 316862 531922 316958 531978
rect 316338 514350 316958 531922
rect 316338 514294 316434 514350
rect 316490 514294 316558 514350
rect 316614 514294 316682 514350
rect 316738 514294 316806 514350
rect 316862 514294 316958 514350
rect 316338 514226 316958 514294
rect 316338 514170 316434 514226
rect 316490 514170 316558 514226
rect 316614 514170 316682 514226
rect 316738 514170 316806 514226
rect 316862 514170 316958 514226
rect 316338 514102 316958 514170
rect 316338 514046 316434 514102
rect 316490 514046 316558 514102
rect 316614 514046 316682 514102
rect 316738 514046 316806 514102
rect 316862 514046 316958 514102
rect 316338 513978 316958 514046
rect 316338 513922 316434 513978
rect 316490 513922 316558 513978
rect 316614 513922 316682 513978
rect 316738 513922 316806 513978
rect 316862 513922 316958 513978
rect 316338 496350 316958 513922
rect 316338 496294 316434 496350
rect 316490 496294 316558 496350
rect 316614 496294 316682 496350
rect 316738 496294 316806 496350
rect 316862 496294 316958 496350
rect 316338 496226 316958 496294
rect 316338 496170 316434 496226
rect 316490 496170 316558 496226
rect 316614 496170 316682 496226
rect 316738 496170 316806 496226
rect 316862 496170 316958 496226
rect 316338 496102 316958 496170
rect 316338 496046 316434 496102
rect 316490 496046 316558 496102
rect 316614 496046 316682 496102
rect 316738 496046 316806 496102
rect 316862 496046 316958 496102
rect 316338 495978 316958 496046
rect 316338 495922 316434 495978
rect 316490 495922 316558 495978
rect 316614 495922 316682 495978
rect 316738 495922 316806 495978
rect 316862 495922 316958 495978
rect 316338 478350 316958 495922
rect 316338 478294 316434 478350
rect 316490 478294 316558 478350
rect 316614 478294 316682 478350
rect 316738 478294 316806 478350
rect 316862 478294 316958 478350
rect 316338 478226 316958 478294
rect 316338 478170 316434 478226
rect 316490 478170 316558 478226
rect 316614 478170 316682 478226
rect 316738 478170 316806 478226
rect 316862 478170 316958 478226
rect 316338 478102 316958 478170
rect 316338 478046 316434 478102
rect 316490 478046 316558 478102
rect 316614 478046 316682 478102
rect 316738 478046 316806 478102
rect 316862 478046 316958 478102
rect 316338 477978 316958 478046
rect 316338 477922 316434 477978
rect 316490 477922 316558 477978
rect 316614 477922 316682 477978
rect 316738 477922 316806 477978
rect 316862 477922 316958 477978
rect 316338 460350 316958 477922
rect 316338 460294 316434 460350
rect 316490 460294 316558 460350
rect 316614 460294 316682 460350
rect 316738 460294 316806 460350
rect 316862 460294 316958 460350
rect 316338 460226 316958 460294
rect 316338 460170 316434 460226
rect 316490 460170 316558 460226
rect 316614 460170 316682 460226
rect 316738 460170 316806 460226
rect 316862 460170 316958 460226
rect 316338 460102 316958 460170
rect 316338 460046 316434 460102
rect 316490 460046 316558 460102
rect 316614 460046 316682 460102
rect 316738 460046 316806 460102
rect 316862 460046 316958 460102
rect 316338 459978 316958 460046
rect 316338 459922 316434 459978
rect 316490 459922 316558 459978
rect 316614 459922 316682 459978
rect 316738 459922 316806 459978
rect 316862 459922 316958 459978
rect 316338 442350 316958 459922
rect 316338 442294 316434 442350
rect 316490 442294 316558 442350
rect 316614 442294 316682 442350
rect 316738 442294 316806 442350
rect 316862 442294 316958 442350
rect 316338 442226 316958 442294
rect 316338 442170 316434 442226
rect 316490 442170 316558 442226
rect 316614 442170 316682 442226
rect 316738 442170 316806 442226
rect 316862 442170 316958 442226
rect 316338 442102 316958 442170
rect 316338 442046 316434 442102
rect 316490 442046 316558 442102
rect 316614 442046 316682 442102
rect 316738 442046 316806 442102
rect 316862 442046 316958 442102
rect 316338 441978 316958 442046
rect 316338 441922 316434 441978
rect 316490 441922 316558 441978
rect 316614 441922 316682 441978
rect 316738 441922 316806 441978
rect 316862 441922 316958 441978
rect 316338 424350 316958 441922
rect 316338 424294 316434 424350
rect 316490 424294 316558 424350
rect 316614 424294 316682 424350
rect 316738 424294 316806 424350
rect 316862 424294 316958 424350
rect 316338 424226 316958 424294
rect 316338 424170 316434 424226
rect 316490 424170 316558 424226
rect 316614 424170 316682 424226
rect 316738 424170 316806 424226
rect 316862 424170 316958 424226
rect 316338 424102 316958 424170
rect 316338 424046 316434 424102
rect 316490 424046 316558 424102
rect 316614 424046 316682 424102
rect 316738 424046 316806 424102
rect 316862 424046 316958 424102
rect 316338 423978 316958 424046
rect 316338 423922 316434 423978
rect 316490 423922 316558 423978
rect 316614 423922 316682 423978
rect 316738 423922 316806 423978
rect 316862 423922 316958 423978
rect 316338 406350 316958 423922
rect 316338 406294 316434 406350
rect 316490 406294 316558 406350
rect 316614 406294 316682 406350
rect 316738 406294 316806 406350
rect 316862 406294 316958 406350
rect 316338 406226 316958 406294
rect 316338 406170 316434 406226
rect 316490 406170 316558 406226
rect 316614 406170 316682 406226
rect 316738 406170 316806 406226
rect 316862 406170 316958 406226
rect 316338 406102 316958 406170
rect 316338 406046 316434 406102
rect 316490 406046 316558 406102
rect 316614 406046 316682 406102
rect 316738 406046 316806 406102
rect 316862 406046 316958 406102
rect 316338 405978 316958 406046
rect 316338 405922 316434 405978
rect 316490 405922 316558 405978
rect 316614 405922 316682 405978
rect 316738 405922 316806 405978
rect 316862 405922 316958 405978
rect 316338 388350 316958 405922
rect 316338 388294 316434 388350
rect 316490 388294 316558 388350
rect 316614 388294 316682 388350
rect 316738 388294 316806 388350
rect 316862 388294 316958 388350
rect 316338 388226 316958 388294
rect 316338 388170 316434 388226
rect 316490 388170 316558 388226
rect 316614 388170 316682 388226
rect 316738 388170 316806 388226
rect 316862 388170 316958 388226
rect 316338 388102 316958 388170
rect 316338 388046 316434 388102
rect 316490 388046 316558 388102
rect 316614 388046 316682 388102
rect 316738 388046 316806 388102
rect 316862 388046 316958 388102
rect 316338 387978 316958 388046
rect 316338 387922 316434 387978
rect 316490 387922 316558 387978
rect 316614 387922 316682 387978
rect 316738 387922 316806 387978
rect 316862 387922 316958 387978
rect 316338 370350 316958 387922
rect 316338 370294 316434 370350
rect 316490 370294 316558 370350
rect 316614 370294 316682 370350
rect 316738 370294 316806 370350
rect 316862 370294 316958 370350
rect 316338 370226 316958 370294
rect 316338 370170 316434 370226
rect 316490 370170 316558 370226
rect 316614 370170 316682 370226
rect 316738 370170 316806 370226
rect 316862 370170 316958 370226
rect 316338 370102 316958 370170
rect 316338 370046 316434 370102
rect 316490 370046 316558 370102
rect 316614 370046 316682 370102
rect 316738 370046 316806 370102
rect 316862 370046 316958 370102
rect 316338 369978 316958 370046
rect 316338 369922 316434 369978
rect 316490 369922 316558 369978
rect 316614 369922 316682 369978
rect 316738 369922 316806 369978
rect 316862 369922 316958 369978
rect 316338 352350 316958 369922
rect 316338 352294 316434 352350
rect 316490 352294 316558 352350
rect 316614 352294 316682 352350
rect 316738 352294 316806 352350
rect 316862 352294 316958 352350
rect 316338 352226 316958 352294
rect 316338 352170 316434 352226
rect 316490 352170 316558 352226
rect 316614 352170 316682 352226
rect 316738 352170 316806 352226
rect 316862 352170 316958 352226
rect 316338 352102 316958 352170
rect 316338 352046 316434 352102
rect 316490 352046 316558 352102
rect 316614 352046 316682 352102
rect 316738 352046 316806 352102
rect 316862 352046 316958 352102
rect 316338 351978 316958 352046
rect 316338 351922 316434 351978
rect 316490 351922 316558 351978
rect 316614 351922 316682 351978
rect 316738 351922 316806 351978
rect 316862 351922 316958 351978
rect 316338 334350 316958 351922
rect 316338 334294 316434 334350
rect 316490 334294 316558 334350
rect 316614 334294 316682 334350
rect 316738 334294 316806 334350
rect 316862 334294 316958 334350
rect 316338 334226 316958 334294
rect 316338 334170 316434 334226
rect 316490 334170 316558 334226
rect 316614 334170 316682 334226
rect 316738 334170 316806 334226
rect 316862 334170 316958 334226
rect 316338 334102 316958 334170
rect 316338 334046 316434 334102
rect 316490 334046 316558 334102
rect 316614 334046 316682 334102
rect 316738 334046 316806 334102
rect 316862 334046 316958 334102
rect 316338 333978 316958 334046
rect 316338 333922 316434 333978
rect 316490 333922 316558 333978
rect 316614 333922 316682 333978
rect 316738 333922 316806 333978
rect 316862 333922 316958 333978
rect 316338 316350 316958 333922
rect 316338 316294 316434 316350
rect 316490 316294 316558 316350
rect 316614 316294 316682 316350
rect 316738 316294 316806 316350
rect 316862 316294 316958 316350
rect 316338 316226 316958 316294
rect 316338 316170 316434 316226
rect 316490 316170 316558 316226
rect 316614 316170 316682 316226
rect 316738 316170 316806 316226
rect 316862 316170 316958 316226
rect 316338 316102 316958 316170
rect 316338 316046 316434 316102
rect 316490 316046 316558 316102
rect 316614 316046 316682 316102
rect 316738 316046 316806 316102
rect 316862 316046 316958 316102
rect 316338 315978 316958 316046
rect 316338 315922 316434 315978
rect 316490 315922 316558 315978
rect 316614 315922 316682 315978
rect 316738 315922 316806 315978
rect 316862 315922 316958 315978
rect 316338 298350 316958 315922
rect 316338 298294 316434 298350
rect 316490 298294 316558 298350
rect 316614 298294 316682 298350
rect 316738 298294 316806 298350
rect 316862 298294 316958 298350
rect 316338 298226 316958 298294
rect 316338 298170 316434 298226
rect 316490 298170 316558 298226
rect 316614 298170 316682 298226
rect 316738 298170 316806 298226
rect 316862 298170 316958 298226
rect 316338 298102 316958 298170
rect 316338 298046 316434 298102
rect 316490 298046 316558 298102
rect 316614 298046 316682 298102
rect 316738 298046 316806 298102
rect 316862 298046 316958 298102
rect 316338 297978 316958 298046
rect 316338 297922 316434 297978
rect 316490 297922 316558 297978
rect 316614 297922 316682 297978
rect 316738 297922 316806 297978
rect 316862 297922 316958 297978
rect 316338 280350 316958 297922
rect 316338 280294 316434 280350
rect 316490 280294 316558 280350
rect 316614 280294 316682 280350
rect 316738 280294 316806 280350
rect 316862 280294 316958 280350
rect 316338 280226 316958 280294
rect 316338 280170 316434 280226
rect 316490 280170 316558 280226
rect 316614 280170 316682 280226
rect 316738 280170 316806 280226
rect 316862 280170 316958 280226
rect 316338 280102 316958 280170
rect 316338 280046 316434 280102
rect 316490 280046 316558 280102
rect 316614 280046 316682 280102
rect 316738 280046 316806 280102
rect 316862 280046 316958 280102
rect 316338 279978 316958 280046
rect 316338 279922 316434 279978
rect 316490 279922 316558 279978
rect 316614 279922 316682 279978
rect 316738 279922 316806 279978
rect 316862 279922 316958 279978
rect 316338 262350 316958 279922
rect 316338 262294 316434 262350
rect 316490 262294 316558 262350
rect 316614 262294 316682 262350
rect 316738 262294 316806 262350
rect 316862 262294 316958 262350
rect 316338 262226 316958 262294
rect 316338 262170 316434 262226
rect 316490 262170 316558 262226
rect 316614 262170 316682 262226
rect 316738 262170 316806 262226
rect 316862 262170 316958 262226
rect 316338 262102 316958 262170
rect 316338 262046 316434 262102
rect 316490 262046 316558 262102
rect 316614 262046 316682 262102
rect 316738 262046 316806 262102
rect 316862 262046 316958 262102
rect 316338 261978 316958 262046
rect 316338 261922 316434 261978
rect 316490 261922 316558 261978
rect 316614 261922 316682 261978
rect 316738 261922 316806 261978
rect 316862 261922 316958 261978
rect 316338 244350 316958 261922
rect 316338 244294 316434 244350
rect 316490 244294 316558 244350
rect 316614 244294 316682 244350
rect 316738 244294 316806 244350
rect 316862 244294 316958 244350
rect 316338 244226 316958 244294
rect 316338 244170 316434 244226
rect 316490 244170 316558 244226
rect 316614 244170 316682 244226
rect 316738 244170 316806 244226
rect 316862 244170 316958 244226
rect 316338 244102 316958 244170
rect 316338 244046 316434 244102
rect 316490 244046 316558 244102
rect 316614 244046 316682 244102
rect 316738 244046 316806 244102
rect 316862 244046 316958 244102
rect 316338 243978 316958 244046
rect 316338 243922 316434 243978
rect 316490 243922 316558 243978
rect 316614 243922 316682 243978
rect 316738 243922 316806 243978
rect 316862 243922 316958 243978
rect 316338 226350 316958 243922
rect 316338 226294 316434 226350
rect 316490 226294 316558 226350
rect 316614 226294 316682 226350
rect 316738 226294 316806 226350
rect 316862 226294 316958 226350
rect 316338 226226 316958 226294
rect 316338 226170 316434 226226
rect 316490 226170 316558 226226
rect 316614 226170 316682 226226
rect 316738 226170 316806 226226
rect 316862 226170 316958 226226
rect 316338 226102 316958 226170
rect 316338 226046 316434 226102
rect 316490 226046 316558 226102
rect 316614 226046 316682 226102
rect 316738 226046 316806 226102
rect 316862 226046 316958 226102
rect 316338 225978 316958 226046
rect 316338 225922 316434 225978
rect 316490 225922 316558 225978
rect 316614 225922 316682 225978
rect 316738 225922 316806 225978
rect 316862 225922 316958 225978
rect 316338 208350 316958 225922
rect 316338 208294 316434 208350
rect 316490 208294 316558 208350
rect 316614 208294 316682 208350
rect 316738 208294 316806 208350
rect 316862 208294 316958 208350
rect 316338 208226 316958 208294
rect 316338 208170 316434 208226
rect 316490 208170 316558 208226
rect 316614 208170 316682 208226
rect 316738 208170 316806 208226
rect 316862 208170 316958 208226
rect 316338 208102 316958 208170
rect 316338 208046 316434 208102
rect 316490 208046 316558 208102
rect 316614 208046 316682 208102
rect 316738 208046 316806 208102
rect 316862 208046 316958 208102
rect 316338 207978 316958 208046
rect 316338 207922 316434 207978
rect 316490 207922 316558 207978
rect 316614 207922 316682 207978
rect 316738 207922 316806 207978
rect 316862 207922 316958 207978
rect 316338 190350 316958 207922
rect 316338 190294 316434 190350
rect 316490 190294 316558 190350
rect 316614 190294 316682 190350
rect 316738 190294 316806 190350
rect 316862 190294 316958 190350
rect 316338 190226 316958 190294
rect 316338 190170 316434 190226
rect 316490 190170 316558 190226
rect 316614 190170 316682 190226
rect 316738 190170 316806 190226
rect 316862 190170 316958 190226
rect 316338 190102 316958 190170
rect 316338 190046 316434 190102
rect 316490 190046 316558 190102
rect 316614 190046 316682 190102
rect 316738 190046 316806 190102
rect 316862 190046 316958 190102
rect 316338 189978 316958 190046
rect 316338 189922 316434 189978
rect 316490 189922 316558 189978
rect 316614 189922 316682 189978
rect 316738 189922 316806 189978
rect 316862 189922 316958 189978
rect 316338 172350 316958 189922
rect 316338 172294 316434 172350
rect 316490 172294 316558 172350
rect 316614 172294 316682 172350
rect 316738 172294 316806 172350
rect 316862 172294 316958 172350
rect 316338 172226 316958 172294
rect 316338 172170 316434 172226
rect 316490 172170 316558 172226
rect 316614 172170 316682 172226
rect 316738 172170 316806 172226
rect 316862 172170 316958 172226
rect 316338 172102 316958 172170
rect 316338 172046 316434 172102
rect 316490 172046 316558 172102
rect 316614 172046 316682 172102
rect 316738 172046 316806 172102
rect 316862 172046 316958 172102
rect 316338 171978 316958 172046
rect 316338 171922 316434 171978
rect 316490 171922 316558 171978
rect 316614 171922 316682 171978
rect 316738 171922 316806 171978
rect 316862 171922 316958 171978
rect 316338 154350 316958 171922
rect 316338 154294 316434 154350
rect 316490 154294 316558 154350
rect 316614 154294 316682 154350
rect 316738 154294 316806 154350
rect 316862 154294 316958 154350
rect 316338 154226 316958 154294
rect 316338 154170 316434 154226
rect 316490 154170 316558 154226
rect 316614 154170 316682 154226
rect 316738 154170 316806 154226
rect 316862 154170 316958 154226
rect 316338 154102 316958 154170
rect 316338 154046 316434 154102
rect 316490 154046 316558 154102
rect 316614 154046 316682 154102
rect 316738 154046 316806 154102
rect 316862 154046 316958 154102
rect 316338 153978 316958 154046
rect 316338 153922 316434 153978
rect 316490 153922 316558 153978
rect 316614 153922 316682 153978
rect 316738 153922 316806 153978
rect 316862 153922 316958 153978
rect 316338 136350 316958 153922
rect 316338 136294 316434 136350
rect 316490 136294 316558 136350
rect 316614 136294 316682 136350
rect 316738 136294 316806 136350
rect 316862 136294 316958 136350
rect 316338 136226 316958 136294
rect 316338 136170 316434 136226
rect 316490 136170 316558 136226
rect 316614 136170 316682 136226
rect 316738 136170 316806 136226
rect 316862 136170 316958 136226
rect 316338 136102 316958 136170
rect 316338 136046 316434 136102
rect 316490 136046 316558 136102
rect 316614 136046 316682 136102
rect 316738 136046 316806 136102
rect 316862 136046 316958 136102
rect 316338 135978 316958 136046
rect 316338 135922 316434 135978
rect 316490 135922 316558 135978
rect 316614 135922 316682 135978
rect 316738 135922 316806 135978
rect 316862 135922 316958 135978
rect 316338 118350 316958 135922
rect 316338 118294 316434 118350
rect 316490 118294 316558 118350
rect 316614 118294 316682 118350
rect 316738 118294 316806 118350
rect 316862 118294 316958 118350
rect 316338 118226 316958 118294
rect 316338 118170 316434 118226
rect 316490 118170 316558 118226
rect 316614 118170 316682 118226
rect 316738 118170 316806 118226
rect 316862 118170 316958 118226
rect 316338 118102 316958 118170
rect 316338 118046 316434 118102
rect 316490 118046 316558 118102
rect 316614 118046 316682 118102
rect 316738 118046 316806 118102
rect 316862 118046 316958 118102
rect 316338 117978 316958 118046
rect 316338 117922 316434 117978
rect 316490 117922 316558 117978
rect 316614 117922 316682 117978
rect 316738 117922 316806 117978
rect 316862 117922 316958 117978
rect 316338 100350 316958 117922
rect 316338 100294 316434 100350
rect 316490 100294 316558 100350
rect 316614 100294 316682 100350
rect 316738 100294 316806 100350
rect 316862 100294 316958 100350
rect 316338 100226 316958 100294
rect 316338 100170 316434 100226
rect 316490 100170 316558 100226
rect 316614 100170 316682 100226
rect 316738 100170 316806 100226
rect 316862 100170 316958 100226
rect 316338 100102 316958 100170
rect 316338 100046 316434 100102
rect 316490 100046 316558 100102
rect 316614 100046 316682 100102
rect 316738 100046 316806 100102
rect 316862 100046 316958 100102
rect 316338 99978 316958 100046
rect 316338 99922 316434 99978
rect 316490 99922 316558 99978
rect 316614 99922 316682 99978
rect 316738 99922 316806 99978
rect 316862 99922 316958 99978
rect 316338 82350 316958 99922
rect 316338 82294 316434 82350
rect 316490 82294 316558 82350
rect 316614 82294 316682 82350
rect 316738 82294 316806 82350
rect 316862 82294 316958 82350
rect 316338 82226 316958 82294
rect 316338 82170 316434 82226
rect 316490 82170 316558 82226
rect 316614 82170 316682 82226
rect 316738 82170 316806 82226
rect 316862 82170 316958 82226
rect 316338 82102 316958 82170
rect 316338 82046 316434 82102
rect 316490 82046 316558 82102
rect 316614 82046 316682 82102
rect 316738 82046 316806 82102
rect 316862 82046 316958 82102
rect 316338 81978 316958 82046
rect 316338 81922 316434 81978
rect 316490 81922 316558 81978
rect 316614 81922 316682 81978
rect 316738 81922 316806 81978
rect 316862 81922 316958 81978
rect 316338 64350 316958 81922
rect 341068 590212 341124 590222
rect 341068 79858 341124 590156
rect 341068 79792 341124 79802
rect 343338 580350 343958 596784
rect 343338 580294 343434 580350
rect 343490 580294 343558 580350
rect 343614 580294 343682 580350
rect 343738 580294 343806 580350
rect 343862 580294 343958 580350
rect 343338 580226 343958 580294
rect 343338 580170 343434 580226
rect 343490 580170 343558 580226
rect 343614 580170 343682 580226
rect 343738 580170 343806 580226
rect 343862 580170 343958 580226
rect 343338 580102 343958 580170
rect 343338 580046 343434 580102
rect 343490 580046 343558 580102
rect 343614 580046 343682 580102
rect 343738 580046 343806 580102
rect 343862 580046 343958 580102
rect 343338 579978 343958 580046
rect 343338 579922 343434 579978
rect 343490 579922 343558 579978
rect 343614 579922 343682 579978
rect 343738 579922 343806 579978
rect 343862 579922 343958 579978
rect 343338 562350 343958 579922
rect 343338 562294 343434 562350
rect 343490 562294 343558 562350
rect 343614 562294 343682 562350
rect 343738 562294 343806 562350
rect 343862 562294 343958 562350
rect 343338 562226 343958 562294
rect 343338 562170 343434 562226
rect 343490 562170 343558 562226
rect 343614 562170 343682 562226
rect 343738 562170 343806 562226
rect 343862 562170 343958 562226
rect 343338 562102 343958 562170
rect 343338 562046 343434 562102
rect 343490 562046 343558 562102
rect 343614 562046 343682 562102
rect 343738 562046 343806 562102
rect 343862 562046 343958 562102
rect 343338 561978 343958 562046
rect 343338 561922 343434 561978
rect 343490 561922 343558 561978
rect 343614 561922 343682 561978
rect 343738 561922 343806 561978
rect 343862 561922 343958 561978
rect 343338 544350 343958 561922
rect 343338 544294 343434 544350
rect 343490 544294 343558 544350
rect 343614 544294 343682 544350
rect 343738 544294 343806 544350
rect 343862 544294 343958 544350
rect 343338 544226 343958 544294
rect 343338 544170 343434 544226
rect 343490 544170 343558 544226
rect 343614 544170 343682 544226
rect 343738 544170 343806 544226
rect 343862 544170 343958 544226
rect 343338 544102 343958 544170
rect 343338 544046 343434 544102
rect 343490 544046 343558 544102
rect 343614 544046 343682 544102
rect 343738 544046 343806 544102
rect 343862 544046 343958 544102
rect 343338 543978 343958 544046
rect 343338 543922 343434 543978
rect 343490 543922 343558 543978
rect 343614 543922 343682 543978
rect 343738 543922 343806 543978
rect 343862 543922 343958 543978
rect 343338 526350 343958 543922
rect 343338 526294 343434 526350
rect 343490 526294 343558 526350
rect 343614 526294 343682 526350
rect 343738 526294 343806 526350
rect 343862 526294 343958 526350
rect 343338 526226 343958 526294
rect 343338 526170 343434 526226
rect 343490 526170 343558 526226
rect 343614 526170 343682 526226
rect 343738 526170 343806 526226
rect 343862 526170 343958 526226
rect 343338 526102 343958 526170
rect 343338 526046 343434 526102
rect 343490 526046 343558 526102
rect 343614 526046 343682 526102
rect 343738 526046 343806 526102
rect 343862 526046 343958 526102
rect 343338 525978 343958 526046
rect 343338 525922 343434 525978
rect 343490 525922 343558 525978
rect 343614 525922 343682 525978
rect 343738 525922 343806 525978
rect 343862 525922 343958 525978
rect 343338 508350 343958 525922
rect 343338 508294 343434 508350
rect 343490 508294 343558 508350
rect 343614 508294 343682 508350
rect 343738 508294 343806 508350
rect 343862 508294 343958 508350
rect 343338 508226 343958 508294
rect 343338 508170 343434 508226
rect 343490 508170 343558 508226
rect 343614 508170 343682 508226
rect 343738 508170 343806 508226
rect 343862 508170 343958 508226
rect 343338 508102 343958 508170
rect 343338 508046 343434 508102
rect 343490 508046 343558 508102
rect 343614 508046 343682 508102
rect 343738 508046 343806 508102
rect 343862 508046 343958 508102
rect 343338 507978 343958 508046
rect 343338 507922 343434 507978
rect 343490 507922 343558 507978
rect 343614 507922 343682 507978
rect 343738 507922 343806 507978
rect 343862 507922 343958 507978
rect 343338 490350 343958 507922
rect 343338 490294 343434 490350
rect 343490 490294 343558 490350
rect 343614 490294 343682 490350
rect 343738 490294 343806 490350
rect 343862 490294 343958 490350
rect 343338 490226 343958 490294
rect 343338 490170 343434 490226
rect 343490 490170 343558 490226
rect 343614 490170 343682 490226
rect 343738 490170 343806 490226
rect 343862 490170 343958 490226
rect 343338 490102 343958 490170
rect 343338 490046 343434 490102
rect 343490 490046 343558 490102
rect 343614 490046 343682 490102
rect 343738 490046 343806 490102
rect 343862 490046 343958 490102
rect 343338 489978 343958 490046
rect 343338 489922 343434 489978
rect 343490 489922 343558 489978
rect 343614 489922 343682 489978
rect 343738 489922 343806 489978
rect 343862 489922 343958 489978
rect 343338 472350 343958 489922
rect 343338 472294 343434 472350
rect 343490 472294 343558 472350
rect 343614 472294 343682 472350
rect 343738 472294 343806 472350
rect 343862 472294 343958 472350
rect 343338 472226 343958 472294
rect 343338 472170 343434 472226
rect 343490 472170 343558 472226
rect 343614 472170 343682 472226
rect 343738 472170 343806 472226
rect 343862 472170 343958 472226
rect 343338 472102 343958 472170
rect 343338 472046 343434 472102
rect 343490 472046 343558 472102
rect 343614 472046 343682 472102
rect 343738 472046 343806 472102
rect 343862 472046 343958 472102
rect 343338 471978 343958 472046
rect 343338 471922 343434 471978
rect 343490 471922 343558 471978
rect 343614 471922 343682 471978
rect 343738 471922 343806 471978
rect 343862 471922 343958 471978
rect 343338 454350 343958 471922
rect 343338 454294 343434 454350
rect 343490 454294 343558 454350
rect 343614 454294 343682 454350
rect 343738 454294 343806 454350
rect 343862 454294 343958 454350
rect 343338 454226 343958 454294
rect 343338 454170 343434 454226
rect 343490 454170 343558 454226
rect 343614 454170 343682 454226
rect 343738 454170 343806 454226
rect 343862 454170 343958 454226
rect 343338 454102 343958 454170
rect 343338 454046 343434 454102
rect 343490 454046 343558 454102
rect 343614 454046 343682 454102
rect 343738 454046 343806 454102
rect 343862 454046 343958 454102
rect 343338 453978 343958 454046
rect 343338 453922 343434 453978
rect 343490 453922 343558 453978
rect 343614 453922 343682 453978
rect 343738 453922 343806 453978
rect 343862 453922 343958 453978
rect 343338 436350 343958 453922
rect 343338 436294 343434 436350
rect 343490 436294 343558 436350
rect 343614 436294 343682 436350
rect 343738 436294 343806 436350
rect 343862 436294 343958 436350
rect 343338 436226 343958 436294
rect 343338 436170 343434 436226
rect 343490 436170 343558 436226
rect 343614 436170 343682 436226
rect 343738 436170 343806 436226
rect 343862 436170 343958 436226
rect 343338 436102 343958 436170
rect 343338 436046 343434 436102
rect 343490 436046 343558 436102
rect 343614 436046 343682 436102
rect 343738 436046 343806 436102
rect 343862 436046 343958 436102
rect 343338 435978 343958 436046
rect 343338 435922 343434 435978
rect 343490 435922 343558 435978
rect 343614 435922 343682 435978
rect 343738 435922 343806 435978
rect 343862 435922 343958 435978
rect 343338 418350 343958 435922
rect 343338 418294 343434 418350
rect 343490 418294 343558 418350
rect 343614 418294 343682 418350
rect 343738 418294 343806 418350
rect 343862 418294 343958 418350
rect 343338 418226 343958 418294
rect 343338 418170 343434 418226
rect 343490 418170 343558 418226
rect 343614 418170 343682 418226
rect 343738 418170 343806 418226
rect 343862 418170 343958 418226
rect 343338 418102 343958 418170
rect 343338 418046 343434 418102
rect 343490 418046 343558 418102
rect 343614 418046 343682 418102
rect 343738 418046 343806 418102
rect 343862 418046 343958 418102
rect 343338 417978 343958 418046
rect 343338 417922 343434 417978
rect 343490 417922 343558 417978
rect 343614 417922 343682 417978
rect 343738 417922 343806 417978
rect 343862 417922 343958 417978
rect 343338 400350 343958 417922
rect 343338 400294 343434 400350
rect 343490 400294 343558 400350
rect 343614 400294 343682 400350
rect 343738 400294 343806 400350
rect 343862 400294 343958 400350
rect 343338 400226 343958 400294
rect 343338 400170 343434 400226
rect 343490 400170 343558 400226
rect 343614 400170 343682 400226
rect 343738 400170 343806 400226
rect 343862 400170 343958 400226
rect 343338 400102 343958 400170
rect 343338 400046 343434 400102
rect 343490 400046 343558 400102
rect 343614 400046 343682 400102
rect 343738 400046 343806 400102
rect 343862 400046 343958 400102
rect 343338 399978 343958 400046
rect 343338 399922 343434 399978
rect 343490 399922 343558 399978
rect 343614 399922 343682 399978
rect 343738 399922 343806 399978
rect 343862 399922 343958 399978
rect 343338 382350 343958 399922
rect 343338 382294 343434 382350
rect 343490 382294 343558 382350
rect 343614 382294 343682 382350
rect 343738 382294 343806 382350
rect 343862 382294 343958 382350
rect 343338 382226 343958 382294
rect 343338 382170 343434 382226
rect 343490 382170 343558 382226
rect 343614 382170 343682 382226
rect 343738 382170 343806 382226
rect 343862 382170 343958 382226
rect 343338 382102 343958 382170
rect 343338 382046 343434 382102
rect 343490 382046 343558 382102
rect 343614 382046 343682 382102
rect 343738 382046 343806 382102
rect 343862 382046 343958 382102
rect 343338 381978 343958 382046
rect 343338 381922 343434 381978
rect 343490 381922 343558 381978
rect 343614 381922 343682 381978
rect 343738 381922 343806 381978
rect 343862 381922 343958 381978
rect 343338 364350 343958 381922
rect 343338 364294 343434 364350
rect 343490 364294 343558 364350
rect 343614 364294 343682 364350
rect 343738 364294 343806 364350
rect 343862 364294 343958 364350
rect 343338 364226 343958 364294
rect 343338 364170 343434 364226
rect 343490 364170 343558 364226
rect 343614 364170 343682 364226
rect 343738 364170 343806 364226
rect 343862 364170 343958 364226
rect 343338 364102 343958 364170
rect 343338 364046 343434 364102
rect 343490 364046 343558 364102
rect 343614 364046 343682 364102
rect 343738 364046 343806 364102
rect 343862 364046 343958 364102
rect 343338 363978 343958 364046
rect 343338 363922 343434 363978
rect 343490 363922 343558 363978
rect 343614 363922 343682 363978
rect 343738 363922 343806 363978
rect 343862 363922 343958 363978
rect 343338 346350 343958 363922
rect 343338 346294 343434 346350
rect 343490 346294 343558 346350
rect 343614 346294 343682 346350
rect 343738 346294 343806 346350
rect 343862 346294 343958 346350
rect 343338 346226 343958 346294
rect 343338 346170 343434 346226
rect 343490 346170 343558 346226
rect 343614 346170 343682 346226
rect 343738 346170 343806 346226
rect 343862 346170 343958 346226
rect 343338 346102 343958 346170
rect 343338 346046 343434 346102
rect 343490 346046 343558 346102
rect 343614 346046 343682 346102
rect 343738 346046 343806 346102
rect 343862 346046 343958 346102
rect 343338 345978 343958 346046
rect 343338 345922 343434 345978
rect 343490 345922 343558 345978
rect 343614 345922 343682 345978
rect 343738 345922 343806 345978
rect 343862 345922 343958 345978
rect 343338 328350 343958 345922
rect 343338 328294 343434 328350
rect 343490 328294 343558 328350
rect 343614 328294 343682 328350
rect 343738 328294 343806 328350
rect 343862 328294 343958 328350
rect 343338 328226 343958 328294
rect 343338 328170 343434 328226
rect 343490 328170 343558 328226
rect 343614 328170 343682 328226
rect 343738 328170 343806 328226
rect 343862 328170 343958 328226
rect 343338 328102 343958 328170
rect 343338 328046 343434 328102
rect 343490 328046 343558 328102
rect 343614 328046 343682 328102
rect 343738 328046 343806 328102
rect 343862 328046 343958 328102
rect 343338 327978 343958 328046
rect 343338 327922 343434 327978
rect 343490 327922 343558 327978
rect 343614 327922 343682 327978
rect 343738 327922 343806 327978
rect 343862 327922 343958 327978
rect 343338 310350 343958 327922
rect 343338 310294 343434 310350
rect 343490 310294 343558 310350
rect 343614 310294 343682 310350
rect 343738 310294 343806 310350
rect 343862 310294 343958 310350
rect 343338 310226 343958 310294
rect 343338 310170 343434 310226
rect 343490 310170 343558 310226
rect 343614 310170 343682 310226
rect 343738 310170 343806 310226
rect 343862 310170 343958 310226
rect 343338 310102 343958 310170
rect 343338 310046 343434 310102
rect 343490 310046 343558 310102
rect 343614 310046 343682 310102
rect 343738 310046 343806 310102
rect 343862 310046 343958 310102
rect 343338 309978 343958 310046
rect 343338 309922 343434 309978
rect 343490 309922 343558 309978
rect 343614 309922 343682 309978
rect 343738 309922 343806 309978
rect 343862 309922 343958 309978
rect 343338 292350 343958 309922
rect 343338 292294 343434 292350
rect 343490 292294 343558 292350
rect 343614 292294 343682 292350
rect 343738 292294 343806 292350
rect 343862 292294 343958 292350
rect 343338 292226 343958 292294
rect 343338 292170 343434 292226
rect 343490 292170 343558 292226
rect 343614 292170 343682 292226
rect 343738 292170 343806 292226
rect 343862 292170 343958 292226
rect 343338 292102 343958 292170
rect 343338 292046 343434 292102
rect 343490 292046 343558 292102
rect 343614 292046 343682 292102
rect 343738 292046 343806 292102
rect 343862 292046 343958 292102
rect 343338 291978 343958 292046
rect 343338 291922 343434 291978
rect 343490 291922 343558 291978
rect 343614 291922 343682 291978
rect 343738 291922 343806 291978
rect 343862 291922 343958 291978
rect 343338 274350 343958 291922
rect 343338 274294 343434 274350
rect 343490 274294 343558 274350
rect 343614 274294 343682 274350
rect 343738 274294 343806 274350
rect 343862 274294 343958 274350
rect 343338 274226 343958 274294
rect 343338 274170 343434 274226
rect 343490 274170 343558 274226
rect 343614 274170 343682 274226
rect 343738 274170 343806 274226
rect 343862 274170 343958 274226
rect 343338 274102 343958 274170
rect 343338 274046 343434 274102
rect 343490 274046 343558 274102
rect 343614 274046 343682 274102
rect 343738 274046 343806 274102
rect 343862 274046 343958 274102
rect 343338 273978 343958 274046
rect 343338 273922 343434 273978
rect 343490 273922 343558 273978
rect 343614 273922 343682 273978
rect 343738 273922 343806 273978
rect 343862 273922 343958 273978
rect 343338 256350 343958 273922
rect 343338 256294 343434 256350
rect 343490 256294 343558 256350
rect 343614 256294 343682 256350
rect 343738 256294 343806 256350
rect 343862 256294 343958 256350
rect 343338 256226 343958 256294
rect 343338 256170 343434 256226
rect 343490 256170 343558 256226
rect 343614 256170 343682 256226
rect 343738 256170 343806 256226
rect 343862 256170 343958 256226
rect 343338 256102 343958 256170
rect 343338 256046 343434 256102
rect 343490 256046 343558 256102
rect 343614 256046 343682 256102
rect 343738 256046 343806 256102
rect 343862 256046 343958 256102
rect 343338 255978 343958 256046
rect 343338 255922 343434 255978
rect 343490 255922 343558 255978
rect 343614 255922 343682 255978
rect 343738 255922 343806 255978
rect 343862 255922 343958 255978
rect 343338 238350 343958 255922
rect 343338 238294 343434 238350
rect 343490 238294 343558 238350
rect 343614 238294 343682 238350
rect 343738 238294 343806 238350
rect 343862 238294 343958 238350
rect 343338 238226 343958 238294
rect 343338 238170 343434 238226
rect 343490 238170 343558 238226
rect 343614 238170 343682 238226
rect 343738 238170 343806 238226
rect 343862 238170 343958 238226
rect 343338 238102 343958 238170
rect 343338 238046 343434 238102
rect 343490 238046 343558 238102
rect 343614 238046 343682 238102
rect 343738 238046 343806 238102
rect 343862 238046 343958 238102
rect 343338 237978 343958 238046
rect 343338 237922 343434 237978
rect 343490 237922 343558 237978
rect 343614 237922 343682 237978
rect 343738 237922 343806 237978
rect 343862 237922 343958 237978
rect 343338 220350 343958 237922
rect 343338 220294 343434 220350
rect 343490 220294 343558 220350
rect 343614 220294 343682 220350
rect 343738 220294 343806 220350
rect 343862 220294 343958 220350
rect 343338 220226 343958 220294
rect 343338 220170 343434 220226
rect 343490 220170 343558 220226
rect 343614 220170 343682 220226
rect 343738 220170 343806 220226
rect 343862 220170 343958 220226
rect 343338 220102 343958 220170
rect 343338 220046 343434 220102
rect 343490 220046 343558 220102
rect 343614 220046 343682 220102
rect 343738 220046 343806 220102
rect 343862 220046 343958 220102
rect 343338 219978 343958 220046
rect 343338 219922 343434 219978
rect 343490 219922 343558 219978
rect 343614 219922 343682 219978
rect 343738 219922 343806 219978
rect 343862 219922 343958 219978
rect 343338 202350 343958 219922
rect 343338 202294 343434 202350
rect 343490 202294 343558 202350
rect 343614 202294 343682 202350
rect 343738 202294 343806 202350
rect 343862 202294 343958 202350
rect 343338 202226 343958 202294
rect 343338 202170 343434 202226
rect 343490 202170 343558 202226
rect 343614 202170 343682 202226
rect 343738 202170 343806 202226
rect 343862 202170 343958 202226
rect 343338 202102 343958 202170
rect 343338 202046 343434 202102
rect 343490 202046 343558 202102
rect 343614 202046 343682 202102
rect 343738 202046 343806 202102
rect 343862 202046 343958 202102
rect 343338 201978 343958 202046
rect 343338 201922 343434 201978
rect 343490 201922 343558 201978
rect 343614 201922 343682 201978
rect 343738 201922 343806 201978
rect 343862 201922 343958 201978
rect 343338 184350 343958 201922
rect 343338 184294 343434 184350
rect 343490 184294 343558 184350
rect 343614 184294 343682 184350
rect 343738 184294 343806 184350
rect 343862 184294 343958 184350
rect 343338 184226 343958 184294
rect 343338 184170 343434 184226
rect 343490 184170 343558 184226
rect 343614 184170 343682 184226
rect 343738 184170 343806 184226
rect 343862 184170 343958 184226
rect 343338 184102 343958 184170
rect 343338 184046 343434 184102
rect 343490 184046 343558 184102
rect 343614 184046 343682 184102
rect 343738 184046 343806 184102
rect 343862 184046 343958 184102
rect 343338 183978 343958 184046
rect 343338 183922 343434 183978
rect 343490 183922 343558 183978
rect 343614 183922 343682 183978
rect 343738 183922 343806 183978
rect 343862 183922 343958 183978
rect 343338 166350 343958 183922
rect 343338 166294 343434 166350
rect 343490 166294 343558 166350
rect 343614 166294 343682 166350
rect 343738 166294 343806 166350
rect 343862 166294 343958 166350
rect 343338 166226 343958 166294
rect 343338 166170 343434 166226
rect 343490 166170 343558 166226
rect 343614 166170 343682 166226
rect 343738 166170 343806 166226
rect 343862 166170 343958 166226
rect 343338 166102 343958 166170
rect 343338 166046 343434 166102
rect 343490 166046 343558 166102
rect 343614 166046 343682 166102
rect 343738 166046 343806 166102
rect 343862 166046 343958 166102
rect 343338 165978 343958 166046
rect 343338 165922 343434 165978
rect 343490 165922 343558 165978
rect 343614 165922 343682 165978
rect 343738 165922 343806 165978
rect 343862 165922 343958 165978
rect 343338 148350 343958 165922
rect 343338 148294 343434 148350
rect 343490 148294 343558 148350
rect 343614 148294 343682 148350
rect 343738 148294 343806 148350
rect 343862 148294 343958 148350
rect 343338 148226 343958 148294
rect 343338 148170 343434 148226
rect 343490 148170 343558 148226
rect 343614 148170 343682 148226
rect 343738 148170 343806 148226
rect 343862 148170 343958 148226
rect 343338 148102 343958 148170
rect 343338 148046 343434 148102
rect 343490 148046 343558 148102
rect 343614 148046 343682 148102
rect 343738 148046 343806 148102
rect 343862 148046 343958 148102
rect 343338 147978 343958 148046
rect 343338 147922 343434 147978
rect 343490 147922 343558 147978
rect 343614 147922 343682 147978
rect 343738 147922 343806 147978
rect 343862 147922 343958 147978
rect 343338 130350 343958 147922
rect 343338 130294 343434 130350
rect 343490 130294 343558 130350
rect 343614 130294 343682 130350
rect 343738 130294 343806 130350
rect 343862 130294 343958 130350
rect 343338 130226 343958 130294
rect 343338 130170 343434 130226
rect 343490 130170 343558 130226
rect 343614 130170 343682 130226
rect 343738 130170 343806 130226
rect 343862 130170 343958 130226
rect 343338 130102 343958 130170
rect 343338 130046 343434 130102
rect 343490 130046 343558 130102
rect 343614 130046 343682 130102
rect 343738 130046 343806 130102
rect 343862 130046 343958 130102
rect 343338 129978 343958 130046
rect 343338 129922 343434 129978
rect 343490 129922 343558 129978
rect 343614 129922 343682 129978
rect 343738 129922 343806 129978
rect 343862 129922 343958 129978
rect 343338 112350 343958 129922
rect 343338 112294 343434 112350
rect 343490 112294 343558 112350
rect 343614 112294 343682 112350
rect 343738 112294 343806 112350
rect 343862 112294 343958 112350
rect 343338 112226 343958 112294
rect 343338 112170 343434 112226
rect 343490 112170 343558 112226
rect 343614 112170 343682 112226
rect 343738 112170 343806 112226
rect 343862 112170 343958 112226
rect 343338 112102 343958 112170
rect 343338 112046 343434 112102
rect 343490 112046 343558 112102
rect 343614 112046 343682 112102
rect 343738 112046 343806 112102
rect 343862 112046 343958 112102
rect 343338 111978 343958 112046
rect 343338 111922 343434 111978
rect 343490 111922 343558 111978
rect 343614 111922 343682 111978
rect 343738 111922 343806 111978
rect 343862 111922 343958 111978
rect 343338 94350 343958 111922
rect 343338 94294 343434 94350
rect 343490 94294 343558 94350
rect 343614 94294 343682 94350
rect 343738 94294 343806 94350
rect 343862 94294 343958 94350
rect 343338 94226 343958 94294
rect 343338 94170 343434 94226
rect 343490 94170 343558 94226
rect 343614 94170 343682 94226
rect 343738 94170 343806 94226
rect 343862 94170 343958 94226
rect 343338 94102 343958 94170
rect 343338 94046 343434 94102
rect 343490 94046 343558 94102
rect 343614 94046 343682 94102
rect 343738 94046 343806 94102
rect 343862 94046 343958 94102
rect 343338 93978 343958 94046
rect 343338 93922 343434 93978
rect 343490 93922 343558 93978
rect 343614 93922 343682 93978
rect 343738 93922 343806 93978
rect 343862 93922 343958 93978
rect 343338 76350 343958 93922
rect 343338 76294 343434 76350
rect 343490 76294 343558 76350
rect 343614 76294 343682 76350
rect 343738 76294 343806 76350
rect 343862 76294 343958 76350
rect 343338 76226 343958 76294
rect 343338 76170 343434 76226
rect 343490 76170 343558 76226
rect 343614 76170 343682 76226
rect 343738 76170 343806 76226
rect 343862 76170 343958 76226
rect 343338 76102 343958 76170
rect 343338 76046 343434 76102
rect 343490 76046 343558 76102
rect 343614 76046 343682 76102
rect 343738 76046 343806 76102
rect 343862 76046 343958 76102
rect 343338 75978 343958 76046
rect 343338 75922 343434 75978
rect 343490 75922 343558 75978
rect 343614 75922 343682 75978
rect 343738 75922 343806 75978
rect 343862 75922 343958 75978
rect 316338 64294 316434 64350
rect 316490 64294 316558 64350
rect 316614 64294 316682 64350
rect 316738 64294 316806 64350
rect 316862 64294 316958 64350
rect 316338 64226 316958 64294
rect 316338 64170 316434 64226
rect 316490 64170 316558 64226
rect 316614 64170 316682 64226
rect 316738 64170 316806 64226
rect 316862 64170 316958 64226
rect 316338 64102 316958 64170
rect 316338 64046 316434 64102
rect 316490 64046 316558 64102
rect 316614 64046 316682 64102
rect 316738 64046 316806 64102
rect 316862 64046 316958 64102
rect 316338 63978 316958 64046
rect 316338 63922 316434 63978
rect 316490 63922 316558 63978
rect 316614 63922 316682 63978
rect 316738 63922 316806 63978
rect 316862 63922 316958 63978
rect 316338 46350 316958 63922
rect 316338 46294 316434 46350
rect 316490 46294 316558 46350
rect 316614 46294 316682 46350
rect 316738 46294 316806 46350
rect 316862 46294 316958 46350
rect 316338 46226 316958 46294
rect 316338 46170 316434 46226
rect 316490 46170 316558 46226
rect 316614 46170 316682 46226
rect 316738 46170 316806 46226
rect 316862 46170 316958 46226
rect 316338 46102 316958 46170
rect 316338 46046 316434 46102
rect 316490 46046 316558 46102
rect 316614 46046 316682 46102
rect 316738 46046 316806 46102
rect 316862 46046 316958 46102
rect 316338 45978 316958 46046
rect 316338 45922 316434 45978
rect 316490 45922 316558 45978
rect 316614 45922 316682 45978
rect 316738 45922 316806 45978
rect 316862 45922 316958 45978
rect 316338 28350 316958 45922
rect 316338 28294 316434 28350
rect 316490 28294 316558 28350
rect 316614 28294 316682 28350
rect 316738 28294 316806 28350
rect 316862 28294 316958 28350
rect 316338 28226 316958 28294
rect 316338 28170 316434 28226
rect 316490 28170 316558 28226
rect 316614 28170 316682 28226
rect 316738 28170 316806 28226
rect 316862 28170 316958 28226
rect 316338 28102 316958 28170
rect 316338 28046 316434 28102
rect 316490 28046 316558 28102
rect 316614 28046 316682 28102
rect 316738 28046 316806 28102
rect 316862 28046 316958 28102
rect 316338 27978 316958 28046
rect 316338 27922 316434 27978
rect 316490 27922 316558 27978
rect 316614 27922 316682 27978
rect 316738 27922 316806 27978
rect 316862 27922 316958 27978
rect 312618 22294 312714 22350
rect 312770 22294 312838 22350
rect 312894 22294 312962 22350
rect 313018 22294 313086 22350
rect 313142 22294 313238 22350
rect 312618 22226 313238 22294
rect 312618 22170 312714 22226
rect 312770 22170 312838 22226
rect 312894 22170 312962 22226
rect 313018 22170 313086 22226
rect 313142 22170 313238 22226
rect 312618 22102 313238 22170
rect 312618 22046 312714 22102
rect 312770 22046 312838 22102
rect 312894 22046 312962 22102
rect 313018 22046 313086 22102
rect 313142 22046 313238 22102
rect 312618 21978 313238 22046
rect 312618 21922 312714 21978
rect 312770 21922 312838 21978
rect 312894 21922 312962 21978
rect 313018 21922 313086 21978
rect 313142 21922 313238 21978
rect 312618 4350 313238 21922
rect 312618 4294 312714 4350
rect 312770 4294 312838 4350
rect 312894 4294 312962 4350
rect 313018 4294 313086 4350
rect 313142 4294 313238 4350
rect 312618 4226 313238 4294
rect 312618 4170 312714 4226
rect 312770 4170 312838 4226
rect 312894 4170 312962 4226
rect 313018 4170 313086 4226
rect 313142 4170 313238 4226
rect 308364 3378 308420 3388
rect 312618 4102 313238 4170
rect 314188 22798 314244 22808
rect 314188 4228 314244 22742
rect 314188 4162 314244 4172
rect 316338 10350 316958 27922
rect 316338 10294 316434 10350
rect 316490 10294 316558 10350
rect 316614 10294 316682 10350
rect 316738 10294 316806 10350
rect 316862 10294 316958 10350
rect 316338 10226 316958 10294
rect 316338 10170 316434 10226
rect 316490 10170 316558 10226
rect 316614 10170 316682 10226
rect 316738 10170 316806 10226
rect 316862 10170 316958 10226
rect 316338 10102 316958 10170
rect 316338 10046 316434 10102
rect 316490 10046 316558 10102
rect 316614 10046 316682 10102
rect 316738 10046 316806 10102
rect 316862 10046 316958 10102
rect 316338 9978 316958 10046
rect 316338 9922 316434 9978
rect 316490 9922 316558 9978
rect 316614 9922 316682 9978
rect 316738 9922 316806 9978
rect 316862 9922 316958 9978
rect 312618 4046 312714 4102
rect 312770 4046 312838 4102
rect 312894 4046 312962 4102
rect 313018 4046 313086 4102
rect 313142 4046 313238 4102
rect 312618 3978 313238 4046
rect 312618 3922 312714 3978
rect 312770 3922 312838 3978
rect 312894 3922 312962 3978
rect 313018 3922 313086 3978
rect 313142 3922 313238 3978
rect 285618 -1176 285714 -1120
rect 285770 -1176 285838 -1120
rect 285894 -1176 285962 -1120
rect 286018 -1176 286086 -1120
rect 286142 -1176 286238 -1120
rect 285618 -1244 286238 -1176
rect 285618 -1300 285714 -1244
rect 285770 -1300 285838 -1244
rect 285894 -1300 285962 -1244
rect 286018 -1300 286086 -1244
rect 286142 -1300 286238 -1244
rect 285618 -1368 286238 -1300
rect 285618 -1424 285714 -1368
rect 285770 -1424 285838 -1368
rect 285894 -1424 285962 -1368
rect 286018 -1424 286086 -1368
rect 286142 -1424 286238 -1368
rect 285618 -1492 286238 -1424
rect 285618 -1548 285714 -1492
rect 285770 -1548 285838 -1492
rect 285894 -1548 285962 -1492
rect 286018 -1548 286086 -1492
rect 286142 -1548 286238 -1492
rect 285618 -1644 286238 -1548
rect 312618 -160 313238 3922
rect 312618 -216 312714 -160
rect 312770 -216 312838 -160
rect 312894 -216 312962 -160
rect 313018 -216 313086 -160
rect 313142 -216 313238 -160
rect 312618 -284 313238 -216
rect 312618 -340 312714 -284
rect 312770 -340 312838 -284
rect 312894 -340 312962 -284
rect 313018 -340 313086 -284
rect 313142 -340 313238 -284
rect 312618 -408 313238 -340
rect 312618 -464 312714 -408
rect 312770 -464 312838 -408
rect 312894 -464 312962 -408
rect 313018 -464 313086 -408
rect 313142 -464 313238 -408
rect 312618 -532 313238 -464
rect 312618 -588 312714 -532
rect 312770 -588 312838 -532
rect 312894 -588 312962 -532
rect 313018 -588 313086 -532
rect 313142 -588 313238 -532
rect 312618 -1644 313238 -588
rect 316338 -1120 316958 9922
rect 317548 65998 317604 66008
rect 317548 4228 317604 65942
rect 324268 62578 324324 62588
rect 322588 59518 322644 59528
rect 317548 4162 317604 4172
rect 319228 44398 319284 44408
rect 319228 4228 319284 44342
rect 319228 4162 319284 4172
rect 322588 4228 322644 59462
rect 322588 4162 322644 4172
rect 324268 4228 324324 62522
rect 343338 58350 343958 75922
rect 343338 58294 343434 58350
rect 343490 58294 343558 58350
rect 343614 58294 343682 58350
rect 343738 58294 343806 58350
rect 343862 58294 343958 58350
rect 343338 58226 343958 58294
rect 343338 58170 343434 58226
rect 343490 58170 343558 58226
rect 343614 58170 343682 58226
rect 343738 58170 343806 58226
rect 343862 58170 343958 58226
rect 343338 58102 343958 58170
rect 343338 58046 343434 58102
rect 343490 58046 343558 58102
rect 343614 58046 343682 58102
rect 343738 58046 343806 58102
rect 343862 58046 343958 58102
rect 343338 57978 343958 58046
rect 343338 57922 343434 57978
rect 343490 57922 343558 57978
rect 343614 57922 343682 57978
rect 343738 57922 343806 57978
rect 343862 57922 343958 57978
rect 330988 40798 331044 40808
rect 330988 20188 331044 40742
rect 343338 40350 343958 57922
rect 347058 598172 347678 598268
rect 347058 598116 347154 598172
rect 347210 598116 347278 598172
rect 347334 598116 347402 598172
rect 347458 598116 347526 598172
rect 347582 598116 347678 598172
rect 347058 598048 347678 598116
rect 347058 597992 347154 598048
rect 347210 597992 347278 598048
rect 347334 597992 347402 598048
rect 347458 597992 347526 598048
rect 347582 597992 347678 598048
rect 347058 597924 347678 597992
rect 347058 597868 347154 597924
rect 347210 597868 347278 597924
rect 347334 597868 347402 597924
rect 347458 597868 347526 597924
rect 347582 597868 347678 597924
rect 347058 597800 347678 597868
rect 347058 597744 347154 597800
rect 347210 597744 347278 597800
rect 347334 597744 347402 597800
rect 347458 597744 347526 597800
rect 347582 597744 347678 597800
rect 347058 586350 347678 597744
rect 347058 586294 347154 586350
rect 347210 586294 347278 586350
rect 347334 586294 347402 586350
rect 347458 586294 347526 586350
rect 347582 586294 347678 586350
rect 347058 586226 347678 586294
rect 347058 586170 347154 586226
rect 347210 586170 347278 586226
rect 347334 586170 347402 586226
rect 347458 586170 347526 586226
rect 347582 586170 347678 586226
rect 347058 586102 347678 586170
rect 347058 586046 347154 586102
rect 347210 586046 347278 586102
rect 347334 586046 347402 586102
rect 347458 586046 347526 586102
rect 347582 586046 347678 586102
rect 347058 585978 347678 586046
rect 347058 585922 347154 585978
rect 347210 585922 347278 585978
rect 347334 585922 347402 585978
rect 347458 585922 347526 585978
rect 347582 585922 347678 585978
rect 347058 568350 347678 585922
rect 347058 568294 347154 568350
rect 347210 568294 347278 568350
rect 347334 568294 347402 568350
rect 347458 568294 347526 568350
rect 347582 568294 347678 568350
rect 347058 568226 347678 568294
rect 347058 568170 347154 568226
rect 347210 568170 347278 568226
rect 347334 568170 347402 568226
rect 347458 568170 347526 568226
rect 347582 568170 347678 568226
rect 347058 568102 347678 568170
rect 347058 568046 347154 568102
rect 347210 568046 347278 568102
rect 347334 568046 347402 568102
rect 347458 568046 347526 568102
rect 347582 568046 347678 568102
rect 347058 567978 347678 568046
rect 347058 567922 347154 567978
rect 347210 567922 347278 567978
rect 347334 567922 347402 567978
rect 347458 567922 347526 567978
rect 347582 567922 347678 567978
rect 347058 550350 347678 567922
rect 347058 550294 347154 550350
rect 347210 550294 347278 550350
rect 347334 550294 347402 550350
rect 347458 550294 347526 550350
rect 347582 550294 347678 550350
rect 347058 550226 347678 550294
rect 347058 550170 347154 550226
rect 347210 550170 347278 550226
rect 347334 550170 347402 550226
rect 347458 550170 347526 550226
rect 347582 550170 347678 550226
rect 347058 550102 347678 550170
rect 347058 550046 347154 550102
rect 347210 550046 347278 550102
rect 347334 550046 347402 550102
rect 347458 550046 347526 550102
rect 347582 550046 347678 550102
rect 347058 549978 347678 550046
rect 347058 549922 347154 549978
rect 347210 549922 347278 549978
rect 347334 549922 347402 549978
rect 347458 549922 347526 549978
rect 347582 549922 347678 549978
rect 347058 532350 347678 549922
rect 347058 532294 347154 532350
rect 347210 532294 347278 532350
rect 347334 532294 347402 532350
rect 347458 532294 347526 532350
rect 347582 532294 347678 532350
rect 347058 532226 347678 532294
rect 347058 532170 347154 532226
rect 347210 532170 347278 532226
rect 347334 532170 347402 532226
rect 347458 532170 347526 532226
rect 347582 532170 347678 532226
rect 347058 532102 347678 532170
rect 347058 532046 347154 532102
rect 347210 532046 347278 532102
rect 347334 532046 347402 532102
rect 347458 532046 347526 532102
rect 347582 532046 347678 532102
rect 347058 531978 347678 532046
rect 347058 531922 347154 531978
rect 347210 531922 347278 531978
rect 347334 531922 347402 531978
rect 347458 531922 347526 531978
rect 347582 531922 347678 531978
rect 347058 514350 347678 531922
rect 347058 514294 347154 514350
rect 347210 514294 347278 514350
rect 347334 514294 347402 514350
rect 347458 514294 347526 514350
rect 347582 514294 347678 514350
rect 347058 514226 347678 514294
rect 347058 514170 347154 514226
rect 347210 514170 347278 514226
rect 347334 514170 347402 514226
rect 347458 514170 347526 514226
rect 347582 514170 347678 514226
rect 347058 514102 347678 514170
rect 347058 514046 347154 514102
rect 347210 514046 347278 514102
rect 347334 514046 347402 514102
rect 347458 514046 347526 514102
rect 347582 514046 347678 514102
rect 347058 513978 347678 514046
rect 347058 513922 347154 513978
rect 347210 513922 347278 513978
rect 347334 513922 347402 513978
rect 347458 513922 347526 513978
rect 347582 513922 347678 513978
rect 347058 496350 347678 513922
rect 347058 496294 347154 496350
rect 347210 496294 347278 496350
rect 347334 496294 347402 496350
rect 347458 496294 347526 496350
rect 347582 496294 347678 496350
rect 347058 496226 347678 496294
rect 347058 496170 347154 496226
rect 347210 496170 347278 496226
rect 347334 496170 347402 496226
rect 347458 496170 347526 496226
rect 347582 496170 347678 496226
rect 347058 496102 347678 496170
rect 347058 496046 347154 496102
rect 347210 496046 347278 496102
rect 347334 496046 347402 496102
rect 347458 496046 347526 496102
rect 347582 496046 347678 496102
rect 347058 495978 347678 496046
rect 347058 495922 347154 495978
rect 347210 495922 347278 495978
rect 347334 495922 347402 495978
rect 347458 495922 347526 495978
rect 347582 495922 347678 495978
rect 347058 478350 347678 495922
rect 347058 478294 347154 478350
rect 347210 478294 347278 478350
rect 347334 478294 347402 478350
rect 347458 478294 347526 478350
rect 347582 478294 347678 478350
rect 347058 478226 347678 478294
rect 347058 478170 347154 478226
rect 347210 478170 347278 478226
rect 347334 478170 347402 478226
rect 347458 478170 347526 478226
rect 347582 478170 347678 478226
rect 347058 478102 347678 478170
rect 347058 478046 347154 478102
rect 347210 478046 347278 478102
rect 347334 478046 347402 478102
rect 347458 478046 347526 478102
rect 347582 478046 347678 478102
rect 347058 477978 347678 478046
rect 347058 477922 347154 477978
rect 347210 477922 347278 477978
rect 347334 477922 347402 477978
rect 347458 477922 347526 477978
rect 347582 477922 347678 477978
rect 347058 460350 347678 477922
rect 347058 460294 347154 460350
rect 347210 460294 347278 460350
rect 347334 460294 347402 460350
rect 347458 460294 347526 460350
rect 347582 460294 347678 460350
rect 347058 460226 347678 460294
rect 347058 460170 347154 460226
rect 347210 460170 347278 460226
rect 347334 460170 347402 460226
rect 347458 460170 347526 460226
rect 347582 460170 347678 460226
rect 347058 460102 347678 460170
rect 347058 460046 347154 460102
rect 347210 460046 347278 460102
rect 347334 460046 347402 460102
rect 347458 460046 347526 460102
rect 347582 460046 347678 460102
rect 347058 459978 347678 460046
rect 347058 459922 347154 459978
rect 347210 459922 347278 459978
rect 347334 459922 347402 459978
rect 347458 459922 347526 459978
rect 347582 459922 347678 459978
rect 347058 442350 347678 459922
rect 347058 442294 347154 442350
rect 347210 442294 347278 442350
rect 347334 442294 347402 442350
rect 347458 442294 347526 442350
rect 347582 442294 347678 442350
rect 347058 442226 347678 442294
rect 347058 442170 347154 442226
rect 347210 442170 347278 442226
rect 347334 442170 347402 442226
rect 347458 442170 347526 442226
rect 347582 442170 347678 442226
rect 347058 442102 347678 442170
rect 347058 442046 347154 442102
rect 347210 442046 347278 442102
rect 347334 442046 347402 442102
rect 347458 442046 347526 442102
rect 347582 442046 347678 442102
rect 347058 441978 347678 442046
rect 347058 441922 347154 441978
rect 347210 441922 347278 441978
rect 347334 441922 347402 441978
rect 347458 441922 347526 441978
rect 347582 441922 347678 441978
rect 347058 424350 347678 441922
rect 347058 424294 347154 424350
rect 347210 424294 347278 424350
rect 347334 424294 347402 424350
rect 347458 424294 347526 424350
rect 347582 424294 347678 424350
rect 347058 424226 347678 424294
rect 347058 424170 347154 424226
rect 347210 424170 347278 424226
rect 347334 424170 347402 424226
rect 347458 424170 347526 424226
rect 347582 424170 347678 424226
rect 347058 424102 347678 424170
rect 347058 424046 347154 424102
rect 347210 424046 347278 424102
rect 347334 424046 347402 424102
rect 347458 424046 347526 424102
rect 347582 424046 347678 424102
rect 347058 423978 347678 424046
rect 347058 423922 347154 423978
rect 347210 423922 347278 423978
rect 347334 423922 347402 423978
rect 347458 423922 347526 423978
rect 347582 423922 347678 423978
rect 347058 406350 347678 423922
rect 347058 406294 347154 406350
rect 347210 406294 347278 406350
rect 347334 406294 347402 406350
rect 347458 406294 347526 406350
rect 347582 406294 347678 406350
rect 347058 406226 347678 406294
rect 347058 406170 347154 406226
rect 347210 406170 347278 406226
rect 347334 406170 347402 406226
rect 347458 406170 347526 406226
rect 347582 406170 347678 406226
rect 347058 406102 347678 406170
rect 347058 406046 347154 406102
rect 347210 406046 347278 406102
rect 347334 406046 347402 406102
rect 347458 406046 347526 406102
rect 347582 406046 347678 406102
rect 347058 405978 347678 406046
rect 347058 405922 347154 405978
rect 347210 405922 347278 405978
rect 347334 405922 347402 405978
rect 347458 405922 347526 405978
rect 347582 405922 347678 405978
rect 347058 388350 347678 405922
rect 347058 388294 347154 388350
rect 347210 388294 347278 388350
rect 347334 388294 347402 388350
rect 347458 388294 347526 388350
rect 347582 388294 347678 388350
rect 347058 388226 347678 388294
rect 347058 388170 347154 388226
rect 347210 388170 347278 388226
rect 347334 388170 347402 388226
rect 347458 388170 347526 388226
rect 347582 388170 347678 388226
rect 347058 388102 347678 388170
rect 347058 388046 347154 388102
rect 347210 388046 347278 388102
rect 347334 388046 347402 388102
rect 347458 388046 347526 388102
rect 347582 388046 347678 388102
rect 347058 387978 347678 388046
rect 347058 387922 347154 387978
rect 347210 387922 347278 387978
rect 347334 387922 347402 387978
rect 347458 387922 347526 387978
rect 347582 387922 347678 387978
rect 347058 370350 347678 387922
rect 347058 370294 347154 370350
rect 347210 370294 347278 370350
rect 347334 370294 347402 370350
rect 347458 370294 347526 370350
rect 347582 370294 347678 370350
rect 347058 370226 347678 370294
rect 347058 370170 347154 370226
rect 347210 370170 347278 370226
rect 347334 370170 347402 370226
rect 347458 370170 347526 370226
rect 347582 370170 347678 370226
rect 347058 370102 347678 370170
rect 347058 370046 347154 370102
rect 347210 370046 347278 370102
rect 347334 370046 347402 370102
rect 347458 370046 347526 370102
rect 347582 370046 347678 370102
rect 347058 369978 347678 370046
rect 347058 369922 347154 369978
rect 347210 369922 347278 369978
rect 347334 369922 347402 369978
rect 347458 369922 347526 369978
rect 347582 369922 347678 369978
rect 347058 352350 347678 369922
rect 347058 352294 347154 352350
rect 347210 352294 347278 352350
rect 347334 352294 347402 352350
rect 347458 352294 347526 352350
rect 347582 352294 347678 352350
rect 347058 352226 347678 352294
rect 347058 352170 347154 352226
rect 347210 352170 347278 352226
rect 347334 352170 347402 352226
rect 347458 352170 347526 352226
rect 347582 352170 347678 352226
rect 347058 352102 347678 352170
rect 347058 352046 347154 352102
rect 347210 352046 347278 352102
rect 347334 352046 347402 352102
rect 347458 352046 347526 352102
rect 347582 352046 347678 352102
rect 347058 351978 347678 352046
rect 347058 351922 347154 351978
rect 347210 351922 347278 351978
rect 347334 351922 347402 351978
rect 347458 351922 347526 351978
rect 347582 351922 347678 351978
rect 347058 334350 347678 351922
rect 347058 334294 347154 334350
rect 347210 334294 347278 334350
rect 347334 334294 347402 334350
rect 347458 334294 347526 334350
rect 347582 334294 347678 334350
rect 347058 334226 347678 334294
rect 347058 334170 347154 334226
rect 347210 334170 347278 334226
rect 347334 334170 347402 334226
rect 347458 334170 347526 334226
rect 347582 334170 347678 334226
rect 347058 334102 347678 334170
rect 347058 334046 347154 334102
rect 347210 334046 347278 334102
rect 347334 334046 347402 334102
rect 347458 334046 347526 334102
rect 347582 334046 347678 334102
rect 347058 333978 347678 334046
rect 347058 333922 347154 333978
rect 347210 333922 347278 333978
rect 347334 333922 347402 333978
rect 347458 333922 347526 333978
rect 347582 333922 347678 333978
rect 347058 316350 347678 333922
rect 347058 316294 347154 316350
rect 347210 316294 347278 316350
rect 347334 316294 347402 316350
rect 347458 316294 347526 316350
rect 347582 316294 347678 316350
rect 347058 316226 347678 316294
rect 347058 316170 347154 316226
rect 347210 316170 347278 316226
rect 347334 316170 347402 316226
rect 347458 316170 347526 316226
rect 347582 316170 347678 316226
rect 347058 316102 347678 316170
rect 347058 316046 347154 316102
rect 347210 316046 347278 316102
rect 347334 316046 347402 316102
rect 347458 316046 347526 316102
rect 347582 316046 347678 316102
rect 347058 315978 347678 316046
rect 347058 315922 347154 315978
rect 347210 315922 347278 315978
rect 347334 315922 347402 315978
rect 347458 315922 347526 315978
rect 347582 315922 347678 315978
rect 347058 298350 347678 315922
rect 347058 298294 347154 298350
rect 347210 298294 347278 298350
rect 347334 298294 347402 298350
rect 347458 298294 347526 298350
rect 347582 298294 347678 298350
rect 347058 298226 347678 298294
rect 347058 298170 347154 298226
rect 347210 298170 347278 298226
rect 347334 298170 347402 298226
rect 347458 298170 347526 298226
rect 347582 298170 347678 298226
rect 347058 298102 347678 298170
rect 347058 298046 347154 298102
rect 347210 298046 347278 298102
rect 347334 298046 347402 298102
rect 347458 298046 347526 298102
rect 347582 298046 347678 298102
rect 347058 297978 347678 298046
rect 347058 297922 347154 297978
rect 347210 297922 347278 297978
rect 347334 297922 347402 297978
rect 347458 297922 347526 297978
rect 347582 297922 347678 297978
rect 347058 280350 347678 297922
rect 347058 280294 347154 280350
rect 347210 280294 347278 280350
rect 347334 280294 347402 280350
rect 347458 280294 347526 280350
rect 347582 280294 347678 280350
rect 347058 280226 347678 280294
rect 347058 280170 347154 280226
rect 347210 280170 347278 280226
rect 347334 280170 347402 280226
rect 347458 280170 347526 280226
rect 347582 280170 347678 280226
rect 347058 280102 347678 280170
rect 347058 280046 347154 280102
rect 347210 280046 347278 280102
rect 347334 280046 347402 280102
rect 347458 280046 347526 280102
rect 347582 280046 347678 280102
rect 347058 279978 347678 280046
rect 347058 279922 347154 279978
rect 347210 279922 347278 279978
rect 347334 279922 347402 279978
rect 347458 279922 347526 279978
rect 347582 279922 347678 279978
rect 347058 262350 347678 279922
rect 347058 262294 347154 262350
rect 347210 262294 347278 262350
rect 347334 262294 347402 262350
rect 347458 262294 347526 262350
rect 347582 262294 347678 262350
rect 347058 262226 347678 262294
rect 347058 262170 347154 262226
rect 347210 262170 347278 262226
rect 347334 262170 347402 262226
rect 347458 262170 347526 262226
rect 347582 262170 347678 262226
rect 347058 262102 347678 262170
rect 347058 262046 347154 262102
rect 347210 262046 347278 262102
rect 347334 262046 347402 262102
rect 347458 262046 347526 262102
rect 347582 262046 347678 262102
rect 347058 261978 347678 262046
rect 347058 261922 347154 261978
rect 347210 261922 347278 261978
rect 347334 261922 347402 261978
rect 347458 261922 347526 261978
rect 347582 261922 347678 261978
rect 347058 244350 347678 261922
rect 347058 244294 347154 244350
rect 347210 244294 347278 244350
rect 347334 244294 347402 244350
rect 347458 244294 347526 244350
rect 347582 244294 347678 244350
rect 347058 244226 347678 244294
rect 347058 244170 347154 244226
rect 347210 244170 347278 244226
rect 347334 244170 347402 244226
rect 347458 244170 347526 244226
rect 347582 244170 347678 244226
rect 347058 244102 347678 244170
rect 347058 244046 347154 244102
rect 347210 244046 347278 244102
rect 347334 244046 347402 244102
rect 347458 244046 347526 244102
rect 347582 244046 347678 244102
rect 347058 243978 347678 244046
rect 347058 243922 347154 243978
rect 347210 243922 347278 243978
rect 347334 243922 347402 243978
rect 347458 243922 347526 243978
rect 347582 243922 347678 243978
rect 347058 226350 347678 243922
rect 347058 226294 347154 226350
rect 347210 226294 347278 226350
rect 347334 226294 347402 226350
rect 347458 226294 347526 226350
rect 347582 226294 347678 226350
rect 347058 226226 347678 226294
rect 347058 226170 347154 226226
rect 347210 226170 347278 226226
rect 347334 226170 347402 226226
rect 347458 226170 347526 226226
rect 347582 226170 347678 226226
rect 347058 226102 347678 226170
rect 347058 226046 347154 226102
rect 347210 226046 347278 226102
rect 347334 226046 347402 226102
rect 347458 226046 347526 226102
rect 347582 226046 347678 226102
rect 347058 225978 347678 226046
rect 347058 225922 347154 225978
rect 347210 225922 347278 225978
rect 347334 225922 347402 225978
rect 347458 225922 347526 225978
rect 347582 225922 347678 225978
rect 347058 208350 347678 225922
rect 347058 208294 347154 208350
rect 347210 208294 347278 208350
rect 347334 208294 347402 208350
rect 347458 208294 347526 208350
rect 347582 208294 347678 208350
rect 347058 208226 347678 208294
rect 347058 208170 347154 208226
rect 347210 208170 347278 208226
rect 347334 208170 347402 208226
rect 347458 208170 347526 208226
rect 347582 208170 347678 208226
rect 347058 208102 347678 208170
rect 347058 208046 347154 208102
rect 347210 208046 347278 208102
rect 347334 208046 347402 208102
rect 347458 208046 347526 208102
rect 347582 208046 347678 208102
rect 347058 207978 347678 208046
rect 347058 207922 347154 207978
rect 347210 207922 347278 207978
rect 347334 207922 347402 207978
rect 347458 207922 347526 207978
rect 347582 207922 347678 207978
rect 347058 190350 347678 207922
rect 347058 190294 347154 190350
rect 347210 190294 347278 190350
rect 347334 190294 347402 190350
rect 347458 190294 347526 190350
rect 347582 190294 347678 190350
rect 347058 190226 347678 190294
rect 347058 190170 347154 190226
rect 347210 190170 347278 190226
rect 347334 190170 347402 190226
rect 347458 190170 347526 190226
rect 347582 190170 347678 190226
rect 347058 190102 347678 190170
rect 347058 190046 347154 190102
rect 347210 190046 347278 190102
rect 347334 190046 347402 190102
rect 347458 190046 347526 190102
rect 347582 190046 347678 190102
rect 347058 189978 347678 190046
rect 347058 189922 347154 189978
rect 347210 189922 347278 189978
rect 347334 189922 347402 189978
rect 347458 189922 347526 189978
rect 347582 189922 347678 189978
rect 347058 172350 347678 189922
rect 347058 172294 347154 172350
rect 347210 172294 347278 172350
rect 347334 172294 347402 172350
rect 347458 172294 347526 172350
rect 347582 172294 347678 172350
rect 347058 172226 347678 172294
rect 347058 172170 347154 172226
rect 347210 172170 347278 172226
rect 347334 172170 347402 172226
rect 347458 172170 347526 172226
rect 347582 172170 347678 172226
rect 347058 172102 347678 172170
rect 347058 172046 347154 172102
rect 347210 172046 347278 172102
rect 347334 172046 347402 172102
rect 347458 172046 347526 172102
rect 347582 172046 347678 172102
rect 347058 171978 347678 172046
rect 347058 171922 347154 171978
rect 347210 171922 347278 171978
rect 347334 171922 347402 171978
rect 347458 171922 347526 171978
rect 347582 171922 347678 171978
rect 347058 154350 347678 171922
rect 347058 154294 347154 154350
rect 347210 154294 347278 154350
rect 347334 154294 347402 154350
rect 347458 154294 347526 154350
rect 347582 154294 347678 154350
rect 347058 154226 347678 154294
rect 347058 154170 347154 154226
rect 347210 154170 347278 154226
rect 347334 154170 347402 154226
rect 347458 154170 347526 154226
rect 347582 154170 347678 154226
rect 347058 154102 347678 154170
rect 347058 154046 347154 154102
rect 347210 154046 347278 154102
rect 347334 154046 347402 154102
rect 347458 154046 347526 154102
rect 347582 154046 347678 154102
rect 347058 153978 347678 154046
rect 347058 153922 347154 153978
rect 347210 153922 347278 153978
rect 347334 153922 347402 153978
rect 347458 153922 347526 153978
rect 347582 153922 347678 153978
rect 347058 136350 347678 153922
rect 347058 136294 347154 136350
rect 347210 136294 347278 136350
rect 347334 136294 347402 136350
rect 347458 136294 347526 136350
rect 347582 136294 347678 136350
rect 347058 136226 347678 136294
rect 347058 136170 347154 136226
rect 347210 136170 347278 136226
rect 347334 136170 347402 136226
rect 347458 136170 347526 136226
rect 347582 136170 347678 136226
rect 347058 136102 347678 136170
rect 347058 136046 347154 136102
rect 347210 136046 347278 136102
rect 347334 136046 347402 136102
rect 347458 136046 347526 136102
rect 347582 136046 347678 136102
rect 347058 135978 347678 136046
rect 347058 135922 347154 135978
rect 347210 135922 347278 135978
rect 347334 135922 347402 135978
rect 347458 135922 347526 135978
rect 347582 135922 347678 135978
rect 347058 118350 347678 135922
rect 347058 118294 347154 118350
rect 347210 118294 347278 118350
rect 347334 118294 347402 118350
rect 347458 118294 347526 118350
rect 347582 118294 347678 118350
rect 347058 118226 347678 118294
rect 347058 118170 347154 118226
rect 347210 118170 347278 118226
rect 347334 118170 347402 118226
rect 347458 118170 347526 118226
rect 347582 118170 347678 118226
rect 347058 118102 347678 118170
rect 347058 118046 347154 118102
rect 347210 118046 347278 118102
rect 347334 118046 347402 118102
rect 347458 118046 347526 118102
rect 347582 118046 347678 118102
rect 347058 117978 347678 118046
rect 347058 117922 347154 117978
rect 347210 117922 347278 117978
rect 347334 117922 347402 117978
rect 347458 117922 347526 117978
rect 347582 117922 347678 117978
rect 347058 100350 347678 117922
rect 347058 100294 347154 100350
rect 347210 100294 347278 100350
rect 347334 100294 347402 100350
rect 347458 100294 347526 100350
rect 347582 100294 347678 100350
rect 347058 100226 347678 100294
rect 347058 100170 347154 100226
rect 347210 100170 347278 100226
rect 347334 100170 347402 100226
rect 347458 100170 347526 100226
rect 347582 100170 347678 100226
rect 347058 100102 347678 100170
rect 347058 100046 347154 100102
rect 347210 100046 347278 100102
rect 347334 100046 347402 100102
rect 347458 100046 347526 100102
rect 347582 100046 347678 100102
rect 347058 99978 347678 100046
rect 347058 99922 347154 99978
rect 347210 99922 347278 99978
rect 347334 99922 347402 99978
rect 347458 99922 347526 99978
rect 347582 99922 347678 99978
rect 347058 82350 347678 99922
rect 347058 82294 347154 82350
rect 347210 82294 347278 82350
rect 347334 82294 347402 82350
rect 347458 82294 347526 82350
rect 347582 82294 347678 82350
rect 347058 82226 347678 82294
rect 347058 82170 347154 82226
rect 347210 82170 347278 82226
rect 347334 82170 347402 82226
rect 347458 82170 347526 82226
rect 347582 82170 347678 82226
rect 347058 82102 347678 82170
rect 347058 82046 347154 82102
rect 347210 82046 347278 82102
rect 347334 82046 347402 82102
rect 347458 82046 347526 82102
rect 347582 82046 347678 82102
rect 347058 81978 347678 82046
rect 347058 81922 347154 81978
rect 347210 81922 347278 81978
rect 347334 81922 347402 81978
rect 347458 81922 347526 81978
rect 347582 81922 347678 81978
rect 347058 64350 347678 81922
rect 347058 64294 347154 64350
rect 347210 64294 347278 64350
rect 347334 64294 347402 64350
rect 347458 64294 347526 64350
rect 347582 64294 347678 64350
rect 347058 64226 347678 64294
rect 347058 64170 347154 64226
rect 347210 64170 347278 64226
rect 347334 64170 347402 64226
rect 347458 64170 347526 64226
rect 347582 64170 347678 64226
rect 347058 64102 347678 64170
rect 347058 64046 347154 64102
rect 347210 64046 347278 64102
rect 347334 64046 347402 64102
rect 347458 64046 347526 64102
rect 347582 64046 347678 64102
rect 347058 63978 347678 64046
rect 347058 63922 347154 63978
rect 347210 63922 347278 63978
rect 347334 63922 347402 63978
rect 347458 63922 347526 63978
rect 347582 63922 347678 63978
rect 347058 46350 347678 63922
rect 347058 46294 347154 46350
rect 347210 46294 347278 46350
rect 347334 46294 347402 46350
rect 347458 46294 347526 46350
rect 347582 46294 347678 46350
rect 347058 46226 347678 46294
rect 347058 46170 347154 46226
rect 347210 46170 347278 46226
rect 347334 46170 347402 46226
rect 347458 46170 347526 46226
rect 347582 46170 347678 46226
rect 347058 46102 347678 46170
rect 347058 46046 347154 46102
rect 347210 46046 347278 46102
rect 347334 46046 347402 46102
rect 347458 46046 347526 46102
rect 347582 46046 347678 46102
rect 347058 45978 347678 46046
rect 347058 45922 347154 45978
rect 347210 45922 347278 45978
rect 347334 45922 347402 45978
rect 347458 45922 347526 45978
rect 347582 45922 347678 45978
rect 343338 40294 343434 40350
rect 343490 40294 343558 40350
rect 343614 40294 343682 40350
rect 343738 40294 343806 40350
rect 343862 40294 343958 40350
rect 343338 40226 343958 40294
rect 343338 40170 343434 40226
rect 343490 40170 343558 40226
rect 343614 40170 343682 40226
rect 343738 40170 343806 40226
rect 343862 40170 343958 40226
rect 343338 40102 343958 40170
rect 343338 40046 343434 40102
rect 343490 40046 343558 40102
rect 343614 40046 343682 40102
rect 343738 40046 343806 40102
rect 343862 40046 343958 40102
rect 343338 39978 343958 40046
rect 343338 39922 343434 39978
rect 343490 39922 343558 39978
rect 343614 39922 343682 39978
rect 343738 39922 343806 39978
rect 343862 39922 343958 39978
rect 342748 30718 342804 30728
rect 339388 30538 339444 30548
rect 330988 20132 331268 20188
rect 324268 4162 324324 4172
rect 331212 4228 331268 20132
rect 331212 4162 331268 4172
rect 336028 17218 336084 17228
rect 336028 4228 336084 17162
rect 336028 4162 336084 4172
rect 339388 4228 339444 30482
rect 339388 4162 339444 4172
rect 342748 4228 342804 30662
rect 342748 4162 342804 4172
rect 343338 22350 343958 39922
rect 343338 22294 343434 22350
rect 343490 22294 343558 22350
rect 343614 22294 343682 22350
rect 343738 22294 343806 22350
rect 343862 22294 343958 22350
rect 343338 22226 343958 22294
rect 343338 22170 343434 22226
rect 343490 22170 343558 22226
rect 343614 22170 343682 22226
rect 343738 22170 343806 22226
rect 343862 22170 343958 22226
rect 343338 22102 343958 22170
rect 343338 22046 343434 22102
rect 343490 22046 343558 22102
rect 343614 22046 343682 22102
rect 343738 22046 343806 22102
rect 343862 22046 343958 22102
rect 343338 21978 343958 22046
rect 343338 21922 343434 21978
rect 343490 21922 343558 21978
rect 343614 21922 343682 21978
rect 343738 21922 343806 21978
rect 343862 21922 343958 21978
rect 343338 4350 343958 21922
rect 343338 4294 343434 4350
rect 343490 4294 343558 4350
rect 343614 4294 343682 4350
rect 343738 4294 343806 4350
rect 343862 4294 343958 4350
rect 343338 4226 343958 4294
rect 343338 4170 343434 4226
rect 343490 4170 343558 4226
rect 343614 4170 343682 4226
rect 343738 4170 343806 4226
rect 343862 4170 343958 4226
rect 316338 -1176 316434 -1120
rect 316490 -1176 316558 -1120
rect 316614 -1176 316682 -1120
rect 316738 -1176 316806 -1120
rect 316862 -1176 316958 -1120
rect 316338 -1244 316958 -1176
rect 316338 -1300 316434 -1244
rect 316490 -1300 316558 -1244
rect 316614 -1300 316682 -1244
rect 316738 -1300 316806 -1244
rect 316862 -1300 316958 -1244
rect 316338 -1368 316958 -1300
rect 316338 -1424 316434 -1368
rect 316490 -1424 316558 -1368
rect 316614 -1424 316682 -1368
rect 316738 -1424 316806 -1368
rect 316862 -1424 316958 -1368
rect 316338 -1492 316958 -1424
rect 316338 -1548 316434 -1492
rect 316490 -1548 316558 -1492
rect 316614 -1548 316682 -1492
rect 316738 -1548 316806 -1492
rect 316862 -1548 316958 -1492
rect 316338 -1644 316958 -1548
rect 343338 4102 343958 4170
rect 346108 42778 346164 42788
rect 346108 4228 346164 42722
rect 346108 4162 346164 4172
rect 347058 28350 347678 45922
rect 374058 597212 374678 598268
rect 374058 597156 374154 597212
rect 374210 597156 374278 597212
rect 374334 597156 374402 597212
rect 374458 597156 374526 597212
rect 374582 597156 374678 597212
rect 374058 597088 374678 597156
rect 374058 597032 374154 597088
rect 374210 597032 374278 597088
rect 374334 597032 374402 597088
rect 374458 597032 374526 597088
rect 374582 597032 374678 597088
rect 374058 596964 374678 597032
rect 374058 596908 374154 596964
rect 374210 596908 374278 596964
rect 374334 596908 374402 596964
rect 374458 596908 374526 596964
rect 374582 596908 374678 596964
rect 374058 596840 374678 596908
rect 374058 596784 374154 596840
rect 374210 596784 374278 596840
rect 374334 596784 374402 596840
rect 374458 596784 374526 596840
rect 374582 596784 374678 596840
rect 374058 580350 374678 596784
rect 374058 580294 374154 580350
rect 374210 580294 374278 580350
rect 374334 580294 374402 580350
rect 374458 580294 374526 580350
rect 374582 580294 374678 580350
rect 374058 580226 374678 580294
rect 374058 580170 374154 580226
rect 374210 580170 374278 580226
rect 374334 580170 374402 580226
rect 374458 580170 374526 580226
rect 374582 580170 374678 580226
rect 374058 580102 374678 580170
rect 374058 580046 374154 580102
rect 374210 580046 374278 580102
rect 374334 580046 374402 580102
rect 374458 580046 374526 580102
rect 374582 580046 374678 580102
rect 374058 579978 374678 580046
rect 374058 579922 374154 579978
rect 374210 579922 374278 579978
rect 374334 579922 374402 579978
rect 374458 579922 374526 579978
rect 374582 579922 374678 579978
rect 374058 562350 374678 579922
rect 374058 562294 374154 562350
rect 374210 562294 374278 562350
rect 374334 562294 374402 562350
rect 374458 562294 374526 562350
rect 374582 562294 374678 562350
rect 374058 562226 374678 562294
rect 374058 562170 374154 562226
rect 374210 562170 374278 562226
rect 374334 562170 374402 562226
rect 374458 562170 374526 562226
rect 374582 562170 374678 562226
rect 374058 562102 374678 562170
rect 374058 562046 374154 562102
rect 374210 562046 374278 562102
rect 374334 562046 374402 562102
rect 374458 562046 374526 562102
rect 374582 562046 374678 562102
rect 374058 561978 374678 562046
rect 374058 561922 374154 561978
rect 374210 561922 374278 561978
rect 374334 561922 374402 561978
rect 374458 561922 374526 561978
rect 374582 561922 374678 561978
rect 374058 544350 374678 561922
rect 374058 544294 374154 544350
rect 374210 544294 374278 544350
rect 374334 544294 374402 544350
rect 374458 544294 374526 544350
rect 374582 544294 374678 544350
rect 374058 544226 374678 544294
rect 374058 544170 374154 544226
rect 374210 544170 374278 544226
rect 374334 544170 374402 544226
rect 374458 544170 374526 544226
rect 374582 544170 374678 544226
rect 374058 544102 374678 544170
rect 374058 544046 374154 544102
rect 374210 544046 374278 544102
rect 374334 544046 374402 544102
rect 374458 544046 374526 544102
rect 374582 544046 374678 544102
rect 374058 543978 374678 544046
rect 374058 543922 374154 543978
rect 374210 543922 374278 543978
rect 374334 543922 374402 543978
rect 374458 543922 374526 543978
rect 374582 543922 374678 543978
rect 374058 526350 374678 543922
rect 374058 526294 374154 526350
rect 374210 526294 374278 526350
rect 374334 526294 374402 526350
rect 374458 526294 374526 526350
rect 374582 526294 374678 526350
rect 374058 526226 374678 526294
rect 374058 526170 374154 526226
rect 374210 526170 374278 526226
rect 374334 526170 374402 526226
rect 374458 526170 374526 526226
rect 374582 526170 374678 526226
rect 374058 526102 374678 526170
rect 374058 526046 374154 526102
rect 374210 526046 374278 526102
rect 374334 526046 374402 526102
rect 374458 526046 374526 526102
rect 374582 526046 374678 526102
rect 374058 525978 374678 526046
rect 374058 525922 374154 525978
rect 374210 525922 374278 525978
rect 374334 525922 374402 525978
rect 374458 525922 374526 525978
rect 374582 525922 374678 525978
rect 374058 508350 374678 525922
rect 374058 508294 374154 508350
rect 374210 508294 374278 508350
rect 374334 508294 374402 508350
rect 374458 508294 374526 508350
rect 374582 508294 374678 508350
rect 374058 508226 374678 508294
rect 374058 508170 374154 508226
rect 374210 508170 374278 508226
rect 374334 508170 374402 508226
rect 374458 508170 374526 508226
rect 374582 508170 374678 508226
rect 374058 508102 374678 508170
rect 374058 508046 374154 508102
rect 374210 508046 374278 508102
rect 374334 508046 374402 508102
rect 374458 508046 374526 508102
rect 374582 508046 374678 508102
rect 374058 507978 374678 508046
rect 374058 507922 374154 507978
rect 374210 507922 374278 507978
rect 374334 507922 374402 507978
rect 374458 507922 374526 507978
rect 374582 507922 374678 507978
rect 374058 490350 374678 507922
rect 374058 490294 374154 490350
rect 374210 490294 374278 490350
rect 374334 490294 374402 490350
rect 374458 490294 374526 490350
rect 374582 490294 374678 490350
rect 374058 490226 374678 490294
rect 374058 490170 374154 490226
rect 374210 490170 374278 490226
rect 374334 490170 374402 490226
rect 374458 490170 374526 490226
rect 374582 490170 374678 490226
rect 374058 490102 374678 490170
rect 374058 490046 374154 490102
rect 374210 490046 374278 490102
rect 374334 490046 374402 490102
rect 374458 490046 374526 490102
rect 374582 490046 374678 490102
rect 374058 489978 374678 490046
rect 374058 489922 374154 489978
rect 374210 489922 374278 489978
rect 374334 489922 374402 489978
rect 374458 489922 374526 489978
rect 374582 489922 374678 489978
rect 374058 472350 374678 489922
rect 374058 472294 374154 472350
rect 374210 472294 374278 472350
rect 374334 472294 374402 472350
rect 374458 472294 374526 472350
rect 374582 472294 374678 472350
rect 374058 472226 374678 472294
rect 374058 472170 374154 472226
rect 374210 472170 374278 472226
rect 374334 472170 374402 472226
rect 374458 472170 374526 472226
rect 374582 472170 374678 472226
rect 374058 472102 374678 472170
rect 374058 472046 374154 472102
rect 374210 472046 374278 472102
rect 374334 472046 374402 472102
rect 374458 472046 374526 472102
rect 374582 472046 374678 472102
rect 374058 471978 374678 472046
rect 374058 471922 374154 471978
rect 374210 471922 374278 471978
rect 374334 471922 374402 471978
rect 374458 471922 374526 471978
rect 374582 471922 374678 471978
rect 374058 454350 374678 471922
rect 374058 454294 374154 454350
rect 374210 454294 374278 454350
rect 374334 454294 374402 454350
rect 374458 454294 374526 454350
rect 374582 454294 374678 454350
rect 374058 454226 374678 454294
rect 374058 454170 374154 454226
rect 374210 454170 374278 454226
rect 374334 454170 374402 454226
rect 374458 454170 374526 454226
rect 374582 454170 374678 454226
rect 374058 454102 374678 454170
rect 374058 454046 374154 454102
rect 374210 454046 374278 454102
rect 374334 454046 374402 454102
rect 374458 454046 374526 454102
rect 374582 454046 374678 454102
rect 374058 453978 374678 454046
rect 374058 453922 374154 453978
rect 374210 453922 374278 453978
rect 374334 453922 374402 453978
rect 374458 453922 374526 453978
rect 374582 453922 374678 453978
rect 374058 436350 374678 453922
rect 374058 436294 374154 436350
rect 374210 436294 374278 436350
rect 374334 436294 374402 436350
rect 374458 436294 374526 436350
rect 374582 436294 374678 436350
rect 374058 436226 374678 436294
rect 374058 436170 374154 436226
rect 374210 436170 374278 436226
rect 374334 436170 374402 436226
rect 374458 436170 374526 436226
rect 374582 436170 374678 436226
rect 374058 436102 374678 436170
rect 374058 436046 374154 436102
rect 374210 436046 374278 436102
rect 374334 436046 374402 436102
rect 374458 436046 374526 436102
rect 374582 436046 374678 436102
rect 374058 435978 374678 436046
rect 374058 435922 374154 435978
rect 374210 435922 374278 435978
rect 374334 435922 374402 435978
rect 374458 435922 374526 435978
rect 374582 435922 374678 435978
rect 374058 418350 374678 435922
rect 374058 418294 374154 418350
rect 374210 418294 374278 418350
rect 374334 418294 374402 418350
rect 374458 418294 374526 418350
rect 374582 418294 374678 418350
rect 374058 418226 374678 418294
rect 374058 418170 374154 418226
rect 374210 418170 374278 418226
rect 374334 418170 374402 418226
rect 374458 418170 374526 418226
rect 374582 418170 374678 418226
rect 374058 418102 374678 418170
rect 374058 418046 374154 418102
rect 374210 418046 374278 418102
rect 374334 418046 374402 418102
rect 374458 418046 374526 418102
rect 374582 418046 374678 418102
rect 374058 417978 374678 418046
rect 374058 417922 374154 417978
rect 374210 417922 374278 417978
rect 374334 417922 374402 417978
rect 374458 417922 374526 417978
rect 374582 417922 374678 417978
rect 374058 400350 374678 417922
rect 374058 400294 374154 400350
rect 374210 400294 374278 400350
rect 374334 400294 374402 400350
rect 374458 400294 374526 400350
rect 374582 400294 374678 400350
rect 374058 400226 374678 400294
rect 374058 400170 374154 400226
rect 374210 400170 374278 400226
rect 374334 400170 374402 400226
rect 374458 400170 374526 400226
rect 374582 400170 374678 400226
rect 374058 400102 374678 400170
rect 374058 400046 374154 400102
rect 374210 400046 374278 400102
rect 374334 400046 374402 400102
rect 374458 400046 374526 400102
rect 374582 400046 374678 400102
rect 374058 399978 374678 400046
rect 374058 399922 374154 399978
rect 374210 399922 374278 399978
rect 374334 399922 374402 399978
rect 374458 399922 374526 399978
rect 374582 399922 374678 399978
rect 374058 382350 374678 399922
rect 374058 382294 374154 382350
rect 374210 382294 374278 382350
rect 374334 382294 374402 382350
rect 374458 382294 374526 382350
rect 374582 382294 374678 382350
rect 374058 382226 374678 382294
rect 374058 382170 374154 382226
rect 374210 382170 374278 382226
rect 374334 382170 374402 382226
rect 374458 382170 374526 382226
rect 374582 382170 374678 382226
rect 374058 382102 374678 382170
rect 374058 382046 374154 382102
rect 374210 382046 374278 382102
rect 374334 382046 374402 382102
rect 374458 382046 374526 382102
rect 374582 382046 374678 382102
rect 374058 381978 374678 382046
rect 374058 381922 374154 381978
rect 374210 381922 374278 381978
rect 374334 381922 374402 381978
rect 374458 381922 374526 381978
rect 374582 381922 374678 381978
rect 374058 364350 374678 381922
rect 374058 364294 374154 364350
rect 374210 364294 374278 364350
rect 374334 364294 374402 364350
rect 374458 364294 374526 364350
rect 374582 364294 374678 364350
rect 374058 364226 374678 364294
rect 374058 364170 374154 364226
rect 374210 364170 374278 364226
rect 374334 364170 374402 364226
rect 374458 364170 374526 364226
rect 374582 364170 374678 364226
rect 374058 364102 374678 364170
rect 374058 364046 374154 364102
rect 374210 364046 374278 364102
rect 374334 364046 374402 364102
rect 374458 364046 374526 364102
rect 374582 364046 374678 364102
rect 374058 363978 374678 364046
rect 374058 363922 374154 363978
rect 374210 363922 374278 363978
rect 374334 363922 374402 363978
rect 374458 363922 374526 363978
rect 374582 363922 374678 363978
rect 374058 346350 374678 363922
rect 374058 346294 374154 346350
rect 374210 346294 374278 346350
rect 374334 346294 374402 346350
rect 374458 346294 374526 346350
rect 374582 346294 374678 346350
rect 374058 346226 374678 346294
rect 374058 346170 374154 346226
rect 374210 346170 374278 346226
rect 374334 346170 374402 346226
rect 374458 346170 374526 346226
rect 374582 346170 374678 346226
rect 374058 346102 374678 346170
rect 374058 346046 374154 346102
rect 374210 346046 374278 346102
rect 374334 346046 374402 346102
rect 374458 346046 374526 346102
rect 374582 346046 374678 346102
rect 374058 345978 374678 346046
rect 374058 345922 374154 345978
rect 374210 345922 374278 345978
rect 374334 345922 374402 345978
rect 374458 345922 374526 345978
rect 374582 345922 374678 345978
rect 374058 328350 374678 345922
rect 374058 328294 374154 328350
rect 374210 328294 374278 328350
rect 374334 328294 374402 328350
rect 374458 328294 374526 328350
rect 374582 328294 374678 328350
rect 374058 328226 374678 328294
rect 374058 328170 374154 328226
rect 374210 328170 374278 328226
rect 374334 328170 374402 328226
rect 374458 328170 374526 328226
rect 374582 328170 374678 328226
rect 374058 328102 374678 328170
rect 374058 328046 374154 328102
rect 374210 328046 374278 328102
rect 374334 328046 374402 328102
rect 374458 328046 374526 328102
rect 374582 328046 374678 328102
rect 374058 327978 374678 328046
rect 374058 327922 374154 327978
rect 374210 327922 374278 327978
rect 374334 327922 374402 327978
rect 374458 327922 374526 327978
rect 374582 327922 374678 327978
rect 374058 310350 374678 327922
rect 374058 310294 374154 310350
rect 374210 310294 374278 310350
rect 374334 310294 374402 310350
rect 374458 310294 374526 310350
rect 374582 310294 374678 310350
rect 374058 310226 374678 310294
rect 374058 310170 374154 310226
rect 374210 310170 374278 310226
rect 374334 310170 374402 310226
rect 374458 310170 374526 310226
rect 374582 310170 374678 310226
rect 374058 310102 374678 310170
rect 374058 310046 374154 310102
rect 374210 310046 374278 310102
rect 374334 310046 374402 310102
rect 374458 310046 374526 310102
rect 374582 310046 374678 310102
rect 374058 309978 374678 310046
rect 374058 309922 374154 309978
rect 374210 309922 374278 309978
rect 374334 309922 374402 309978
rect 374458 309922 374526 309978
rect 374582 309922 374678 309978
rect 374058 292350 374678 309922
rect 374058 292294 374154 292350
rect 374210 292294 374278 292350
rect 374334 292294 374402 292350
rect 374458 292294 374526 292350
rect 374582 292294 374678 292350
rect 374058 292226 374678 292294
rect 374058 292170 374154 292226
rect 374210 292170 374278 292226
rect 374334 292170 374402 292226
rect 374458 292170 374526 292226
rect 374582 292170 374678 292226
rect 374058 292102 374678 292170
rect 374058 292046 374154 292102
rect 374210 292046 374278 292102
rect 374334 292046 374402 292102
rect 374458 292046 374526 292102
rect 374582 292046 374678 292102
rect 374058 291978 374678 292046
rect 374058 291922 374154 291978
rect 374210 291922 374278 291978
rect 374334 291922 374402 291978
rect 374458 291922 374526 291978
rect 374582 291922 374678 291978
rect 374058 274350 374678 291922
rect 374058 274294 374154 274350
rect 374210 274294 374278 274350
rect 374334 274294 374402 274350
rect 374458 274294 374526 274350
rect 374582 274294 374678 274350
rect 374058 274226 374678 274294
rect 374058 274170 374154 274226
rect 374210 274170 374278 274226
rect 374334 274170 374402 274226
rect 374458 274170 374526 274226
rect 374582 274170 374678 274226
rect 374058 274102 374678 274170
rect 374058 274046 374154 274102
rect 374210 274046 374278 274102
rect 374334 274046 374402 274102
rect 374458 274046 374526 274102
rect 374582 274046 374678 274102
rect 374058 273978 374678 274046
rect 374058 273922 374154 273978
rect 374210 273922 374278 273978
rect 374334 273922 374402 273978
rect 374458 273922 374526 273978
rect 374582 273922 374678 273978
rect 374058 256350 374678 273922
rect 374058 256294 374154 256350
rect 374210 256294 374278 256350
rect 374334 256294 374402 256350
rect 374458 256294 374526 256350
rect 374582 256294 374678 256350
rect 374058 256226 374678 256294
rect 374058 256170 374154 256226
rect 374210 256170 374278 256226
rect 374334 256170 374402 256226
rect 374458 256170 374526 256226
rect 374582 256170 374678 256226
rect 374058 256102 374678 256170
rect 374058 256046 374154 256102
rect 374210 256046 374278 256102
rect 374334 256046 374402 256102
rect 374458 256046 374526 256102
rect 374582 256046 374678 256102
rect 374058 255978 374678 256046
rect 374058 255922 374154 255978
rect 374210 255922 374278 255978
rect 374334 255922 374402 255978
rect 374458 255922 374526 255978
rect 374582 255922 374678 255978
rect 374058 238350 374678 255922
rect 374058 238294 374154 238350
rect 374210 238294 374278 238350
rect 374334 238294 374402 238350
rect 374458 238294 374526 238350
rect 374582 238294 374678 238350
rect 374058 238226 374678 238294
rect 374058 238170 374154 238226
rect 374210 238170 374278 238226
rect 374334 238170 374402 238226
rect 374458 238170 374526 238226
rect 374582 238170 374678 238226
rect 374058 238102 374678 238170
rect 374058 238046 374154 238102
rect 374210 238046 374278 238102
rect 374334 238046 374402 238102
rect 374458 238046 374526 238102
rect 374582 238046 374678 238102
rect 374058 237978 374678 238046
rect 374058 237922 374154 237978
rect 374210 237922 374278 237978
rect 374334 237922 374402 237978
rect 374458 237922 374526 237978
rect 374582 237922 374678 237978
rect 374058 220350 374678 237922
rect 374058 220294 374154 220350
rect 374210 220294 374278 220350
rect 374334 220294 374402 220350
rect 374458 220294 374526 220350
rect 374582 220294 374678 220350
rect 374058 220226 374678 220294
rect 374058 220170 374154 220226
rect 374210 220170 374278 220226
rect 374334 220170 374402 220226
rect 374458 220170 374526 220226
rect 374582 220170 374678 220226
rect 374058 220102 374678 220170
rect 374058 220046 374154 220102
rect 374210 220046 374278 220102
rect 374334 220046 374402 220102
rect 374458 220046 374526 220102
rect 374582 220046 374678 220102
rect 374058 219978 374678 220046
rect 374058 219922 374154 219978
rect 374210 219922 374278 219978
rect 374334 219922 374402 219978
rect 374458 219922 374526 219978
rect 374582 219922 374678 219978
rect 374058 202350 374678 219922
rect 374058 202294 374154 202350
rect 374210 202294 374278 202350
rect 374334 202294 374402 202350
rect 374458 202294 374526 202350
rect 374582 202294 374678 202350
rect 374058 202226 374678 202294
rect 374058 202170 374154 202226
rect 374210 202170 374278 202226
rect 374334 202170 374402 202226
rect 374458 202170 374526 202226
rect 374582 202170 374678 202226
rect 374058 202102 374678 202170
rect 374058 202046 374154 202102
rect 374210 202046 374278 202102
rect 374334 202046 374402 202102
rect 374458 202046 374526 202102
rect 374582 202046 374678 202102
rect 374058 201978 374678 202046
rect 374058 201922 374154 201978
rect 374210 201922 374278 201978
rect 374334 201922 374402 201978
rect 374458 201922 374526 201978
rect 374582 201922 374678 201978
rect 374058 184350 374678 201922
rect 374058 184294 374154 184350
rect 374210 184294 374278 184350
rect 374334 184294 374402 184350
rect 374458 184294 374526 184350
rect 374582 184294 374678 184350
rect 374058 184226 374678 184294
rect 374058 184170 374154 184226
rect 374210 184170 374278 184226
rect 374334 184170 374402 184226
rect 374458 184170 374526 184226
rect 374582 184170 374678 184226
rect 374058 184102 374678 184170
rect 374058 184046 374154 184102
rect 374210 184046 374278 184102
rect 374334 184046 374402 184102
rect 374458 184046 374526 184102
rect 374582 184046 374678 184102
rect 374058 183978 374678 184046
rect 374058 183922 374154 183978
rect 374210 183922 374278 183978
rect 374334 183922 374402 183978
rect 374458 183922 374526 183978
rect 374582 183922 374678 183978
rect 374058 166350 374678 183922
rect 374058 166294 374154 166350
rect 374210 166294 374278 166350
rect 374334 166294 374402 166350
rect 374458 166294 374526 166350
rect 374582 166294 374678 166350
rect 374058 166226 374678 166294
rect 374058 166170 374154 166226
rect 374210 166170 374278 166226
rect 374334 166170 374402 166226
rect 374458 166170 374526 166226
rect 374582 166170 374678 166226
rect 374058 166102 374678 166170
rect 374058 166046 374154 166102
rect 374210 166046 374278 166102
rect 374334 166046 374402 166102
rect 374458 166046 374526 166102
rect 374582 166046 374678 166102
rect 374058 165978 374678 166046
rect 374058 165922 374154 165978
rect 374210 165922 374278 165978
rect 374334 165922 374402 165978
rect 374458 165922 374526 165978
rect 374582 165922 374678 165978
rect 374058 148350 374678 165922
rect 374058 148294 374154 148350
rect 374210 148294 374278 148350
rect 374334 148294 374402 148350
rect 374458 148294 374526 148350
rect 374582 148294 374678 148350
rect 374058 148226 374678 148294
rect 374058 148170 374154 148226
rect 374210 148170 374278 148226
rect 374334 148170 374402 148226
rect 374458 148170 374526 148226
rect 374582 148170 374678 148226
rect 374058 148102 374678 148170
rect 374058 148046 374154 148102
rect 374210 148046 374278 148102
rect 374334 148046 374402 148102
rect 374458 148046 374526 148102
rect 374582 148046 374678 148102
rect 374058 147978 374678 148046
rect 374058 147922 374154 147978
rect 374210 147922 374278 147978
rect 374334 147922 374402 147978
rect 374458 147922 374526 147978
rect 374582 147922 374678 147978
rect 374058 130350 374678 147922
rect 374058 130294 374154 130350
rect 374210 130294 374278 130350
rect 374334 130294 374402 130350
rect 374458 130294 374526 130350
rect 374582 130294 374678 130350
rect 374058 130226 374678 130294
rect 374058 130170 374154 130226
rect 374210 130170 374278 130226
rect 374334 130170 374402 130226
rect 374458 130170 374526 130226
rect 374582 130170 374678 130226
rect 374058 130102 374678 130170
rect 374058 130046 374154 130102
rect 374210 130046 374278 130102
rect 374334 130046 374402 130102
rect 374458 130046 374526 130102
rect 374582 130046 374678 130102
rect 374058 129978 374678 130046
rect 374058 129922 374154 129978
rect 374210 129922 374278 129978
rect 374334 129922 374402 129978
rect 374458 129922 374526 129978
rect 374582 129922 374678 129978
rect 374058 112350 374678 129922
rect 374058 112294 374154 112350
rect 374210 112294 374278 112350
rect 374334 112294 374402 112350
rect 374458 112294 374526 112350
rect 374582 112294 374678 112350
rect 374058 112226 374678 112294
rect 374058 112170 374154 112226
rect 374210 112170 374278 112226
rect 374334 112170 374402 112226
rect 374458 112170 374526 112226
rect 374582 112170 374678 112226
rect 374058 112102 374678 112170
rect 374058 112046 374154 112102
rect 374210 112046 374278 112102
rect 374334 112046 374402 112102
rect 374458 112046 374526 112102
rect 374582 112046 374678 112102
rect 374058 111978 374678 112046
rect 374058 111922 374154 111978
rect 374210 111922 374278 111978
rect 374334 111922 374402 111978
rect 374458 111922 374526 111978
rect 374582 111922 374678 111978
rect 374058 94350 374678 111922
rect 374058 94294 374154 94350
rect 374210 94294 374278 94350
rect 374334 94294 374402 94350
rect 374458 94294 374526 94350
rect 374582 94294 374678 94350
rect 374058 94226 374678 94294
rect 374058 94170 374154 94226
rect 374210 94170 374278 94226
rect 374334 94170 374402 94226
rect 374458 94170 374526 94226
rect 374582 94170 374678 94226
rect 374058 94102 374678 94170
rect 374058 94046 374154 94102
rect 374210 94046 374278 94102
rect 374334 94046 374402 94102
rect 374458 94046 374526 94102
rect 374582 94046 374678 94102
rect 374058 93978 374678 94046
rect 374058 93922 374154 93978
rect 374210 93922 374278 93978
rect 374334 93922 374402 93978
rect 374458 93922 374526 93978
rect 374582 93922 374678 93978
rect 374058 76350 374678 93922
rect 374058 76294 374154 76350
rect 374210 76294 374278 76350
rect 374334 76294 374402 76350
rect 374458 76294 374526 76350
rect 374582 76294 374678 76350
rect 374058 76226 374678 76294
rect 374058 76170 374154 76226
rect 374210 76170 374278 76226
rect 374334 76170 374402 76226
rect 374458 76170 374526 76226
rect 374582 76170 374678 76226
rect 374058 76102 374678 76170
rect 374058 76046 374154 76102
rect 374210 76046 374278 76102
rect 374334 76046 374402 76102
rect 374458 76046 374526 76102
rect 374582 76046 374678 76102
rect 374058 75978 374678 76046
rect 374058 75922 374154 75978
rect 374210 75922 374278 75978
rect 374334 75922 374402 75978
rect 374458 75922 374526 75978
rect 374582 75922 374678 75978
rect 374058 58350 374678 75922
rect 374058 58294 374154 58350
rect 374210 58294 374278 58350
rect 374334 58294 374402 58350
rect 374458 58294 374526 58350
rect 374582 58294 374678 58350
rect 374058 58226 374678 58294
rect 374058 58170 374154 58226
rect 374210 58170 374278 58226
rect 374334 58170 374402 58226
rect 374458 58170 374526 58226
rect 374582 58170 374678 58226
rect 374058 58102 374678 58170
rect 374058 58046 374154 58102
rect 374210 58046 374278 58102
rect 374334 58046 374402 58102
rect 374458 58046 374526 58102
rect 374582 58046 374678 58102
rect 374058 57978 374678 58046
rect 374058 57922 374154 57978
rect 374210 57922 374278 57978
rect 374334 57922 374402 57978
rect 374458 57922 374526 57978
rect 374582 57922 374678 57978
rect 364588 44218 364644 44228
rect 352828 44038 352884 44048
rect 347058 28294 347154 28350
rect 347210 28294 347278 28350
rect 347334 28294 347402 28350
rect 347458 28294 347526 28350
rect 347582 28294 347678 28350
rect 347058 28226 347678 28294
rect 347058 28170 347154 28226
rect 347210 28170 347278 28226
rect 347334 28170 347402 28226
rect 347458 28170 347526 28226
rect 347582 28170 347678 28226
rect 347058 28102 347678 28170
rect 347058 28046 347154 28102
rect 347210 28046 347278 28102
rect 347334 28046 347402 28102
rect 347458 28046 347526 28102
rect 347582 28046 347678 28102
rect 347058 27978 347678 28046
rect 347058 27922 347154 27978
rect 347210 27922 347278 27978
rect 347334 27922 347402 27978
rect 347458 27922 347526 27978
rect 347582 27922 347678 27978
rect 347058 10350 347678 27922
rect 351148 43858 351204 43868
rect 347058 10294 347154 10350
rect 347210 10294 347278 10350
rect 347334 10294 347402 10350
rect 347458 10294 347526 10350
rect 347582 10294 347678 10350
rect 347058 10226 347678 10294
rect 347058 10170 347154 10226
rect 347210 10170 347278 10226
rect 347334 10170 347402 10226
rect 347458 10170 347526 10226
rect 347582 10170 347678 10226
rect 347058 10102 347678 10170
rect 347058 10046 347154 10102
rect 347210 10046 347278 10102
rect 347334 10046 347402 10102
rect 347458 10046 347526 10102
rect 347582 10046 347678 10102
rect 347058 9978 347678 10046
rect 347058 9922 347154 9978
rect 347210 9922 347278 9978
rect 347334 9922 347402 9978
rect 347458 9922 347526 9978
rect 347582 9922 347678 9978
rect 343338 4046 343434 4102
rect 343490 4046 343558 4102
rect 343614 4046 343682 4102
rect 343738 4046 343806 4102
rect 343862 4046 343958 4102
rect 343338 3978 343958 4046
rect 343338 3922 343434 3978
rect 343490 3922 343558 3978
rect 343614 3922 343682 3978
rect 343738 3922 343806 3978
rect 343862 3922 343958 3978
rect 343338 -160 343958 3922
rect 343338 -216 343434 -160
rect 343490 -216 343558 -160
rect 343614 -216 343682 -160
rect 343738 -216 343806 -160
rect 343862 -216 343958 -160
rect 343338 -284 343958 -216
rect 343338 -340 343434 -284
rect 343490 -340 343558 -284
rect 343614 -340 343682 -284
rect 343738 -340 343806 -284
rect 343862 -340 343958 -284
rect 343338 -408 343958 -340
rect 343338 -464 343434 -408
rect 343490 -464 343558 -408
rect 343614 -464 343682 -408
rect 343738 -464 343806 -408
rect 343862 -464 343958 -408
rect 343338 -532 343958 -464
rect 343338 -588 343434 -532
rect 343490 -588 343558 -532
rect 343614 -588 343682 -532
rect 343738 -588 343806 -532
rect 343862 -588 343958 -532
rect 343338 -1644 343958 -588
rect 347058 -1120 347678 9922
rect 347788 24058 347844 24068
rect 347788 4228 347844 24002
rect 347788 4162 347844 4172
rect 351148 4228 351204 43802
rect 351148 4162 351204 4172
rect 352828 4228 352884 43982
rect 362908 42238 362964 42248
rect 359548 20278 359604 20288
rect 359548 20188 359604 20222
rect 359548 20132 359828 20188
rect 352828 4162 352884 4172
rect 359772 4228 359828 20132
rect 359772 4162 359828 4172
rect 362908 4228 362964 42182
rect 362908 4162 362964 4172
rect 364588 4228 364644 44162
rect 374058 40350 374678 57922
rect 377778 598172 378398 598268
rect 377778 598116 377874 598172
rect 377930 598116 377998 598172
rect 378054 598116 378122 598172
rect 378178 598116 378246 598172
rect 378302 598116 378398 598172
rect 377778 598048 378398 598116
rect 377778 597992 377874 598048
rect 377930 597992 377998 598048
rect 378054 597992 378122 598048
rect 378178 597992 378246 598048
rect 378302 597992 378398 598048
rect 377778 597924 378398 597992
rect 377778 597868 377874 597924
rect 377930 597868 377998 597924
rect 378054 597868 378122 597924
rect 378178 597868 378246 597924
rect 378302 597868 378398 597924
rect 377778 597800 378398 597868
rect 377778 597744 377874 597800
rect 377930 597744 377998 597800
rect 378054 597744 378122 597800
rect 378178 597744 378246 597800
rect 378302 597744 378398 597800
rect 377778 586350 378398 597744
rect 377778 586294 377874 586350
rect 377930 586294 377998 586350
rect 378054 586294 378122 586350
rect 378178 586294 378246 586350
rect 378302 586294 378398 586350
rect 377778 586226 378398 586294
rect 377778 586170 377874 586226
rect 377930 586170 377998 586226
rect 378054 586170 378122 586226
rect 378178 586170 378246 586226
rect 378302 586170 378398 586226
rect 377778 586102 378398 586170
rect 377778 586046 377874 586102
rect 377930 586046 377998 586102
rect 378054 586046 378122 586102
rect 378178 586046 378246 586102
rect 378302 586046 378398 586102
rect 377778 585978 378398 586046
rect 377778 585922 377874 585978
rect 377930 585922 377998 585978
rect 378054 585922 378122 585978
rect 378178 585922 378246 585978
rect 378302 585922 378398 585978
rect 377778 568350 378398 585922
rect 377778 568294 377874 568350
rect 377930 568294 377998 568350
rect 378054 568294 378122 568350
rect 378178 568294 378246 568350
rect 378302 568294 378398 568350
rect 377778 568226 378398 568294
rect 377778 568170 377874 568226
rect 377930 568170 377998 568226
rect 378054 568170 378122 568226
rect 378178 568170 378246 568226
rect 378302 568170 378398 568226
rect 377778 568102 378398 568170
rect 377778 568046 377874 568102
rect 377930 568046 377998 568102
rect 378054 568046 378122 568102
rect 378178 568046 378246 568102
rect 378302 568046 378398 568102
rect 377778 567978 378398 568046
rect 377778 567922 377874 567978
rect 377930 567922 377998 567978
rect 378054 567922 378122 567978
rect 378178 567922 378246 567978
rect 378302 567922 378398 567978
rect 377778 550350 378398 567922
rect 377778 550294 377874 550350
rect 377930 550294 377998 550350
rect 378054 550294 378122 550350
rect 378178 550294 378246 550350
rect 378302 550294 378398 550350
rect 377778 550226 378398 550294
rect 377778 550170 377874 550226
rect 377930 550170 377998 550226
rect 378054 550170 378122 550226
rect 378178 550170 378246 550226
rect 378302 550170 378398 550226
rect 377778 550102 378398 550170
rect 377778 550046 377874 550102
rect 377930 550046 377998 550102
rect 378054 550046 378122 550102
rect 378178 550046 378246 550102
rect 378302 550046 378398 550102
rect 377778 549978 378398 550046
rect 377778 549922 377874 549978
rect 377930 549922 377998 549978
rect 378054 549922 378122 549978
rect 378178 549922 378246 549978
rect 378302 549922 378398 549978
rect 377778 532350 378398 549922
rect 377778 532294 377874 532350
rect 377930 532294 377998 532350
rect 378054 532294 378122 532350
rect 378178 532294 378246 532350
rect 378302 532294 378398 532350
rect 377778 532226 378398 532294
rect 377778 532170 377874 532226
rect 377930 532170 377998 532226
rect 378054 532170 378122 532226
rect 378178 532170 378246 532226
rect 378302 532170 378398 532226
rect 377778 532102 378398 532170
rect 377778 532046 377874 532102
rect 377930 532046 377998 532102
rect 378054 532046 378122 532102
rect 378178 532046 378246 532102
rect 378302 532046 378398 532102
rect 377778 531978 378398 532046
rect 377778 531922 377874 531978
rect 377930 531922 377998 531978
rect 378054 531922 378122 531978
rect 378178 531922 378246 531978
rect 378302 531922 378398 531978
rect 377778 514350 378398 531922
rect 377778 514294 377874 514350
rect 377930 514294 377998 514350
rect 378054 514294 378122 514350
rect 378178 514294 378246 514350
rect 378302 514294 378398 514350
rect 377778 514226 378398 514294
rect 377778 514170 377874 514226
rect 377930 514170 377998 514226
rect 378054 514170 378122 514226
rect 378178 514170 378246 514226
rect 378302 514170 378398 514226
rect 377778 514102 378398 514170
rect 377778 514046 377874 514102
rect 377930 514046 377998 514102
rect 378054 514046 378122 514102
rect 378178 514046 378246 514102
rect 378302 514046 378398 514102
rect 377778 513978 378398 514046
rect 377778 513922 377874 513978
rect 377930 513922 377998 513978
rect 378054 513922 378122 513978
rect 378178 513922 378246 513978
rect 378302 513922 378398 513978
rect 377778 496350 378398 513922
rect 377778 496294 377874 496350
rect 377930 496294 377998 496350
rect 378054 496294 378122 496350
rect 378178 496294 378246 496350
rect 378302 496294 378398 496350
rect 377778 496226 378398 496294
rect 377778 496170 377874 496226
rect 377930 496170 377998 496226
rect 378054 496170 378122 496226
rect 378178 496170 378246 496226
rect 378302 496170 378398 496226
rect 377778 496102 378398 496170
rect 377778 496046 377874 496102
rect 377930 496046 377998 496102
rect 378054 496046 378122 496102
rect 378178 496046 378246 496102
rect 378302 496046 378398 496102
rect 377778 495978 378398 496046
rect 377778 495922 377874 495978
rect 377930 495922 377998 495978
rect 378054 495922 378122 495978
rect 378178 495922 378246 495978
rect 378302 495922 378398 495978
rect 377778 478350 378398 495922
rect 377778 478294 377874 478350
rect 377930 478294 377998 478350
rect 378054 478294 378122 478350
rect 378178 478294 378246 478350
rect 378302 478294 378398 478350
rect 377778 478226 378398 478294
rect 377778 478170 377874 478226
rect 377930 478170 377998 478226
rect 378054 478170 378122 478226
rect 378178 478170 378246 478226
rect 378302 478170 378398 478226
rect 377778 478102 378398 478170
rect 377778 478046 377874 478102
rect 377930 478046 377998 478102
rect 378054 478046 378122 478102
rect 378178 478046 378246 478102
rect 378302 478046 378398 478102
rect 377778 477978 378398 478046
rect 377778 477922 377874 477978
rect 377930 477922 377998 477978
rect 378054 477922 378122 477978
rect 378178 477922 378246 477978
rect 378302 477922 378398 477978
rect 377778 460350 378398 477922
rect 377778 460294 377874 460350
rect 377930 460294 377998 460350
rect 378054 460294 378122 460350
rect 378178 460294 378246 460350
rect 378302 460294 378398 460350
rect 377778 460226 378398 460294
rect 377778 460170 377874 460226
rect 377930 460170 377998 460226
rect 378054 460170 378122 460226
rect 378178 460170 378246 460226
rect 378302 460170 378398 460226
rect 377778 460102 378398 460170
rect 377778 460046 377874 460102
rect 377930 460046 377998 460102
rect 378054 460046 378122 460102
rect 378178 460046 378246 460102
rect 378302 460046 378398 460102
rect 377778 459978 378398 460046
rect 377778 459922 377874 459978
rect 377930 459922 377998 459978
rect 378054 459922 378122 459978
rect 378178 459922 378246 459978
rect 378302 459922 378398 459978
rect 377778 442350 378398 459922
rect 377778 442294 377874 442350
rect 377930 442294 377998 442350
rect 378054 442294 378122 442350
rect 378178 442294 378246 442350
rect 378302 442294 378398 442350
rect 377778 442226 378398 442294
rect 377778 442170 377874 442226
rect 377930 442170 377998 442226
rect 378054 442170 378122 442226
rect 378178 442170 378246 442226
rect 378302 442170 378398 442226
rect 377778 442102 378398 442170
rect 377778 442046 377874 442102
rect 377930 442046 377998 442102
rect 378054 442046 378122 442102
rect 378178 442046 378246 442102
rect 378302 442046 378398 442102
rect 377778 441978 378398 442046
rect 377778 441922 377874 441978
rect 377930 441922 377998 441978
rect 378054 441922 378122 441978
rect 378178 441922 378246 441978
rect 378302 441922 378398 441978
rect 377778 424350 378398 441922
rect 377778 424294 377874 424350
rect 377930 424294 377998 424350
rect 378054 424294 378122 424350
rect 378178 424294 378246 424350
rect 378302 424294 378398 424350
rect 377778 424226 378398 424294
rect 377778 424170 377874 424226
rect 377930 424170 377998 424226
rect 378054 424170 378122 424226
rect 378178 424170 378246 424226
rect 378302 424170 378398 424226
rect 377778 424102 378398 424170
rect 377778 424046 377874 424102
rect 377930 424046 377998 424102
rect 378054 424046 378122 424102
rect 378178 424046 378246 424102
rect 378302 424046 378398 424102
rect 377778 423978 378398 424046
rect 377778 423922 377874 423978
rect 377930 423922 377998 423978
rect 378054 423922 378122 423978
rect 378178 423922 378246 423978
rect 378302 423922 378398 423978
rect 377778 406350 378398 423922
rect 377778 406294 377874 406350
rect 377930 406294 377998 406350
rect 378054 406294 378122 406350
rect 378178 406294 378246 406350
rect 378302 406294 378398 406350
rect 377778 406226 378398 406294
rect 377778 406170 377874 406226
rect 377930 406170 377998 406226
rect 378054 406170 378122 406226
rect 378178 406170 378246 406226
rect 378302 406170 378398 406226
rect 377778 406102 378398 406170
rect 377778 406046 377874 406102
rect 377930 406046 377998 406102
rect 378054 406046 378122 406102
rect 378178 406046 378246 406102
rect 378302 406046 378398 406102
rect 377778 405978 378398 406046
rect 377778 405922 377874 405978
rect 377930 405922 377998 405978
rect 378054 405922 378122 405978
rect 378178 405922 378246 405978
rect 378302 405922 378398 405978
rect 377778 388350 378398 405922
rect 377778 388294 377874 388350
rect 377930 388294 377998 388350
rect 378054 388294 378122 388350
rect 378178 388294 378246 388350
rect 378302 388294 378398 388350
rect 377778 388226 378398 388294
rect 377778 388170 377874 388226
rect 377930 388170 377998 388226
rect 378054 388170 378122 388226
rect 378178 388170 378246 388226
rect 378302 388170 378398 388226
rect 377778 388102 378398 388170
rect 377778 388046 377874 388102
rect 377930 388046 377998 388102
rect 378054 388046 378122 388102
rect 378178 388046 378246 388102
rect 378302 388046 378398 388102
rect 377778 387978 378398 388046
rect 377778 387922 377874 387978
rect 377930 387922 377998 387978
rect 378054 387922 378122 387978
rect 378178 387922 378246 387978
rect 378302 387922 378398 387978
rect 377778 370350 378398 387922
rect 377778 370294 377874 370350
rect 377930 370294 377998 370350
rect 378054 370294 378122 370350
rect 378178 370294 378246 370350
rect 378302 370294 378398 370350
rect 377778 370226 378398 370294
rect 377778 370170 377874 370226
rect 377930 370170 377998 370226
rect 378054 370170 378122 370226
rect 378178 370170 378246 370226
rect 378302 370170 378398 370226
rect 377778 370102 378398 370170
rect 377778 370046 377874 370102
rect 377930 370046 377998 370102
rect 378054 370046 378122 370102
rect 378178 370046 378246 370102
rect 378302 370046 378398 370102
rect 377778 369978 378398 370046
rect 377778 369922 377874 369978
rect 377930 369922 377998 369978
rect 378054 369922 378122 369978
rect 378178 369922 378246 369978
rect 378302 369922 378398 369978
rect 377778 352350 378398 369922
rect 377778 352294 377874 352350
rect 377930 352294 377998 352350
rect 378054 352294 378122 352350
rect 378178 352294 378246 352350
rect 378302 352294 378398 352350
rect 377778 352226 378398 352294
rect 377778 352170 377874 352226
rect 377930 352170 377998 352226
rect 378054 352170 378122 352226
rect 378178 352170 378246 352226
rect 378302 352170 378398 352226
rect 377778 352102 378398 352170
rect 377778 352046 377874 352102
rect 377930 352046 377998 352102
rect 378054 352046 378122 352102
rect 378178 352046 378246 352102
rect 378302 352046 378398 352102
rect 377778 351978 378398 352046
rect 377778 351922 377874 351978
rect 377930 351922 377998 351978
rect 378054 351922 378122 351978
rect 378178 351922 378246 351978
rect 378302 351922 378398 351978
rect 377778 334350 378398 351922
rect 377778 334294 377874 334350
rect 377930 334294 377998 334350
rect 378054 334294 378122 334350
rect 378178 334294 378246 334350
rect 378302 334294 378398 334350
rect 377778 334226 378398 334294
rect 377778 334170 377874 334226
rect 377930 334170 377998 334226
rect 378054 334170 378122 334226
rect 378178 334170 378246 334226
rect 378302 334170 378398 334226
rect 377778 334102 378398 334170
rect 377778 334046 377874 334102
rect 377930 334046 377998 334102
rect 378054 334046 378122 334102
rect 378178 334046 378246 334102
rect 378302 334046 378398 334102
rect 377778 333978 378398 334046
rect 377778 333922 377874 333978
rect 377930 333922 377998 333978
rect 378054 333922 378122 333978
rect 378178 333922 378246 333978
rect 378302 333922 378398 333978
rect 377778 316350 378398 333922
rect 377778 316294 377874 316350
rect 377930 316294 377998 316350
rect 378054 316294 378122 316350
rect 378178 316294 378246 316350
rect 378302 316294 378398 316350
rect 377778 316226 378398 316294
rect 377778 316170 377874 316226
rect 377930 316170 377998 316226
rect 378054 316170 378122 316226
rect 378178 316170 378246 316226
rect 378302 316170 378398 316226
rect 377778 316102 378398 316170
rect 377778 316046 377874 316102
rect 377930 316046 377998 316102
rect 378054 316046 378122 316102
rect 378178 316046 378246 316102
rect 378302 316046 378398 316102
rect 377778 315978 378398 316046
rect 377778 315922 377874 315978
rect 377930 315922 377998 315978
rect 378054 315922 378122 315978
rect 378178 315922 378246 315978
rect 378302 315922 378398 315978
rect 377778 298350 378398 315922
rect 377778 298294 377874 298350
rect 377930 298294 377998 298350
rect 378054 298294 378122 298350
rect 378178 298294 378246 298350
rect 378302 298294 378398 298350
rect 377778 298226 378398 298294
rect 377778 298170 377874 298226
rect 377930 298170 377998 298226
rect 378054 298170 378122 298226
rect 378178 298170 378246 298226
rect 378302 298170 378398 298226
rect 377778 298102 378398 298170
rect 377778 298046 377874 298102
rect 377930 298046 377998 298102
rect 378054 298046 378122 298102
rect 378178 298046 378246 298102
rect 378302 298046 378398 298102
rect 377778 297978 378398 298046
rect 377778 297922 377874 297978
rect 377930 297922 377998 297978
rect 378054 297922 378122 297978
rect 378178 297922 378246 297978
rect 378302 297922 378398 297978
rect 377778 280350 378398 297922
rect 377778 280294 377874 280350
rect 377930 280294 377998 280350
rect 378054 280294 378122 280350
rect 378178 280294 378246 280350
rect 378302 280294 378398 280350
rect 377778 280226 378398 280294
rect 377778 280170 377874 280226
rect 377930 280170 377998 280226
rect 378054 280170 378122 280226
rect 378178 280170 378246 280226
rect 378302 280170 378398 280226
rect 377778 280102 378398 280170
rect 377778 280046 377874 280102
rect 377930 280046 377998 280102
rect 378054 280046 378122 280102
rect 378178 280046 378246 280102
rect 378302 280046 378398 280102
rect 377778 279978 378398 280046
rect 377778 279922 377874 279978
rect 377930 279922 377998 279978
rect 378054 279922 378122 279978
rect 378178 279922 378246 279978
rect 378302 279922 378398 279978
rect 377778 262350 378398 279922
rect 377778 262294 377874 262350
rect 377930 262294 377998 262350
rect 378054 262294 378122 262350
rect 378178 262294 378246 262350
rect 378302 262294 378398 262350
rect 377778 262226 378398 262294
rect 377778 262170 377874 262226
rect 377930 262170 377998 262226
rect 378054 262170 378122 262226
rect 378178 262170 378246 262226
rect 378302 262170 378398 262226
rect 377778 262102 378398 262170
rect 377778 262046 377874 262102
rect 377930 262046 377998 262102
rect 378054 262046 378122 262102
rect 378178 262046 378246 262102
rect 378302 262046 378398 262102
rect 377778 261978 378398 262046
rect 377778 261922 377874 261978
rect 377930 261922 377998 261978
rect 378054 261922 378122 261978
rect 378178 261922 378246 261978
rect 378302 261922 378398 261978
rect 377778 244350 378398 261922
rect 377778 244294 377874 244350
rect 377930 244294 377998 244350
rect 378054 244294 378122 244350
rect 378178 244294 378246 244350
rect 378302 244294 378398 244350
rect 377778 244226 378398 244294
rect 377778 244170 377874 244226
rect 377930 244170 377998 244226
rect 378054 244170 378122 244226
rect 378178 244170 378246 244226
rect 378302 244170 378398 244226
rect 377778 244102 378398 244170
rect 377778 244046 377874 244102
rect 377930 244046 377998 244102
rect 378054 244046 378122 244102
rect 378178 244046 378246 244102
rect 378302 244046 378398 244102
rect 377778 243978 378398 244046
rect 377778 243922 377874 243978
rect 377930 243922 377998 243978
rect 378054 243922 378122 243978
rect 378178 243922 378246 243978
rect 378302 243922 378398 243978
rect 377778 226350 378398 243922
rect 377778 226294 377874 226350
rect 377930 226294 377998 226350
rect 378054 226294 378122 226350
rect 378178 226294 378246 226350
rect 378302 226294 378398 226350
rect 377778 226226 378398 226294
rect 377778 226170 377874 226226
rect 377930 226170 377998 226226
rect 378054 226170 378122 226226
rect 378178 226170 378246 226226
rect 378302 226170 378398 226226
rect 377778 226102 378398 226170
rect 377778 226046 377874 226102
rect 377930 226046 377998 226102
rect 378054 226046 378122 226102
rect 378178 226046 378246 226102
rect 378302 226046 378398 226102
rect 377778 225978 378398 226046
rect 377778 225922 377874 225978
rect 377930 225922 377998 225978
rect 378054 225922 378122 225978
rect 378178 225922 378246 225978
rect 378302 225922 378398 225978
rect 377778 208350 378398 225922
rect 377778 208294 377874 208350
rect 377930 208294 377998 208350
rect 378054 208294 378122 208350
rect 378178 208294 378246 208350
rect 378302 208294 378398 208350
rect 377778 208226 378398 208294
rect 377778 208170 377874 208226
rect 377930 208170 377998 208226
rect 378054 208170 378122 208226
rect 378178 208170 378246 208226
rect 378302 208170 378398 208226
rect 377778 208102 378398 208170
rect 377778 208046 377874 208102
rect 377930 208046 377998 208102
rect 378054 208046 378122 208102
rect 378178 208046 378246 208102
rect 378302 208046 378398 208102
rect 377778 207978 378398 208046
rect 377778 207922 377874 207978
rect 377930 207922 377998 207978
rect 378054 207922 378122 207978
rect 378178 207922 378246 207978
rect 378302 207922 378398 207978
rect 377778 190350 378398 207922
rect 377778 190294 377874 190350
rect 377930 190294 377998 190350
rect 378054 190294 378122 190350
rect 378178 190294 378246 190350
rect 378302 190294 378398 190350
rect 377778 190226 378398 190294
rect 377778 190170 377874 190226
rect 377930 190170 377998 190226
rect 378054 190170 378122 190226
rect 378178 190170 378246 190226
rect 378302 190170 378398 190226
rect 377778 190102 378398 190170
rect 377778 190046 377874 190102
rect 377930 190046 377998 190102
rect 378054 190046 378122 190102
rect 378178 190046 378246 190102
rect 378302 190046 378398 190102
rect 377778 189978 378398 190046
rect 377778 189922 377874 189978
rect 377930 189922 377998 189978
rect 378054 189922 378122 189978
rect 378178 189922 378246 189978
rect 378302 189922 378398 189978
rect 377778 172350 378398 189922
rect 377778 172294 377874 172350
rect 377930 172294 377998 172350
rect 378054 172294 378122 172350
rect 378178 172294 378246 172350
rect 378302 172294 378398 172350
rect 377778 172226 378398 172294
rect 377778 172170 377874 172226
rect 377930 172170 377998 172226
rect 378054 172170 378122 172226
rect 378178 172170 378246 172226
rect 378302 172170 378398 172226
rect 377778 172102 378398 172170
rect 377778 172046 377874 172102
rect 377930 172046 377998 172102
rect 378054 172046 378122 172102
rect 378178 172046 378246 172102
rect 378302 172046 378398 172102
rect 377778 171978 378398 172046
rect 377778 171922 377874 171978
rect 377930 171922 377998 171978
rect 378054 171922 378122 171978
rect 378178 171922 378246 171978
rect 378302 171922 378398 171978
rect 377778 154350 378398 171922
rect 377778 154294 377874 154350
rect 377930 154294 377998 154350
rect 378054 154294 378122 154350
rect 378178 154294 378246 154350
rect 378302 154294 378398 154350
rect 377778 154226 378398 154294
rect 377778 154170 377874 154226
rect 377930 154170 377998 154226
rect 378054 154170 378122 154226
rect 378178 154170 378246 154226
rect 378302 154170 378398 154226
rect 377778 154102 378398 154170
rect 377778 154046 377874 154102
rect 377930 154046 377998 154102
rect 378054 154046 378122 154102
rect 378178 154046 378246 154102
rect 378302 154046 378398 154102
rect 377778 153978 378398 154046
rect 377778 153922 377874 153978
rect 377930 153922 377998 153978
rect 378054 153922 378122 153978
rect 378178 153922 378246 153978
rect 378302 153922 378398 153978
rect 377778 136350 378398 153922
rect 377778 136294 377874 136350
rect 377930 136294 377998 136350
rect 378054 136294 378122 136350
rect 378178 136294 378246 136350
rect 378302 136294 378398 136350
rect 377778 136226 378398 136294
rect 377778 136170 377874 136226
rect 377930 136170 377998 136226
rect 378054 136170 378122 136226
rect 378178 136170 378246 136226
rect 378302 136170 378398 136226
rect 377778 136102 378398 136170
rect 377778 136046 377874 136102
rect 377930 136046 377998 136102
rect 378054 136046 378122 136102
rect 378178 136046 378246 136102
rect 378302 136046 378398 136102
rect 377778 135978 378398 136046
rect 377778 135922 377874 135978
rect 377930 135922 377998 135978
rect 378054 135922 378122 135978
rect 378178 135922 378246 135978
rect 378302 135922 378398 135978
rect 377778 118350 378398 135922
rect 377778 118294 377874 118350
rect 377930 118294 377998 118350
rect 378054 118294 378122 118350
rect 378178 118294 378246 118350
rect 378302 118294 378398 118350
rect 377778 118226 378398 118294
rect 377778 118170 377874 118226
rect 377930 118170 377998 118226
rect 378054 118170 378122 118226
rect 378178 118170 378246 118226
rect 378302 118170 378398 118226
rect 377778 118102 378398 118170
rect 377778 118046 377874 118102
rect 377930 118046 377998 118102
rect 378054 118046 378122 118102
rect 378178 118046 378246 118102
rect 378302 118046 378398 118102
rect 377778 117978 378398 118046
rect 377778 117922 377874 117978
rect 377930 117922 377998 117978
rect 378054 117922 378122 117978
rect 378178 117922 378246 117978
rect 378302 117922 378398 117978
rect 377778 100350 378398 117922
rect 377778 100294 377874 100350
rect 377930 100294 377998 100350
rect 378054 100294 378122 100350
rect 378178 100294 378246 100350
rect 378302 100294 378398 100350
rect 377778 100226 378398 100294
rect 377778 100170 377874 100226
rect 377930 100170 377998 100226
rect 378054 100170 378122 100226
rect 378178 100170 378246 100226
rect 378302 100170 378398 100226
rect 377778 100102 378398 100170
rect 377778 100046 377874 100102
rect 377930 100046 377998 100102
rect 378054 100046 378122 100102
rect 378178 100046 378246 100102
rect 378302 100046 378398 100102
rect 377778 99978 378398 100046
rect 377778 99922 377874 99978
rect 377930 99922 377998 99978
rect 378054 99922 378122 99978
rect 378178 99922 378246 99978
rect 378302 99922 378398 99978
rect 377778 82350 378398 99922
rect 377778 82294 377874 82350
rect 377930 82294 377998 82350
rect 378054 82294 378122 82350
rect 378178 82294 378246 82350
rect 378302 82294 378398 82350
rect 377778 82226 378398 82294
rect 377778 82170 377874 82226
rect 377930 82170 377998 82226
rect 378054 82170 378122 82226
rect 378178 82170 378246 82226
rect 378302 82170 378398 82226
rect 377778 82102 378398 82170
rect 377778 82046 377874 82102
rect 377930 82046 377998 82102
rect 378054 82046 378122 82102
rect 378178 82046 378246 82102
rect 378302 82046 378398 82102
rect 377778 81978 378398 82046
rect 377778 81922 377874 81978
rect 377930 81922 377998 81978
rect 378054 81922 378122 81978
rect 378178 81922 378246 81978
rect 378302 81922 378398 81978
rect 377778 64350 378398 81922
rect 404778 597212 405398 598268
rect 404778 597156 404874 597212
rect 404930 597156 404998 597212
rect 405054 597156 405122 597212
rect 405178 597156 405246 597212
rect 405302 597156 405398 597212
rect 404778 597088 405398 597156
rect 404778 597032 404874 597088
rect 404930 597032 404998 597088
rect 405054 597032 405122 597088
rect 405178 597032 405246 597088
rect 405302 597032 405398 597088
rect 404778 596964 405398 597032
rect 404778 596908 404874 596964
rect 404930 596908 404998 596964
rect 405054 596908 405122 596964
rect 405178 596908 405246 596964
rect 405302 596908 405398 596964
rect 404778 596840 405398 596908
rect 404778 596784 404874 596840
rect 404930 596784 404998 596840
rect 405054 596784 405122 596840
rect 405178 596784 405246 596840
rect 405302 596784 405398 596840
rect 404778 580350 405398 596784
rect 404778 580294 404874 580350
rect 404930 580294 404998 580350
rect 405054 580294 405122 580350
rect 405178 580294 405246 580350
rect 405302 580294 405398 580350
rect 404778 580226 405398 580294
rect 404778 580170 404874 580226
rect 404930 580170 404998 580226
rect 405054 580170 405122 580226
rect 405178 580170 405246 580226
rect 405302 580170 405398 580226
rect 404778 580102 405398 580170
rect 404778 580046 404874 580102
rect 404930 580046 404998 580102
rect 405054 580046 405122 580102
rect 405178 580046 405246 580102
rect 405302 580046 405398 580102
rect 404778 579978 405398 580046
rect 404778 579922 404874 579978
rect 404930 579922 404998 579978
rect 405054 579922 405122 579978
rect 405178 579922 405246 579978
rect 405302 579922 405398 579978
rect 404778 562350 405398 579922
rect 404778 562294 404874 562350
rect 404930 562294 404998 562350
rect 405054 562294 405122 562350
rect 405178 562294 405246 562350
rect 405302 562294 405398 562350
rect 404778 562226 405398 562294
rect 404778 562170 404874 562226
rect 404930 562170 404998 562226
rect 405054 562170 405122 562226
rect 405178 562170 405246 562226
rect 405302 562170 405398 562226
rect 404778 562102 405398 562170
rect 404778 562046 404874 562102
rect 404930 562046 404998 562102
rect 405054 562046 405122 562102
rect 405178 562046 405246 562102
rect 405302 562046 405398 562102
rect 404778 561978 405398 562046
rect 404778 561922 404874 561978
rect 404930 561922 404998 561978
rect 405054 561922 405122 561978
rect 405178 561922 405246 561978
rect 405302 561922 405398 561978
rect 404778 544350 405398 561922
rect 404778 544294 404874 544350
rect 404930 544294 404998 544350
rect 405054 544294 405122 544350
rect 405178 544294 405246 544350
rect 405302 544294 405398 544350
rect 404778 544226 405398 544294
rect 404778 544170 404874 544226
rect 404930 544170 404998 544226
rect 405054 544170 405122 544226
rect 405178 544170 405246 544226
rect 405302 544170 405398 544226
rect 404778 544102 405398 544170
rect 404778 544046 404874 544102
rect 404930 544046 404998 544102
rect 405054 544046 405122 544102
rect 405178 544046 405246 544102
rect 405302 544046 405398 544102
rect 404778 543978 405398 544046
rect 404778 543922 404874 543978
rect 404930 543922 404998 543978
rect 405054 543922 405122 543978
rect 405178 543922 405246 543978
rect 405302 543922 405398 543978
rect 404778 526350 405398 543922
rect 404778 526294 404874 526350
rect 404930 526294 404998 526350
rect 405054 526294 405122 526350
rect 405178 526294 405246 526350
rect 405302 526294 405398 526350
rect 404778 526226 405398 526294
rect 404778 526170 404874 526226
rect 404930 526170 404998 526226
rect 405054 526170 405122 526226
rect 405178 526170 405246 526226
rect 405302 526170 405398 526226
rect 404778 526102 405398 526170
rect 404778 526046 404874 526102
rect 404930 526046 404998 526102
rect 405054 526046 405122 526102
rect 405178 526046 405246 526102
rect 405302 526046 405398 526102
rect 404778 525978 405398 526046
rect 404778 525922 404874 525978
rect 404930 525922 404998 525978
rect 405054 525922 405122 525978
rect 405178 525922 405246 525978
rect 405302 525922 405398 525978
rect 404778 508350 405398 525922
rect 404778 508294 404874 508350
rect 404930 508294 404998 508350
rect 405054 508294 405122 508350
rect 405178 508294 405246 508350
rect 405302 508294 405398 508350
rect 404778 508226 405398 508294
rect 404778 508170 404874 508226
rect 404930 508170 404998 508226
rect 405054 508170 405122 508226
rect 405178 508170 405246 508226
rect 405302 508170 405398 508226
rect 404778 508102 405398 508170
rect 404778 508046 404874 508102
rect 404930 508046 404998 508102
rect 405054 508046 405122 508102
rect 405178 508046 405246 508102
rect 405302 508046 405398 508102
rect 404778 507978 405398 508046
rect 404778 507922 404874 507978
rect 404930 507922 404998 507978
rect 405054 507922 405122 507978
rect 405178 507922 405246 507978
rect 405302 507922 405398 507978
rect 404778 490350 405398 507922
rect 404778 490294 404874 490350
rect 404930 490294 404998 490350
rect 405054 490294 405122 490350
rect 405178 490294 405246 490350
rect 405302 490294 405398 490350
rect 404778 490226 405398 490294
rect 404778 490170 404874 490226
rect 404930 490170 404998 490226
rect 405054 490170 405122 490226
rect 405178 490170 405246 490226
rect 405302 490170 405398 490226
rect 404778 490102 405398 490170
rect 404778 490046 404874 490102
rect 404930 490046 404998 490102
rect 405054 490046 405122 490102
rect 405178 490046 405246 490102
rect 405302 490046 405398 490102
rect 404778 489978 405398 490046
rect 404778 489922 404874 489978
rect 404930 489922 404998 489978
rect 405054 489922 405122 489978
rect 405178 489922 405246 489978
rect 405302 489922 405398 489978
rect 404778 472350 405398 489922
rect 404778 472294 404874 472350
rect 404930 472294 404998 472350
rect 405054 472294 405122 472350
rect 405178 472294 405246 472350
rect 405302 472294 405398 472350
rect 404778 472226 405398 472294
rect 404778 472170 404874 472226
rect 404930 472170 404998 472226
rect 405054 472170 405122 472226
rect 405178 472170 405246 472226
rect 405302 472170 405398 472226
rect 404778 472102 405398 472170
rect 404778 472046 404874 472102
rect 404930 472046 404998 472102
rect 405054 472046 405122 472102
rect 405178 472046 405246 472102
rect 405302 472046 405398 472102
rect 404778 471978 405398 472046
rect 404778 471922 404874 471978
rect 404930 471922 404998 471978
rect 405054 471922 405122 471978
rect 405178 471922 405246 471978
rect 405302 471922 405398 471978
rect 404778 454350 405398 471922
rect 404778 454294 404874 454350
rect 404930 454294 404998 454350
rect 405054 454294 405122 454350
rect 405178 454294 405246 454350
rect 405302 454294 405398 454350
rect 404778 454226 405398 454294
rect 404778 454170 404874 454226
rect 404930 454170 404998 454226
rect 405054 454170 405122 454226
rect 405178 454170 405246 454226
rect 405302 454170 405398 454226
rect 404778 454102 405398 454170
rect 404778 454046 404874 454102
rect 404930 454046 404998 454102
rect 405054 454046 405122 454102
rect 405178 454046 405246 454102
rect 405302 454046 405398 454102
rect 404778 453978 405398 454046
rect 404778 453922 404874 453978
rect 404930 453922 404998 453978
rect 405054 453922 405122 453978
rect 405178 453922 405246 453978
rect 405302 453922 405398 453978
rect 404778 436350 405398 453922
rect 404778 436294 404874 436350
rect 404930 436294 404998 436350
rect 405054 436294 405122 436350
rect 405178 436294 405246 436350
rect 405302 436294 405398 436350
rect 404778 436226 405398 436294
rect 404778 436170 404874 436226
rect 404930 436170 404998 436226
rect 405054 436170 405122 436226
rect 405178 436170 405246 436226
rect 405302 436170 405398 436226
rect 404778 436102 405398 436170
rect 404778 436046 404874 436102
rect 404930 436046 404998 436102
rect 405054 436046 405122 436102
rect 405178 436046 405246 436102
rect 405302 436046 405398 436102
rect 404778 435978 405398 436046
rect 404778 435922 404874 435978
rect 404930 435922 404998 435978
rect 405054 435922 405122 435978
rect 405178 435922 405246 435978
rect 405302 435922 405398 435978
rect 404778 418350 405398 435922
rect 404778 418294 404874 418350
rect 404930 418294 404998 418350
rect 405054 418294 405122 418350
rect 405178 418294 405246 418350
rect 405302 418294 405398 418350
rect 404778 418226 405398 418294
rect 404778 418170 404874 418226
rect 404930 418170 404998 418226
rect 405054 418170 405122 418226
rect 405178 418170 405246 418226
rect 405302 418170 405398 418226
rect 404778 418102 405398 418170
rect 404778 418046 404874 418102
rect 404930 418046 404998 418102
rect 405054 418046 405122 418102
rect 405178 418046 405246 418102
rect 405302 418046 405398 418102
rect 404778 417978 405398 418046
rect 404778 417922 404874 417978
rect 404930 417922 404998 417978
rect 405054 417922 405122 417978
rect 405178 417922 405246 417978
rect 405302 417922 405398 417978
rect 404778 400350 405398 417922
rect 404778 400294 404874 400350
rect 404930 400294 404998 400350
rect 405054 400294 405122 400350
rect 405178 400294 405246 400350
rect 405302 400294 405398 400350
rect 404778 400226 405398 400294
rect 404778 400170 404874 400226
rect 404930 400170 404998 400226
rect 405054 400170 405122 400226
rect 405178 400170 405246 400226
rect 405302 400170 405398 400226
rect 404778 400102 405398 400170
rect 404778 400046 404874 400102
rect 404930 400046 404998 400102
rect 405054 400046 405122 400102
rect 405178 400046 405246 400102
rect 405302 400046 405398 400102
rect 404778 399978 405398 400046
rect 404778 399922 404874 399978
rect 404930 399922 404998 399978
rect 405054 399922 405122 399978
rect 405178 399922 405246 399978
rect 405302 399922 405398 399978
rect 404778 382350 405398 399922
rect 404778 382294 404874 382350
rect 404930 382294 404998 382350
rect 405054 382294 405122 382350
rect 405178 382294 405246 382350
rect 405302 382294 405398 382350
rect 404778 382226 405398 382294
rect 404778 382170 404874 382226
rect 404930 382170 404998 382226
rect 405054 382170 405122 382226
rect 405178 382170 405246 382226
rect 405302 382170 405398 382226
rect 404778 382102 405398 382170
rect 404778 382046 404874 382102
rect 404930 382046 404998 382102
rect 405054 382046 405122 382102
rect 405178 382046 405246 382102
rect 405302 382046 405398 382102
rect 404778 381978 405398 382046
rect 404778 381922 404874 381978
rect 404930 381922 404998 381978
rect 405054 381922 405122 381978
rect 405178 381922 405246 381978
rect 405302 381922 405398 381978
rect 404778 364350 405398 381922
rect 404778 364294 404874 364350
rect 404930 364294 404998 364350
rect 405054 364294 405122 364350
rect 405178 364294 405246 364350
rect 405302 364294 405398 364350
rect 404778 364226 405398 364294
rect 404778 364170 404874 364226
rect 404930 364170 404998 364226
rect 405054 364170 405122 364226
rect 405178 364170 405246 364226
rect 405302 364170 405398 364226
rect 404778 364102 405398 364170
rect 404778 364046 404874 364102
rect 404930 364046 404998 364102
rect 405054 364046 405122 364102
rect 405178 364046 405246 364102
rect 405302 364046 405398 364102
rect 404778 363978 405398 364046
rect 404778 363922 404874 363978
rect 404930 363922 404998 363978
rect 405054 363922 405122 363978
rect 405178 363922 405246 363978
rect 405302 363922 405398 363978
rect 404778 346350 405398 363922
rect 404778 346294 404874 346350
rect 404930 346294 404998 346350
rect 405054 346294 405122 346350
rect 405178 346294 405246 346350
rect 405302 346294 405398 346350
rect 404778 346226 405398 346294
rect 404778 346170 404874 346226
rect 404930 346170 404998 346226
rect 405054 346170 405122 346226
rect 405178 346170 405246 346226
rect 405302 346170 405398 346226
rect 404778 346102 405398 346170
rect 404778 346046 404874 346102
rect 404930 346046 404998 346102
rect 405054 346046 405122 346102
rect 405178 346046 405246 346102
rect 405302 346046 405398 346102
rect 404778 345978 405398 346046
rect 404778 345922 404874 345978
rect 404930 345922 404998 345978
rect 405054 345922 405122 345978
rect 405178 345922 405246 345978
rect 405302 345922 405398 345978
rect 404778 328350 405398 345922
rect 404778 328294 404874 328350
rect 404930 328294 404998 328350
rect 405054 328294 405122 328350
rect 405178 328294 405246 328350
rect 405302 328294 405398 328350
rect 404778 328226 405398 328294
rect 404778 328170 404874 328226
rect 404930 328170 404998 328226
rect 405054 328170 405122 328226
rect 405178 328170 405246 328226
rect 405302 328170 405398 328226
rect 404778 328102 405398 328170
rect 404778 328046 404874 328102
rect 404930 328046 404998 328102
rect 405054 328046 405122 328102
rect 405178 328046 405246 328102
rect 405302 328046 405398 328102
rect 404778 327978 405398 328046
rect 404778 327922 404874 327978
rect 404930 327922 404998 327978
rect 405054 327922 405122 327978
rect 405178 327922 405246 327978
rect 405302 327922 405398 327978
rect 404778 310350 405398 327922
rect 404778 310294 404874 310350
rect 404930 310294 404998 310350
rect 405054 310294 405122 310350
rect 405178 310294 405246 310350
rect 405302 310294 405398 310350
rect 404778 310226 405398 310294
rect 404778 310170 404874 310226
rect 404930 310170 404998 310226
rect 405054 310170 405122 310226
rect 405178 310170 405246 310226
rect 405302 310170 405398 310226
rect 404778 310102 405398 310170
rect 404778 310046 404874 310102
rect 404930 310046 404998 310102
rect 405054 310046 405122 310102
rect 405178 310046 405246 310102
rect 405302 310046 405398 310102
rect 404778 309978 405398 310046
rect 404778 309922 404874 309978
rect 404930 309922 404998 309978
rect 405054 309922 405122 309978
rect 405178 309922 405246 309978
rect 405302 309922 405398 309978
rect 404778 292350 405398 309922
rect 404778 292294 404874 292350
rect 404930 292294 404998 292350
rect 405054 292294 405122 292350
rect 405178 292294 405246 292350
rect 405302 292294 405398 292350
rect 404778 292226 405398 292294
rect 404778 292170 404874 292226
rect 404930 292170 404998 292226
rect 405054 292170 405122 292226
rect 405178 292170 405246 292226
rect 405302 292170 405398 292226
rect 404778 292102 405398 292170
rect 404778 292046 404874 292102
rect 404930 292046 404998 292102
rect 405054 292046 405122 292102
rect 405178 292046 405246 292102
rect 405302 292046 405398 292102
rect 404778 291978 405398 292046
rect 404778 291922 404874 291978
rect 404930 291922 404998 291978
rect 405054 291922 405122 291978
rect 405178 291922 405246 291978
rect 405302 291922 405398 291978
rect 404778 274350 405398 291922
rect 404778 274294 404874 274350
rect 404930 274294 404998 274350
rect 405054 274294 405122 274350
rect 405178 274294 405246 274350
rect 405302 274294 405398 274350
rect 404778 274226 405398 274294
rect 404778 274170 404874 274226
rect 404930 274170 404998 274226
rect 405054 274170 405122 274226
rect 405178 274170 405246 274226
rect 405302 274170 405398 274226
rect 404778 274102 405398 274170
rect 404778 274046 404874 274102
rect 404930 274046 404998 274102
rect 405054 274046 405122 274102
rect 405178 274046 405246 274102
rect 405302 274046 405398 274102
rect 404778 273978 405398 274046
rect 404778 273922 404874 273978
rect 404930 273922 404998 273978
rect 405054 273922 405122 273978
rect 405178 273922 405246 273978
rect 405302 273922 405398 273978
rect 404778 256350 405398 273922
rect 404778 256294 404874 256350
rect 404930 256294 404998 256350
rect 405054 256294 405122 256350
rect 405178 256294 405246 256350
rect 405302 256294 405398 256350
rect 404778 256226 405398 256294
rect 404778 256170 404874 256226
rect 404930 256170 404998 256226
rect 405054 256170 405122 256226
rect 405178 256170 405246 256226
rect 405302 256170 405398 256226
rect 404778 256102 405398 256170
rect 404778 256046 404874 256102
rect 404930 256046 404998 256102
rect 405054 256046 405122 256102
rect 405178 256046 405246 256102
rect 405302 256046 405398 256102
rect 404778 255978 405398 256046
rect 404778 255922 404874 255978
rect 404930 255922 404998 255978
rect 405054 255922 405122 255978
rect 405178 255922 405246 255978
rect 405302 255922 405398 255978
rect 404778 238350 405398 255922
rect 404778 238294 404874 238350
rect 404930 238294 404998 238350
rect 405054 238294 405122 238350
rect 405178 238294 405246 238350
rect 405302 238294 405398 238350
rect 404778 238226 405398 238294
rect 404778 238170 404874 238226
rect 404930 238170 404998 238226
rect 405054 238170 405122 238226
rect 405178 238170 405246 238226
rect 405302 238170 405398 238226
rect 404778 238102 405398 238170
rect 404778 238046 404874 238102
rect 404930 238046 404998 238102
rect 405054 238046 405122 238102
rect 405178 238046 405246 238102
rect 405302 238046 405398 238102
rect 404778 237978 405398 238046
rect 404778 237922 404874 237978
rect 404930 237922 404998 237978
rect 405054 237922 405122 237978
rect 405178 237922 405246 237978
rect 405302 237922 405398 237978
rect 404778 220350 405398 237922
rect 404778 220294 404874 220350
rect 404930 220294 404998 220350
rect 405054 220294 405122 220350
rect 405178 220294 405246 220350
rect 405302 220294 405398 220350
rect 404778 220226 405398 220294
rect 404778 220170 404874 220226
rect 404930 220170 404998 220226
rect 405054 220170 405122 220226
rect 405178 220170 405246 220226
rect 405302 220170 405398 220226
rect 404778 220102 405398 220170
rect 404778 220046 404874 220102
rect 404930 220046 404998 220102
rect 405054 220046 405122 220102
rect 405178 220046 405246 220102
rect 405302 220046 405398 220102
rect 404778 219978 405398 220046
rect 404778 219922 404874 219978
rect 404930 219922 404998 219978
rect 405054 219922 405122 219978
rect 405178 219922 405246 219978
rect 405302 219922 405398 219978
rect 404778 202350 405398 219922
rect 404778 202294 404874 202350
rect 404930 202294 404998 202350
rect 405054 202294 405122 202350
rect 405178 202294 405246 202350
rect 405302 202294 405398 202350
rect 404778 202226 405398 202294
rect 404778 202170 404874 202226
rect 404930 202170 404998 202226
rect 405054 202170 405122 202226
rect 405178 202170 405246 202226
rect 405302 202170 405398 202226
rect 404778 202102 405398 202170
rect 404778 202046 404874 202102
rect 404930 202046 404998 202102
rect 405054 202046 405122 202102
rect 405178 202046 405246 202102
rect 405302 202046 405398 202102
rect 404778 201978 405398 202046
rect 404778 201922 404874 201978
rect 404930 201922 404998 201978
rect 405054 201922 405122 201978
rect 405178 201922 405246 201978
rect 405302 201922 405398 201978
rect 404778 184350 405398 201922
rect 404778 184294 404874 184350
rect 404930 184294 404998 184350
rect 405054 184294 405122 184350
rect 405178 184294 405246 184350
rect 405302 184294 405398 184350
rect 404778 184226 405398 184294
rect 404778 184170 404874 184226
rect 404930 184170 404998 184226
rect 405054 184170 405122 184226
rect 405178 184170 405246 184226
rect 405302 184170 405398 184226
rect 404778 184102 405398 184170
rect 404778 184046 404874 184102
rect 404930 184046 404998 184102
rect 405054 184046 405122 184102
rect 405178 184046 405246 184102
rect 405302 184046 405398 184102
rect 404778 183978 405398 184046
rect 404778 183922 404874 183978
rect 404930 183922 404998 183978
rect 405054 183922 405122 183978
rect 405178 183922 405246 183978
rect 405302 183922 405398 183978
rect 404778 166350 405398 183922
rect 404778 166294 404874 166350
rect 404930 166294 404998 166350
rect 405054 166294 405122 166350
rect 405178 166294 405246 166350
rect 405302 166294 405398 166350
rect 404778 166226 405398 166294
rect 404778 166170 404874 166226
rect 404930 166170 404998 166226
rect 405054 166170 405122 166226
rect 405178 166170 405246 166226
rect 405302 166170 405398 166226
rect 404778 166102 405398 166170
rect 404778 166046 404874 166102
rect 404930 166046 404998 166102
rect 405054 166046 405122 166102
rect 405178 166046 405246 166102
rect 405302 166046 405398 166102
rect 404778 165978 405398 166046
rect 404778 165922 404874 165978
rect 404930 165922 404998 165978
rect 405054 165922 405122 165978
rect 405178 165922 405246 165978
rect 405302 165922 405398 165978
rect 404778 148350 405398 165922
rect 404778 148294 404874 148350
rect 404930 148294 404998 148350
rect 405054 148294 405122 148350
rect 405178 148294 405246 148350
rect 405302 148294 405398 148350
rect 404778 148226 405398 148294
rect 404778 148170 404874 148226
rect 404930 148170 404998 148226
rect 405054 148170 405122 148226
rect 405178 148170 405246 148226
rect 405302 148170 405398 148226
rect 404778 148102 405398 148170
rect 404778 148046 404874 148102
rect 404930 148046 404998 148102
rect 405054 148046 405122 148102
rect 405178 148046 405246 148102
rect 405302 148046 405398 148102
rect 404778 147978 405398 148046
rect 404778 147922 404874 147978
rect 404930 147922 404998 147978
rect 405054 147922 405122 147978
rect 405178 147922 405246 147978
rect 405302 147922 405398 147978
rect 404778 130350 405398 147922
rect 404778 130294 404874 130350
rect 404930 130294 404998 130350
rect 405054 130294 405122 130350
rect 405178 130294 405246 130350
rect 405302 130294 405398 130350
rect 404778 130226 405398 130294
rect 404778 130170 404874 130226
rect 404930 130170 404998 130226
rect 405054 130170 405122 130226
rect 405178 130170 405246 130226
rect 405302 130170 405398 130226
rect 404778 130102 405398 130170
rect 404778 130046 404874 130102
rect 404930 130046 404998 130102
rect 405054 130046 405122 130102
rect 405178 130046 405246 130102
rect 405302 130046 405398 130102
rect 404778 129978 405398 130046
rect 404778 129922 404874 129978
rect 404930 129922 404998 129978
rect 405054 129922 405122 129978
rect 405178 129922 405246 129978
rect 405302 129922 405398 129978
rect 404778 112350 405398 129922
rect 404778 112294 404874 112350
rect 404930 112294 404998 112350
rect 405054 112294 405122 112350
rect 405178 112294 405246 112350
rect 405302 112294 405398 112350
rect 404778 112226 405398 112294
rect 404778 112170 404874 112226
rect 404930 112170 404998 112226
rect 405054 112170 405122 112226
rect 405178 112170 405246 112226
rect 405302 112170 405398 112226
rect 404778 112102 405398 112170
rect 404778 112046 404874 112102
rect 404930 112046 404998 112102
rect 405054 112046 405122 112102
rect 405178 112046 405246 112102
rect 405302 112046 405398 112102
rect 404778 111978 405398 112046
rect 404778 111922 404874 111978
rect 404930 111922 404998 111978
rect 405054 111922 405122 111978
rect 405178 111922 405246 111978
rect 405302 111922 405398 111978
rect 404778 94350 405398 111922
rect 404778 94294 404874 94350
rect 404930 94294 404998 94350
rect 405054 94294 405122 94350
rect 405178 94294 405246 94350
rect 405302 94294 405398 94350
rect 404778 94226 405398 94294
rect 404778 94170 404874 94226
rect 404930 94170 404998 94226
rect 405054 94170 405122 94226
rect 405178 94170 405246 94226
rect 405302 94170 405398 94226
rect 404778 94102 405398 94170
rect 404778 94046 404874 94102
rect 404930 94046 404998 94102
rect 405054 94046 405122 94102
rect 405178 94046 405246 94102
rect 405302 94046 405398 94102
rect 404778 93978 405398 94046
rect 404778 93922 404874 93978
rect 404930 93922 404998 93978
rect 405054 93922 405122 93978
rect 405178 93922 405246 93978
rect 405302 93922 405398 93978
rect 404778 76350 405398 93922
rect 404778 76294 404874 76350
rect 404930 76294 404998 76350
rect 405054 76294 405122 76350
rect 405178 76294 405246 76350
rect 405302 76294 405398 76350
rect 404778 76226 405398 76294
rect 404778 76170 404874 76226
rect 404930 76170 404998 76226
rect 405054 76170 405122 76226
rect 405178 76170 405246 76226
rect 405302 76170 405398 76226
rect 404778 76102 405398 76170
rect 404778 76046 404874 76102
rect 404930 76046 404998 76102
rect 405054 76046 405122 76102
rect 405178 76046 405246 76102
rect 405302 76046 405398 76102
rect 404778 75978 405398 76046
rect 404778 75922 404874 75978
rect 404930 75922 404998 75978
rect 405054 75922 405122 75978
rect 405178 75922 405246 75978
rect 405302 75922 405398 75978
rect 377778 64294 377874 64350
rect 377930 64294 377998 64350
rect 378054 64294 378122 64350
rect 378178 64294 378246 64350
rect 378302 64294 378398 64350
rect 377778 64226 378398 64294
rect 377778 64170 377874 64226
rect 377930 64170 377998 64226
rect 378054 64170 378122 64226
rect 378178 64170 378246 64226
rect 378302 64170 378398 64226
rect 377778 64102 378398 64170
rect 377778 64046 377874 64102
rect 377930 64046 377998 64102
rect 378054 64046 378122 64102
rect 378178 64046 378246 64102
rect 378302 64046 378398 64102
rect 377778 63978 378398 64046
rect 377778 63922 377874 63978
rect 377930 63922 377998 63978
rect 378054 63922 378122 63978
rect 378178 63922 378246 63978
rect 378302 63922 378398 63978
rect 374058 40294 374154 40350
rect 374210 40294 374278 40350
rect 374334 40294 374402 40350
rect 374458 40294 374526 40350
rect 374582 40294 374678 40350
rect 374058 40226 374678 40294
rect 374058 40170 374154 40226
rect 374210 40170 374278 40226
rect 374334 40170 374402 40226
rect 374458 40170 374526 40226
rect 374582 40170 374678 40226
rect 374058 40102 374678 40170
rect 374058 40046 374154 40102
rect 374210 40046 374278 40102
rect 374334 40046 374402 40102
rect 374458 40046 374526 40102
rect 374582 40046 374678 40102
rect 374058 39978 374678 40046
rect 374058 39922 374154 39978
rect 374210 39922 374278 39978
rect 374334 39922 374402 39978
rect 374458 39922 374526 39978
rect 374582 39922 374678 39978
rect 364588 4162 364644 4172
rect 371308 25678 371364 25688
rect 371308 4228 371364 25622
rect 371308 4162 371364 4172
rect 374058 22350 374678 39922
rect 376348 55918 376404 55928
rect 374058 22294 374154 22350
rect 374210 22294 374278 22350
rect 374334 22294 374402 22350
rect 374458 22294 374526 22350
rect 374582 22294 374678 22350
rect 374058 22226 374678 22294
rect 374058 22170 374154 22226
rect 374210 22170 374278 22226
rect 374334 22170 374402 22226
rect 374458 22170 374526 22226
rect 374582 22170 374678 22226
rect 374058 22102 374678 22170
rect 374058 22046 374154 22102
rect 374210 22046 374278 22102
rect 374334 22046 374402 22102
rect 374458 22046 374526 22102
rect 374582 22046 374678 22102
rect 374058 21978 374678 22046
rect 374058 21922 374154 21978
rect 374210 21922 374278 21978
rect 374334 21922 374402 21978
rect 374458 21922 374526 21978
rect 374582 21922 374678 21978
rect 374058 4350 374678 21922
rect 374780 37198 374836 37208
rect 374780 20188 374836 37142
rect 374780 20132 375060 20188
rect 374058 4294 374154 4350
rect 374210 4294 374278 4350
rect 374334 4294 374402 4350
rect 374458 4294 374526 4350
rect 374582 4294 374678 4350
rect 374058 4226 374678 4294
rect 374058 4170 374154 4226
rect 374210 4170 374278 4226
rect 374334 4170 374402 4226
rect 374458 4170 374526 4226
rect 374582 4170 374678 4226
rect 347058 -1176 347154 -1120
rect 347210 -1176 347278 -1120
rect 347334 -1176 347402 -1120
rect 347458 -1176 347526 -1120
rect 347582 -1176 347678 -1120
rect 347058 -1244 347678 -1176
rect 347058 -1300 347154 -1244
rect 347210 -1300 347278 -1244
rect 347334 -1300 347402 -1244
rect 347458 -1300 347526 -1244
rect 347582 -1300 347678 -1244
rect 347058 -1368 347678 -1300
rect 347058 -1424 347154 -1368
rect 347210 -1424 347278 -1368
rect 347334 -1424 347402 -1368
rect 347458 -1424 347526 -1368
rect 347582 -1424 347678 -1368
rect 347058 -1492 347678 -1424
rect 347058 -1548 347154 -1492
rect 347210 -1548 347278 -1492
rect 347334 -1548 347402 -1492
rect 347458 -1548 347526 -1492
rect 347582 -1548 347678 -1492
rect 347058 -1644 347678 -1548
rect 374058 4102 374678 4170
rect 375004 4228 375060 20132
rect 375004 4162 375060 4172
rect 376348 4228 376404 55862
rect 376348 4162 376404 4172
rect 377778 46350 378398 63922
rect 377778 46294 377874 46350
rect 377930 46294 377998 46350
rect 378054 46294 378122 46350
rect 378178 46294 378246 46350
rect 378302 46294 378398 46350
rect 377778 46226 378398 46294
rect 377778 46170 377874 46226
rect 377930 46170 377998 46226
rect 378054 46170 378122 46226
rect 378178 46170 378246 46226
rect 378302 46170 378398 46226
rect 377778 46102 378398 46170
rect 377778 46046 377874 46102
rect 377930 46046 377998 46102
rect 378054 46046 378122 46102
rect 378178 46046 378246 46102
rect 378302 46046 378398 46102
rect 377778 45978 378398 46046
rect 377778 45922 377874 45978
rect 377930 45922 377998 45978
rect 378054 45922 378122 45978
rect 378178 45922 378246 45978
rect 378302 45922 378398 45978
rect 377778 28350 378398 45922
rect 383068 72658 383124 72668
rect 377778 28294 377874 28350
rect 377930 28294 377998 28350
rect 378054 28294 378122 28350
rect 378178 28294 378246 28350
rect 378302 28294 378398 28350
rect 377778 28226 378398 28294
rect 377778 28170 377874 28226
rect 377930 28170 377998 28226
rect 378054 28170 378122 28226
rect 378178 28170 378246 28226
rect 378302 28170 378398 28226
rect 377778 28102 378398 28170
rect 377778 28046 377874 28102
rect 377930 28046 377998 28102
rect 378054 28046 378122 28102
rect 378178 28046 378246 28102
rect 378302 28046 378398 28102
rect 377778 27978 378398 28046
rect 377778 27922 377874 27978
rect 377930 27922 377998 27978
rect 378054 27922 378122 27978
rect 378178 27922 378246 27978
rect 378302 27922 378398 27978
rect 377778 10350 378398 27922
rect 377778 10294 377874 10350
rect 377930 10294 377998 10350
rect 378054 10294 378122 10350
rect 378178 10294 378246 10350
rect 378302 10294 378398 10350
rect 377778 10226 378398 10294
rect 377778 10170 377874 10226
rect 377930 10170 377998 10226
rect 378054 10170 378122 10226
rect 378178 10170 378246 10226
rect 378302 10170 378398 10226
rect 377778 10102 378398 10170
rect 377778 10046 377874 10102
rect 377930 10046 377998 10102
rect 378054 10046 378122 10102
rect 378178 10046 378246 10102
rect 378302 10046 378398 10102
rect 377778 9978 378398 10046
rect 377778 9922 377874 9978
rect 377930 9922 377998 9978
rect 378054 9922 378122 9978
rect 378178 9922 378246 9978
rect 378302 9922 378398 9978
rect 374058 4046 374154 4102
rect 374210 4046 374278 4102
rect 374334 4046 374402 4102
rect 374458 4046 374526 4102
rect 374582 4046 374678 4102
rect 374058 3978 374678 4046
rect 374058 3922 374154 3978
rect 374210 3922 374278 3978
rect 374334 3922 374402 3978
rect 374458 3922 374526 3978
rect 374582 3922 374678 3978
rect 374058 -160 374678 3922
rect 374058 -216 374154 -160
rect 374210 -216 374278 -160
rect 374334 -216 374402 -160
rect 374458 -216 374526 -160
rect 374582 -216 374678 -160
rect 374058 -284 374678 -216
rect 374058 -340 374154 -284
rect 374210 -340 374278 -284
rect 374334 -340 374402 -284
rect 374458 -340 374526 -284
rect 374582 -340 374678 -284
rect 374058 -408 374678 -340
rect 374058 -464 374154 -408
rect 374210 -464 374278 -408
rect 374334 -464 374402 -408
rect 374458 -464 374526 -408
rect 374582 -464 374678 -408
rect 374058 -532 374678 -464
rect 374058 -588 374154 -532
rect 374210 -588 374278 -532
rect 374334 -588 374402 -532
rect 374458 -588 374526 -532
rect 374582 -588 374678 -532
rect 374058 -1644 374678 -588
rect 377778 -1120 378398 9922
rect 379708 34138 379764 34148
rect 379708 4228 379764 34082
rect 379708 4162 379764 4172
rect 383068 4228 383124 72602
rect 396508 60958 396564 60968
rect 383068 4162 383124 4172
rect 386428 37018 386484 37028
rect 386428 4228 386484 36962
rect 388108 23878 388164 23888
rect 388108 20188 388164 23822
rect 391468 23698 391524 23708
rect 388108 20132 388388 20188
rect 386428 4162 386484 4172
rect 388332 4228 388388 20132
rect 388332 4162 388388 4172
rect 391468 4228 391524 23642
rect 391468 4162 391524 4172
rect 393148 12358 393204 12368
rect 393148 4228 393204 12302
rect 393148 4162 393204 4172
rect 394828 12178 394884 12188
rect 394828 4228 394884 12122
rect 394828 4162 394884 4172
rect 396508 4228 396564 60902
rect 404778 58350 405398 75922
rect 408498 598172 409118 598268
rect 408498 598116 408594 598172
rect 408650 598116 408718 598172
rect 408774 598116 408842 598172
rect 408898 598116 408966 598172
rect 409022 598116 409118 598172
rect 408498 598048 409118 598116
rect 408498 597992 408594 598048
rect 408650 597992 408718 598048
rect 408774 597992 408842 598048
rect 408898 597992 408966 598048
rect 409022 597992 409118 598048
rect 408498 597924 409118 597992
rect 408498 597868 408594 597924
rect 408650 597868 408718 597924
rect 408774 597868 408842 597924
rect 408898 597868 408966 597924
rect 409022 597868 409118 597924
rect 408498 597800 409118 597868
rect 408498 597744 408594 597800
rect 408650 597744 408718 597800
rect 408774 597744 408842 597800
rect 408898 597744 408966 597800
rect 409022 597744 409118 597800
rect 408498 586350 409118 597744
rect 408498 586294 408594 586350
rect 408650 586294 408718 586350
rect 408774 586294 408842 586350
rect 408898 586294 408966 586350
rect 409022 586294 409118 586350
rect 408498 586226 409118 586294
rect 408498 586170 408594 586226
rect 408650 586170 408718 586226
rect 408774 586170 408842 586226
rect 408898 586170 408966 586226
rect 409022 586170 409118 586226
rect 408498 586102 409118 586170
rect 408498 586046 408594 586102
rect 408650 586046 408718 586102
rect 408774 586046 408842 586102
rect 408898 586046 408966 586102
rect 409022 586046 409118 586102
rect 408498 585978 409118 586046
rect 408498 585922 408594 585978
rect 408650 585922 408718 585978
rect 408774 585922 408842 585978
rect 408898 585922 408966 585978
rect 409022 585922 409118 585978
rect 408498 568350 409118 585922
rect 408498 568294 408594 568350
rect 408650 568294 408718 568350
rect 408774 568294 408842 568350
rect 408898 568294 408966 568350
rect 409022 568294 409118 568350
rect 408498 568226 409118 568294
rect 408498 568170 408594 568226
rect 408650 568170 408718 568226
rect 408774 568170 408842 568226
rect 408898 568170 408966 568226
rect 409022 568170 409118 568226
rect 408498 568102 409118 568170
rect 408498 568046 408594 568102
rect 408650 568046 408718 568102
rect 408774 568046 408842 568102
rect 408898 568046 408966 568102
rect 409022 568046 409118 568102
rect 408498 567978 409118 568046
rect 408498 567922 408594 567978
rect 408650 567922 408718 567978
rect 408774 567922 408842 567978
rect 408898 567922 408966 567978
rect 409022 567922 409118 567978
rect 408498 550350 409118 567922
rect 408498 550294 408594 550350
rect 408650 550294 408718 550350
rect 408774 550294 408842 550350
rect 408898 550294 408966 550350
rect 409022 550294 409118 550350
rect 408498 550226 409118 550294
rect 408498 550170 408594 550226
rect 408650 550170 408718 550226
rect 408774 550170 408842 550226
rect 408898 550170 408966 550226
rect 409022 550170 409118 550226
rect 408498 550102 409118 550170
rect 408498 550046 408594 550102
rect 408650 550046 408718 550102
rect 408774 550046 408842 550102
rect 408898 550046 408966 550102
rect 409022 550046 409118 550102
rect 408498 549978 409118 550046
rect 408498 549922 408594 549978
rect 408650 549922 408718 549978
rect 408774 549922 408842 549978
rect 408898 549922 408966 549978
rect 409022 549922 409118 549978
rect 408498 532350 409118 549922
rect 408498 532294 408594 532350
rect 408650 532294 408718 532350
rect 408774 532294 408842 532350
rect 408898 532294 408966 532350
rect 409022 532294 409118 532350
rect 408498 532226 409118 532294
rect 408498 532170 408594 532226
rect 408650 532170 408718 532226
rect 408774 532170 408842 532226
rect 408898 532170 408966 532226
rect 409022 532170 409118 532226
rect 408498 532102 409118 532170
rect 408498 532046 408594 532102
rect 408650 532046 408718 532102
rect 408774 532046 408842 532102
rect 408898 532046 408966 532102
rect 409022 532046 409118 532102
rect 408498 531978 409118 532046
rect 408498 531922 408594 531978
rect 408650 531922 408718 531978
rect 408774 531922 408842 531978
rect 408898 531922 408966 531978
rect 409022 531922 409118 531978
rect 408498 514350 409118 531922
rect 408498 514294 408594 514350
rect 408650 514294 408718 514350
rect 408774 514294 408842 514350
rect 408898 514294 408966 514350
rect 409022 514294 409118 514350
rect 408498 514226 409118 514294
rect 408498 514170 408594 514226
rect 408650 514170 408718 514226
rect 408774 514170 408842 514226
rect 408898 514170 408966 514226
rect 409022 514170 409118 514226
rect 408498 514102 409118 514170
rect 408498 514046 408594 514102
rect 408650 514046 408718 514102
rect 408774 514046 408842 514102
rect 408898 514046 408966 514102
rect 409022 514046 409118 514102
rect 408498 513978 409118 514046
rect 408498 513922 408594 513978
rect 408650 513922 408718 513978
rect 408774 513922 408842 513978
rect 408898 513922 408966 513978
rect 409022 513922 409118 513978
rect 408498 496350 409118 513922
rect 408498 496294 408594 496350
rect 408650 496294 408718 496350
rect 408774 496294 408842 496350
rect 408898 496294 408966 496350
rect 409022 496294 409118 496350
rect 408498 496226 409118 496294
rect 408498 496170 408594 496226
rect 408650 496170 408718 496226
rect 408774 496170 408842 496226
rect 408898 496170 408966 496226
rect 409022 496170 409118 496226
rect 408498 496102 409118 496170
rect 408498 496046 408594 496102
rect 408650 496046 408718 496102
rect 408774 496046 408842 496102
rect 408898 496046 408966 496102
rect 409022 496046 409118 496102
rect 408498 495978 409118 496046
rect 408498 495922 408594 495978
rect 408650 495922 408718 495978
rect 408774 495922 408842 495978
rect 408898 495922 408966 495978
rect 409022 495922 409118 495978
rect 408498 478350 409118 495922
rect 408498 478294 408594 478350
rect 408650 478294 408718 478350
rect 408774 478294 408842 478350
rect 408898 478294 408966 478350
rect 409022 478294 409118 478350
rect 408498 478226 409118 478294
rect 408498 478170 408594 478226
rect 408650 478170 408718 478226
rect 408774 478170 408842 478226
rect 408898 478170 408966 478226
rect 409022 478170 409118 478226
rect 408498 478102 409118 478170
rect 408498 478046 408594 478102
rect 408650 478046 408718 478102
rect 408774 478046 408842 478102
rect 408898 478046 408966 478102
rect 409022 478046 409118 478102
rect 408498 477978 409118 478046
rect 408498 477922 408594 477978
rect 408650 477922 408718 477978
rect 408774 477922 408842 477978
rect 408898 477922 408966 477978
rect 409022 477922 409118 477978
rect 408498 460350 409118 477922
rect 408498 460294 408594 460350
rect 408650 460294 408718 460350
rect 408774 460294 408842 460350
rect 408898 460294 408966 460350
rect 409022 460294 409118 460350
rect 408498 460226 409118 460294
rect 408498 460170 408594 460226
rect 408650 460170 408718 460226
rect 408774 460170 408842 460226
rect 408898 460170 408966 460226
rect 409022 460170 409118 460226
rect 408498 460102 409118 460170
rect 408498 460046 408594 460102
rect 408650 460046 408718 460102
rect 408774 460046 408842 460102
rect 408898 460046 408966 460102
rect 409022 460046 409118 460102
rect 408498 459978 409118 460046
rect 408498 459922 408594 459978
rect 408650 459922 408718 459978
rect 408774 459922 408842 459978
rect 408898 459922 408966 459978
rect 409022 459922 409118 459978
rect 408498 442350 409118 459922
rect 408498 442294 408594 442350
rect 408650 442294 408718 442350
rect 408774 442294 408842 442350
rect 408898 442294 408966 442350
rect 409022 442294 409118 442350
rect 408498 442226 409118 442294
rect 408498 442170 408594 442226
rect 408650 442170 408718 442226
rect 408774 442170 408842 442226
rect 408898 442170 408966 442226
rect 409022 442170 409118 442226
rect 408498 442102 409118 442170
rect 408498 442046 408594 442102
rect 408650 442046 408718 442102
rect 408774 442046 408842 442102
rect 408898 442046 408966 442102
rect 409022 442046 409118 442102
rect 408498 441978 409118 442046
rect 408498 441922 408594 441978
rect 408650 441922 408718 441978
rect 408774 441922 408842 441978
rect 408898 441922 408966 441978
rect 409022 441922 409118 441978
rect 408498 424350 409118 441922
rect 408498 424294 408594 424350
rect 408650 424294 408718 424350
rect 408774 424294 408842 424350
rect 408898 424294 408966 424350
rect 409022 424294 409118 424350
rect 408498 424226 409118 424294
rect 408498 424170 408594 424226
rect 408650 424170 408718 424226
rect 408774 424170 408842 424226
rect 408898 424170 408966 424226
rect 409022 424170 409118 424226
rect 408498 424102 409118 424170
rect 408498 424046 408594 424102
rect 408650 424046 408718 424102
rect 408774 424046 408842 424102
rect 408898 424046 408966 424102
rect 409022 424046 409118 424102
rect 408498 423978 409118 424046
rect 408498 423922 408594 423978
rect 408650 423922 408718 423978
rect 408774 423922 408842 423978
rect 408898 423922 408966 423978
rect 409022 423922 409118 423978
rect 408498 406350 409118 423922
rect 408498 406294 408594 406350
rect 408650 406294 408718 406350
rect 408774 406294 408842 406350
rect 408898 406294 408966 406350
rect 409022 406294 409118 406350
rect 408498 406226 409118 406294
rect 408498 406170 408594 406226
rect 408650 406170 408718 406226
rect 408774 406170 408842 406226
rect 408898 406170 408966 406226
rect 409022 406170 409118 406226
rect 408498 406102 409118 406170
rect 408498 406046 408594 406102
rect 408650 406046 408718 406102
rect 408774 406046 408842 406102
rect 408898 406046 408966 406102
rect 409022 406046 409118 406102
rect 408498 405978 409118 406046
rect 408498 405922 408594 405978
rect 408650 405922 408718 405978
rect 408774 405922 408842 405978
rect 408898 405922 408966 405978
rect 409022 405922 409118 405978
rect 408498 388350 409118 405922
rect 408498 388294 408594 388350
rect 408650 388294 408718 388350
rect 408774 388294 408842 388350
rect 408898 388294 408966 388350
rect 409022 388294 409118 388350
rect 408498 388226 409118 388294
rect 408498 388170 408594 388226
rect 408650 388170 408718 388226
rect 408774 388170 408842 388226
rect 408898 388170 408966 388226
rect 409022 388170 409118 388226
rect 408498 388102 409118 388170
rect 408498 388046 408594 388102
rect 408650 388046 408718 388102
rect 408774 388046 408842 388102
rect 408898 388046 408966 388102
rect 409022 388046 409118 388102
rect 408498 387978 409118 388046
rect 408498 387922 408594 387978
rect 408650 387922 408718 387978
rect 408774 387922 408842 387978
rect 408898 387922 408966 387978
rect 409022 387922 409118 387978
rect 408498 370350 409118 387922
rect 408498 370294 408594 370350
rect 408650 370294 408718 370350
rect 408774 370294 408842 370350
rect 408898 370294 408966 370350
rect 409022 370294 409118 370350
rect 408498 370226 409118 370294
rect 408498 370170 408594 370226
rect 408650 370170 408718 370226
rect 408774 370170 408842 370226
rect 408898 370170 408966 370226
rect 409022 370170 409118 370226
rect 408498 370102 409118 370170
rect 408498 370046 408594 370102
rect 408650 370046 408718 370102
rect 408774 370046 408842 370102
rect 408898 370046 408966 370102
rect 409022 370046 409118 370102
rect 408498 369978 409118 370046
rect 408498 369922 408594 369978
rect 408650 369922 408718 369978
rect 408774 369922 408842 369978
rect 408898 369922 408966 369978
rect 409022 369922 409118 369978
rect 408498 352350 409118 369922
rect 408498 352294 408594 352350
rect 408650 352294 408718 352350
rect 408774 352294 408842 352350
rect 408898 352294 408966 352350
rect 409022 352294 409118 352350
rect 408498 352226 409118 352294
rect 408498 352170 408594 352226
rect 408650 352170 408718 352226
rect 408774 352170 408842 352226
rect 408898 352170 408966 352226
rect 409022 352170 409118 352226
rect 408498 352102 409118 352170
rect 408498 352046 408594 352102
rect 408650 352046 408718 352102
rect 408774 352046 408842 352102
rect 408898 352046 408966 352102
rect 409022 352046 409118 352102
rect 408498 351978 409118 352046
rect 408498 351922 408594 351978
rect 408650 351922 408718 351978
rect 408774 351922 408842 351978
rect 408898 351922 408966 351978
rect 409022 351922 409118 351978
rect 408498 334350 409118 351922
rect 408498 334294 408594 334350
rect 408650 334294 408718 334350
rect 408774 334294 408842 334350
rect 408898 334294 408966 334350
rect 409022 334294 409118 334350
rect 408498 334226 409118 334294
rect 408498 334170 408594 334226
rect 408650 334170 408718 334226
rect 408774 334170 408842 334226
rect 408898 334170 408966 334226
rect 409022 334170 409118 334226
rect 408498 334102 409118 334170
rect 408498 334046 408594 334102
rect 408650 334046 408718 334102
rect 408774 334046 408842 334102
rect 408898 334046 408966 334102
rect 409022 334046 409118 334102
rect 408498 333978 409118 334046
rect 408498 333922 408594 333978
rect 408650 333922 408718 333978
rect 408774 333922 408842 333978
rect 408898 333922 408966 333978
rect 409022 333922 409118 333978
rect 408498 316350 409118 333922
rect 408498 316294 408594 316350
rect 408650 316294 408718 316350
rect 408774 316294 408842 316350
rect 408898 316294 408966 316350
rect 409022 316294 409118 316350
rect 408498 316226 409118 316294
rect 408498 316170 408594 316226
rect 408650 316170 408718 316226
rect 408774 316170 408842 316226
rect 408898 316170 408966 316226
rect 409022 316170 409118 316226
rect 408498 316102 409118 316170
rect 408498 316046 408594 316102
rect 408650 316046 408718 316102
rect 408774 316046 408842 316102
rect 408898 316046 408966 316102
rect 409022 316046 409118 316102
rect 408498 315978 409118 316046
rect 408498 315922 408594 315978
rect 408650 315922 408718 315978
rect 408774 315922 408842 315978
rect 408898 315922 408966 315978
rect 409022 315922 409118 315978
rect 408498 298350 409118 315922
rect 408498 298294 408594 298350
rect 408650 298294 408718 298350
rect 408774 298294 408842 298350
rect 408898 298294 408966 298350
rect 409022 298294 409118 298350
rect 408498 298226 409118 298294
rect 408498 298170 408594 298226
rect 408650 298170 408718 298226
rect 408774 298170 408842 298226
rect 408898 298170 408966 298226
rect 409022 298170 409118 298226
rect 408498 298102 409118 298170
rect 408498 298046 408594 298102
rect 408650 298046 408718 298102
rect 408774 298046 408842 298102
rect 408898 298046 408966 298102
rect 409022 298046 409118 298102
rect 408498 297978 409118 298046
rect 408498 297922 408594 297978
rect 408650 297922 408718 297978
rect 408774 297922 408842 297978
rect 408898 297922 408966 297978
rect 409022 297922 409118 297978
rect 408498 280350 409118 297922
rect 408498 280294 408594 280350
rect 408650 280294 408718 280350
rect 408774 280294 408842 280350
rect 408898 280294 408966 280350
rect 409022 280294 409118 280350
rect 408498 280226 409118 280294
rect 408498 280170 408594 280226
rect 408650 280170 408718 280226
rect 408774 280170 408842 280226
rect 408898 280170 408966 280226
rect 409022 280170 409118 280226
rect 408498 280102 409118 280170
rect 408498 280046 408594 280102
rect 408650 280046 408718 280102
rect 408774 280046 408842 280102
rect 408898 280046 408966 280102
rect 409022 280046 409118 280102
rect 408498 279978 409118 280046
rect 408498 279922 408594 279978
rect 408650 279922 408718 279978
rect 408774 279922 408842 279978
rect 408898 279922 408966 279978
rect 409022 279922 409118 279978
rect 408498 262350 409118 279922
rect 408498 262294 408594 262350
rect 408650 262294 408718 262350
rect 408774 262294 408842 262350
rect 408898 262294 408966 262350
rect 409022 262294 409118 262350
rect 408498 262226 409118 262294
rect 408498 262170 408594 262226
rect 408650 262170 408718 262226
rect 408774 262170 408842 262226
rect 408898 262170 408966 262226
rect 409022 262170 409118 262226
rect 408498 262102 409118 262170
rect 408498 262046 408594 262102
rect 408650 262046 408718 262102
rect 408774 262046 408842 262102
rect 408898 262046 408966 262102
rect 409022 262046 409118 262102
rect 408498 261978 409118 262046
rect 408498 261922 408594 261978
rect 408650 261922 408718 261978
rect 408774 261922 408842 261978
rect 408898 261922 408966 261978
rect 409022 261922 409118 261978
rect 408498 244350 409118 261922
rect 408498 244294 408594 244350
rect 408650 244294 408718 244350
rect 408774 244294 408842 244350
rect 408898 244294 408966 244350
rect 409022 244294 409118 244350
rect 408498 244226 409118 244294
rect 408498 244170 408594 244226
rect 408650 244170 408718 244226
rect 408774 244170 408842 244226
rect 408898 244170 408966 244226
rect 409022 244170 409118 244226
rect 408498 244102 409118 244170
rect 408498 244046 408594 244102
rect 408650 244046 408718 244102
rect 408774 244046 408842 244102
rect 408898 244046 408966 244102
rect 409022 244046 409118 244102
rect 408498 243978 409118 244046
rect 408498 243922 408594 243978
rect 408650 243922 408718 243978
rect 408774 243922 408842 243978
rect 408898 243922 408966 243978
rect 409022 243922 409118 243978
rect 408498 226350 409118 243922
rect 408498 226294 408594 226350
rect 408650 226294 408718 226350
rect 408774 226294 408842 226350
rect 408898 226294 408966 226350
rect 409022 226294 409118 226350
rect 408498 226226 409118 226294
rect 408498 226170 408594 226226
rect 408650 226170 408718 226226
rect 408774 226170 408842 226226
rect 408898 226170 408966 226226
rect 409022 226170 409118 226226
rect 408498 226102 409118 226170
rect 408498 226046 408594 226102
rect 408650 226046 408718 226102
rect 408774 226046 408842 226102
rect 408898 226046 408966 226102
rect 409022 226046 409118 226102
rect 408498 225978 409118 226046
rect 408498 225922 408594 225978
rect 408650 225922 408718 225978
rect 408774 225922 408842 225978
rect 408898 225922 408966 225978
rect 409022 225922 409118 225978
rect 408498 208350 409118 225922
rect 408498 208294 408594 208350
rect 408650 208294 408718 208350
rect 408774 208294 408842 208350
rect 408898 208294 408966 208350
rect 409022 208294 409118 208350
rect 408498 208226 409118 208294
rect 408498 208170 408594 208226
rect 408650 208170 408718 208226
rect 408774 208170 408842 208226
rect 408898 208170 408966 208226
rect 409022 208170 409118 208226
rect 408498 208102 409118 208170
rect 408498 208046 408594 208102
rect 408650 208046 408718 208102
rect 408774 208046 408842 208102
rect 408898 208046 408966 208102
rect 409022 208046 409118 208102
rect 408498 207978 409118 208046
rect 408498 207922 408594 207978
rect 408650 207922 408718 207978
rect 408774 207922 408842 207978
rect 408898 207922 408966 207978
rect 409022 207922 409118 207978
rect 408498 190350 409118 207922
rect 408498 190294 408594 190350
rect 408650 190294 408718 190350
rect 408774 190294 408842 190350
rect 408898 190294 408966 190350
rect 409022 190294 409118 190350
rect 408498 190226 409118 190294
rect 408498 190170 408594 190226
rect 408650 190170 408718 190226
rect 408774 190170 408842 190226
rect 408898 190170 408966 190226
rect 409022 190170 409118 190226
rect 408498 190102 409118 190170
rect 408498 190046 408594 190102
rect 408650 190046 408718 190102
rect 408774 190046 408842 190102
rect 408898 190046 408966 190102
rect 409022 190046 409118 190102
rect 408498 189978 409118 190046
rect 408498 189922 408594 189978
rect 408650 189922 408718 189978
rect 408774 189922 408842 189978
rect 408898 189922 408966 189978
rect 409022 189922 409118 189978
rect 408498 172350 409118 189922
rect 408498 172294 408594 172350
rect 408650 172294 408718 172350
rect 408774 172294 408842 172350
rect 408898 172294 408966 172350
rect 409022 172294 409118 172350
rect 408498 172226 409118 172294
rect 408498 172170 408594 172226
rect 408650 172170 408718 172226
rect 408774 172170 408842 172226
rect 408898 172170 408966 172226
rect 409022 172170 409118 172226
rect 408498 172102 409118 172170
rect 408498 172046 408594 172102
rect 408650 172046 408718 172102
rect 408774 172046 408842 172102
rect 408898 172046 408966 172102
rect 409022 172046 409118 172102
rect 408498 171978 409118 172046
rect 408498 171922 408594 171978
rect 408650 171922 408718 171978
rect 408774 171922 408842 171978
rect 408898 171922 408966 171978
rect 409022 171922 409118 171978
rect 408498 154350 409118 171922
rect 408498 154294 408594 154350
rect 408650 154294 408718 154350
rect 408774 154294 408842 154350
rect 408898 154294 408966 154350
rect 409022 154294 409118 154350
rect 408498 154226 409118 154294
rect 408498 154170 408594 154226
rect 408650 154170 408718 154226
rect 408774 154170 408842 154226
rect 408898 154170 408966 154226
rect 409022 154170 409118 154226
rect 408498 154102 409118 154170
rect 408498 154046 408594 154102
rect 408650 154046 408718 154102
rect 408774 154046 408842 154102
rect 408898 154046 408966 154102
rect 409022 154046 409118 154102
rect 408498 153978 409118 154046
rect 408498 153922 408594 153978
rect 408650 153922 408718 153978
rect 408774 153922 408842 153978
rect 408898 153922 408966 153978
rect 409022 153922 409118 153978
rect 408498 136350 409118 153922
rect 408498 136294 408594 136350
rect 408650 136294 408718 136350
rect 408774 136294 408842 136350
rect 408898 136294 408966 136350
rect 409022 136294 409118 136350
rect 408498 136226 409118 136294
rect 408498 136170 408594 136226
rect 408650 136170 408718 136226
rect 408774 136170 408842 136226
rect 408898 136170 408966 136226
rect 409022 136170 409118 136226
rect 408498 136102 409118 136170
rect 408498 136046 408594 136102
rect 408650 136046 408718 136102
rect 408774 136046 408842 136102
rect 408898 136046 408966 136102
rect 409022 136046 409118 136102
rect 408498 135978 409118 136046
rect 408498 135922 408594 135978
rect 408650 135922 408718 135978
rect 408774 135922 408842 135978
rect 408898 135922 408966 135978
rect 409022 135922 409118 135978
rect 408498 118350 409118 135922
rect 408498 118294 408594 118350
rect 408650 118294 408718 118350
rect 408774 118294 408842 118350
rect 408898 118294 408966 118350
rect 409022 118294 409118 118350
rect 408498 118226 409118 118294
rect 408498 118170 408594 118226
rect 408650 118170 408718 118226
rect 408774 118170 408842 118226
rect 408898 118170 408966 118226
rect 409022 118170 409118 118226
rect 408498 118102 409118 118170
rect 408498 118046 408594 118102
rect 408650 118046 408718 118102
rect 408774 118046 408842 118102
rect 408898 118046 408966 118102
rect 409022 118046 409118 118102
rect 408498 117978 409118 118046
rect 408498 117922 408594 117978
rect 408650 117922 408718 117978
rect 408774 117922 408842 117978
rect 408898 117922 408966 117978
rect 409022 117922 409118 117978
rect 408498 100350 409118 117922
rect 408498 100294 408594 100350
rect 408650 100294 408718 100350
rect 408774 100294 408842 100350
rect 408898 100294 408966 100350
rect 409022 100294 409118 100350
rect 408498 100226 409118 100294
rect 408498 100170 408594 100226
rect 408650 100170 408718 100226
rect 408774 100170 408842 100226
rect 408898 100170 408966 100226
rect 409022 100170 409118 100226
rect 408498 100102 409118 100170
rect 408498 100046 408594 100102
rect 408650 100046 408718 100102
rect 408774 100046 408842 100102
rect 408898 100046 408966 100102
rect 409022 100046 409118 100102
rect 408498 99978 409118 100046
rect 408498 99922 408594 99978
rect 408650 99922 408718 99978
rect 408774 99922 408842 99978
rect 408898 99922 408966 99978
rect 409022 99922 409118 99978
rect 408498 82350 409118 99922
rect 408498 82294 408594 82350
rect 408650 82294 408718 82350
rect 408774 82294 408842 82350
rect 408898 82294 408966 82350
rect 409022 82294 409118 82350
rect 408498 82226 409118 82294
rect 408498 82170 408594 82226
rect 408650 82170 408718 82226
rect 408774 82170 408842 82226
rect 408898 82170 408966 82226
rect 409022 82170 409118 82226
rect 408498 82102 409118 82170
rect 408498 82046 408594 82102
rect 408650 82046 408718 82102
rect 408774 82046 408842 82102
rect 408898 82046 408966 82102
rect 409022 82046 409118 82102
rect 408498 81978 409118 82046
rect 408498 81922 408594 81978
rect 408650 81922 408718 81978
rect 408774 81922 408842 81978
rect 408898 81922 408966 81978
rect 409022 81922 409118 81978
rect 404778 58294 404874 58350
rect 404930 58294 404998 58350
rect 405054 58294 405122 58350
rect 405178 58294 405246 58350
rect 405302 58294 405398 58350
rect 404778 58226 405398 58294
rect 404778 58170 404874 58226
rect 404930 58170 404998 58226
rect 405054 58170 405122 58226
rect 405178 58170 405246 58226
rect 405302 58170 405398 58226
rect 404778 58102 405398 58170
rect 404778 58046 404874 58102
rect 404930 58046 404998 58102
rect 405054 58046 405122 58102
rect 405178 58046 405246 58102
rect 405302 58046 405398 58102
rect 404778 57978 405398 58046
rect 404778 57922 404874 57978
rect 404930 57922 404998 57978
rect 405054 57922 405122 57978
rect 405178 57922 405246 57978
rect 405302 57922 405398 57978
rect 404778 40350 405398 57922
rect 404778 40294 404874 40350
rect 404930 40294 404998 40350
rect 405054 40294 405122 40350
rect 405178 40294 405246 40350
rect 405302 40294 405398 40350
rect 404778 40226 405398 40294
rect 404778 40170 404874 40226
rect 404930 40170 404998 40226
rect 405054 40170 405122 40226
rect 405178 40170 405246 40226
rect 405302 40170 405398 40226
rect 404778 40102 405398 40170
rect 404778 40046 404874 40102
rect 404930 40046 404998 40102
rect 405054 40046 405122 40102
rect 405178 40046 405246 40102
rect 405302 40046 405398 40102
rect 404778 39978 405398 40046
rect 404778 39922 404874 39978
rect 404930 39922 404998 39978
rect 405054 39922 405122 39978
rect 405178 39922 405246 39978
rect 405302 39922 405398 39978
rect 396508 4162 396564 4172
rect 403228 33778 403284 33788
rect 403228 4228 403284 33722
rect 403228 4162 403284 4172
rect 404778 22350 405398 39922
rect 404778 22294 404874 22350
rect 404930 22294 404998 22350
rect 405054 22294 405122 22350
rect 405178 22294 405246 22350
rect 405302 22294 405398 22350
rect 404778 22226 405398 22294
rect 404778 22170 404874 22226
rect 404930 22170 404998 22226
rect 405054 22170 405122 22226
rect 405178 22170 405246 22226
rect 405302 22170 405398 22226
rect 404778 22102 405398 22170
rect 404778 22046 404874 22102
rect 404930 22046 404998 22102
rect 405054 22046 405122 22102
rect 405178 22046 405246 22102
rect 405302 22046 405398 22102
rect 404778 21978 405398 22046
rect 404778 21922 404874 21978
rect 404930 21922 404998 21978
rect 405054 21922 405122 21978
rect 405178 21922 405246 21978
rect 405302 21922 405398 21978
rect 404778 4350 405398 21922
rect 404778 4294 404874 4350
rect 404930 4294 404998 4350
rect 405054 4294 405122 4350
rect 405178 4294 405246 4350
rect 405302 4294 405398 4350
rect 404778 4226 405398 4294
rect 404778 4170 404874 4226
rect 404930 4170 404998 4226
rect 405054 4170 405122 4226
rect 405178 4170 405246 4226
rect 405302 4170 405398 4226
rect 377778 -1176 377874 -1120
rect 377930 -1176 377998 -1120
rect 378054 -1176 378122 -1120
rect 378178 -1176 378246 -1120
rect 378302 -1176 378398 -1120
rect 377778 -1244 378398 -1176
rect 377778 -1300 377874 -1244
rect 377930 -1300 377998 -1244
rect 378054 -1300 378122 -1244
rect 378178 -1300 378246 -1244
rect 378302 -1300 378398 -1244
rect 377778 -1368 378398 -1300
rect 377778 -1424 377874 -1368
rect 377930 -1424 377998 -1368
rect 378054 -1424 378122 -1368
rect 378178 -1424 378246 -1368
rect 378302 -1424 378398 -1368
rect 377778 -1492 378398 -1424
rect 377778 -1548 377874 -1492
rect 377930 -1548 377998 -1492
rect 378054 -1548 378122 -1492
rect 378178 -1548 378246 -1492
rect 378302 -1548 378398 -1492
rect 377778 -1644 378398 -1548
rect 404778 4102 405398 4170
rect 406588 65818 406644 65828
rect 406588 4228 406644 65762
rect 406588 4162 406644 4172
rect 408498 64350 409118 81922
rect 435498 597212 436118 598268
rect 435498 597156 435594 597212
rect 435650 597156 435718 597212
rect 435774 597156 435842 597212
rect 435898 597156 435966 597212
rect 436022 597156 436118 597212
rect 435498 597088 436118 597156
rect 435498 597032 435594 597088
rect 435650 597032 435718 597088
rect 435774 597032 435842 597088
rect 435898 597032 435966 597088
rect 436022 597032 436118 597088
rect 435498 596964 436118 597032
rect 435498 596908 435594 596964
rect 435650 596908 435718 596964
rect 435774 596908 435842 596964
rect 435898 596908 435966 596964
rect 436022 596908 436118 596964
rect 435498 596840 436118 596908
rect 435498 596784 435594 596840
rect 435650 596784 435718 596840
rect 435774 596784 435842 596840
rect 435898 596784 435966 596840
rect 436022 596784 436118 596840
rect 435498 580350 436118 596784
rect 435498 580294 435594 580350
rect 435650 580294 435718 580350
rect 435774 580294 435842 580350
rect 435898 580294 435966 580350
rect 436022 580294 436118 580350
rect 435498 580226 436118 580294
rect 435498 580170 435594 580226
rect 435650 580170 435718 580226
rect 435774 580170 435842 580226
rect 435898 580170 435966 580226
rect 436022 580170 436118 580226
rect 435498 580102 436118 580170
rect 435498 580046 435594 580102
rect 435650 580046 435718 580102
rect 435774 580046 435842 580102
rect 435898 580046 435966 580102
rect 436022 580046 436118 580102
rect 435498 579978 436118 580046
rect 435498 579922 435594 579978
rect 435650 579922 435718 579978
rect 435774 579922 435842 579978
rect 435898 579922 435966 579978
rect 436022 579922 436118 579978
rect 435498 562350 436118 579922
rect 435498 562294 435594 562350
rect 435650 562294 435718 562350
rect 435774 562294 435842 562350
rect 435898 562294 435966 562350
rect 436022 562294 436118 562350
rect 435498 562226 436118 562294
rect 435498 562170 435594 562226
rect 435650 562170 435718 562226
rect 435774 562170 435842 562226
rect 435898 562170 435966 562226
rect 436022 562170 436118 562226
rect 435498 562102 436118 562170
rect 435498 562046 435594 562102
rect 435650 562046 435718 562102
rect 435774 562046 435842 562102
rect 435898 562046 435966 562102
rect 436022 562046 436118 562102
rect 435498 561978 436118 562046
rect 435498 561922 435594 561978
rect 435650 561922 435718 561978
rect 435774 561922 435842 561978
rect 435898 561922 435966 561978
rect 436022 561922 436118 561978
rect 435498 544350 436118 561922
rect 435498 544294 435594 544350
rect 435650 544294 435718 544350
rect 435774 544294 435842 544350
rect 435898 544294 435966 544350
rect 436022 544294 436118 544350
rect 435498 544226 436118 544294
rect 435498 544170 435594 544226
rect 435650 544170 435718 544226
rect 435774 544170 435842 544226
rect 435898 544170 435966 544226
rect 436022 544170 436118 544226
rect 435498 544102 436118 544170
rect 435498 544046 435594 544102
rect 435650 544046 435718 544102
rect 435774 544046 435842 544102
rect 435898 544046 435966 544102
rect 436022 544046 436118 544102
rect 435498 543978 436118 544046
rect 435498 543922 435594 543978
rect 435650 543922 435718 543978
rect 435774 543922 435842 543978
rect 435898 543922 435966 543978
rect 436022 543922 436118 543978
rect 435498 526350 436118 543922
rect 435498 526294 435594 526350
rect 435650 526294 435718 526350
rect 435774 526294 435842 526350
rect 435898 526294 435966 526350
rect 436022 526294 436118 526350
rect 435498 526226 436118 526294
rect 435498 526170 435594 526226
rect 435650 526170 435718 526226
rect 435774 526170 435842 526226
rect 435898 526170 435966 526226
rect 436022 526170 436118 526226
rect 435498 526102 436118 526170
rect 435498 526046 435594 526102
rect 435650 526046 435718 526102
rect 435774 526046 435842 526102
rect 435898 526046 435966 526102
rect 436022 526046 436118 526102
rect 435498 525978 436118 526046
rect 435498 525922 435594 525978
rect 435650 525922 435718 525978
rect 435774 525922 435842 525978
rect 435898 525922 435966 525978
rect 436022 525922 436118 525978
rect 435498 508350 436118 525922
rect 435498 508294 435594 508350
rect 435650 508294 435718 508350
rect 435774 508294 435842 508350
rect 435898 508294 435966 508350
rect 436022 508294 436118 508350
rect 435498 508226 436118 508294
rect 435498 508170 435594 508226
rect 435650 508170 435718 508226
rect 435774 508170 435842 508226
rect 435898 508170 435966 508226
rect 436022 508170 436118 508226
rect 435498 508102 436118 508170
rect 435498 508046 435594 508102
rect 435650 508046 435718 508102
rect 435774 508046 435842 508102
rect 435898 508046 435966 508102
rect 436022 508046 436118 508102
rect 435498 507978 436118 508046
rect 435498 507922 435594 507978
rect 435650 507922 435718 507978
rect 435774 507922 435842 507978
rect 435898 507922 435966 507978
rect 436022 507922 436118 507978
rect 435498 490350 436118 507922
rect 435498 490294 435594 490350
rect 435650 490294 435718 490350
rect 435774 490294 435842 490350
rect 435898 490294 435966 490350
rect 436022 490294 436118 490350
rect 435498 490226 436118 490294
rect 435498 490170 435594 490226
rect 435650 490170 435718 490226
rect 435774 490170 435842 490226
rect 435898 490170 435966 490226
rect 436022 490170 436118 490226
rect 435498 490102 436118 490170
rect 435498 490046 435594 490102
rect 435650 490046 435718 490102
rect 435774 490046 435842 490102
rect 435898 490046 435966 490102
rect 436022 490046 436118 490102
rect 435498 489978 436118 490046
rect 435498 489922 435594 489978
rect 435650 489922 435718 489978
rect 435774 489922 435842 489978
rect 435898 489922 435966 489978
rect 436022 489922 436118 489978
rect 435498 472350 436118 489922
rect 435498 472294 435594 472350
rect 435650 472294 435718 472350
rect 435774 472294 435842 472350
rect 435898 472294 435966 472350
rect 436022 472294 436118 472350
rect 435498 472226 436118 472294
rect 435498 472170 435594 472226
rect 435650 472170 435718 472226
rect 435774 472170 435842 472226
rect 435898 472170 435966 472226
rect 436022 472170 436118 472226
rect 435498 472102 436118 472170
rect 435498 472046 435594 472102
rect 435650 472046 435718 472102
rect 435774 472046 435842 472102
rect 435898 472046 435966 472102
rect 436022 472046 436118 472102
rect 435498 471978 436118 472046
rect 435498 471922 435594 471978
rect 435650 471922 435718 471978
rect 435774 471922 435842 471978
rect 435898 471922 435966 471978
rect 436022 471922 436118 471978
rect 435498 454350 436118 471922
rect 435498 454294 435594 454350
rect 435650 454294 435718 454350
rect 435774 454294 435842 454350
rect 435898 454294 435966 454350
rect 436022 454294 436118 454350
rect 435498 454226 436118 454294
rect 435498 454170 435594 454226
rect 435650 454170 435718 454226
rect 435774 454170 435842 454226
rect 435898 454170 435966 454226
rect 436022 454170 436118 454226
rect 435498 454102 436118 454170
rect 435498 454046 435594 454102
rect 435650 454046 435718 454102
rect 435774 454046 435842 454102
rect 435898 454046 435966 454102
rect 436022 454046 436118 454102
rect 435498 453978 436118 454046
rect 435498 453922 435594 453978
rect 435650 453922 435718 453978
rect 435774 453922 435842 453978
rect 435898 453922 435966 453978
rect 436022 453922 436118 453978
rect 435498 436350 436118 453922
rect 435498 436294 435594 436350
rect 435650 436294 435718 436350
rect 435774 436294 435842 436350
rect 435898 436294 435966 436350
rect 436022 436294 436118 436350
rect 435498 436226 436118 436294
rect 435498 436170 435594 436226
rect 435650 436170 435718 436226
rect 435774 436170 435842 436226
rect 435898 436170 435966 436226
rect 436022 436170 436118 436226
rect 435498 436102 436118 436170
rect 435498 436046 435594 436102
rect 435650 436046 435718 436102
rect 435774 436046 435842 436102
rect 435898 436046 435966 436102
rect 436022 436046 436118 436102
rect 435498 435978 436118 436046
rect 435498 435922 435594 435978
rect 435650 435922 435718 435978
rect 435774 435922 435842 435978
rect 435898 435922 435966 435978
rect 436022 435922 436118 435978
rect 435498 418350 436118 435922
rect 435498 418294 435594 418350
rect 435650 418294 435718 418350
rect 435774 418294 435842 418350
rect 435898 418294 435966 418350
rect 436022 418294 436118 418350
rect 435498 418226 436118 418294
rect 435498 418170 435594 418226
rect 435650 418170 435718 418226
rect 435774 418170 435842 418226
rect 435898 418170 435966 418226
rect 436022 418170 436118 418226
rect 435498 418102 436118 418170
rect 435498 418046 435594 418102
rect 435650 418046 435718 418102
rect 435774 418046 435842 418102
rect 435898 418046 435966 418102
rect 436022 418046 436118 418102
rect 435498 417978 436118 418046
rect 435498 417922 435594 417978
rect 435650 417922 435718 417978
rect 435774 417922 435842 417978
rect 435898 417922 435966 417978
rect 436022 417922 436118 417978
rect 435498 400350 436118 417922
rect 435498 400294 435594 400350
rect 435650 400294 435718 400350
rect 435774 400294 435842 400350
rect 435898 400294 435966 400350
rect 436022 400294 436118 400350
rect 435498 400226 436118 400294
rect 435498 400170 435594 400226
rect 435650 400170 435718 400226
rect 435774 400170 435842 400226
rect 435898 400170 435966 400226
rect 436022 400170 436118 400226
rect 435498 400102 436118 400170
rect 435498 400046 435594 400102
rect 435650 400046 435718 400102
rect 435774 400046 435842 400102
rect 435898 400046 435966 400102
rect 436022 400046 436118 400102
rect 435498 399978 436118 400046
rect 435498 399922 435594 399978
rect 435650 399922 435718 399978
rect 435774 399922 435842 399978
rect 435898 399922 435966 399978
rect 436022 399922 436118 399978
rect 435498 382350 436118 399922
rect 435498 382294 435594 382350
rect 435650 382294 435718 382350
rect 435774 382294 435842 382350
rect 435898 382294 435966 382350
rect 436022 382294 436118 382350
rect 435498 382226 436118 382294
rect 435498 382170 435594 382226
rect 435650 382170 435718 382226
rect 435774 382170 435842 382226
rect 435898 382170 435966 382226
rect 436022 382170 436118 382226
rect 435498 382102 436118 382170
rect 435498 382046 435594 382102
rect 435650 382046 435718 382102
rect 435774 382046 435842 382102
rect 435898 382046 435966 382102
rect 436022 382046 436118 382102
rect 435498 381978 436118 382046
rect 435498 381922 435594 381978
rect 435650 381922 435718 381978
rect 435774 381922 435842 381978
rect 435898 381922 435966 381978
rect 436022 381922 436118 381978
rect 435498 364350 436118 381922
rect 435498 364294 435594 364350
rect 435650 364294 435718 364350
rect 435774 364294 435842 364350
rect 435898 364294 435966 364350
rect 436022 364294 436118 364350
rect 435498 364226 436118 364294
rect 435498 364170 435594 364226
rect 435650 364170 435718 364226
rect 435774 364170 435842 364226
rect 435898 364170 435966 364226
rect 436022 364170 436118 364226
rect 435498 364102 436118 364170
rect 435498 364046 435594 364102
rect 435650 364046 435718 364102
rect 435774 364046 435842 364102
rect 435898 364046 435966 364102
rect 436022 364046 436118 364102
rect 435498 363978 436118 364046
rect 435498 363922 435594 363978
rect 435650 363922 435718 363978
rect 435774 363922 435842 363978
rect 435898 363922 435966 363978
rect 436022 363922 436118 363978
rect 435498 346350 436118 363922
rect 435498 346294 435594 346350
rect 435650 346294 435718 346350
rect 435774 346294 435842 346350
rect 435898 346294 435966 346350
rect 436022 346294 436118 346350
rect 435498 346226 436118 346294
rect 435498 346170 435594 346226
rect 435650 346170 435718 346226
rect 435774 346170 435842 346226
rect 435898 346170 435966 346226
rect 436022 346170 436118 346226
rect 435498 346102 436118 346170
rect 435498 346046 435594 346102
rect 435650 346046 435718 346102
rect 435774 346046 435842 346102
rect 435898 346046 435966 346102
rect 436022 346046 436118 346102
rect 435498 345978 436118 346046
rect 435498 345922 435594 345978
rect 435650 345922 435718 345978
rect 435774 345922 435842 345978
rect 435898 345922 435966 345978
rect 436022 345922 436118 345978
rect 435498 328350 436118 345922
rect 435498 328294 435594 328350
rect 435650 328294 435718 328350
rect 435774 328294 435842 328350
rect 435898 328294 435966 328350
rect 436022 328294 436118 328350
rect 435498 328226 436118 328294
rect 435498 328170 435594 328226
rect 435650 328170 435718 328226
rect 435774 328170 435842 328226
rect 435898 328170 435966 328226
rect 436022 328170 436118 328226
rect 435498 328102 436118 328170
rect 435498 328046 435594 328102
rect 435650 328046 435718 328102
rect 435774 328046 435842 328102
rect 435898 328046 435966 328102
rect 436022 328046 436118 328102
rect 435498 327978 436118 328046
rect 435498 327922 435594 327978
rect 435650 327922 435718 327978
rect 435774 327922 435842 327978
rect 435898 327922 435966 327978
rect 436022 327922 436118 327978
rect 435498 310350 436118 327922
rect 435498 310294 435594 310350
rect 435650 310294 435718 310350
rect 435774 310294 435842 310350
rect 435898 310294 435966 310350
rect 436022 310294 436118 310350
rect 435498 310226 436118 310294
rect 435498 310170 435594 310226
rect 435650 310170 435718 310226
rect 435774 310170 435842 310226
rect 435898 310170 435966 310226
rect 436022 310170 436118 310226
rect 435498 310102 436118 310170
rect 435498 310046 435594 310102
rect 435650 310046 435718 310102
rect 435774 310046 435842 310102
rect 435898 310046 435966 310102
rect 436022 310046 436118 310102
rect 435498 309978 436118 310046
rect 435498 309922 435594 309978
rect 435650 309922 435718 309978
rect 435774 309922 435842 309978
rect 435898 309922 435966 309978
rect 436022 309922 436118 309978
rect 435498 292350 436118 309922
rect 435498 292294 435594 292350
rect 435650 292294 435718 292350
rect 435774 292294 435842 292350
rect 435898 292294 435966 292350
rect 436022 292294 436118 292350
rect 435498 292226 436118 292294
rect 435498 292170 435594 292226
rect 435650 292170 435718 292226
rect 435774 292170 435842 292226
rect 435898 292170 435966 292226
rect 436022 292170 436118 292226
rect 435498 292102 436118 292170
rect 435498 292046 435594 292102
rect 435650 292046 435718 292102
rect 435774 292046 435842 292102
rect 435898 292046 435966 292102
rect 436022 292046 436118 292102
rect 435498 291978 436118 292046
rect 435498 291922 435594 291978
rect 435650 291922 435718 291978
rect 435774 291922 435842 291978
rect 435898 291922 435966 291978
rect 436022 291922 436118 291978
rect 435498 274350 436118 291922
rect 435498 274294 435594 274350
rect 435650 274294 435718 274350
rect 435774 274294 435842 274350
rect 435898 274294 435966 274350
rect 436022 274294 436118 274350
rect 435498 274226 436118 274294
rect 435498 274170 435594 274226
rect 435650 274170 435718 274226
rect 435774 274170 435842 274226
rect 435898 274170 435966 274226
rect 436022 274170 436118 274226
rect 435498 274102 436118 274170
rect 435498 274046 435594 274102
rect 435650 274046 435718 274102
rect 435774 274046 435842 274102
rect 435898 274046 435966 274102
rect 436022 274046 436118 274102
rect 435498 273978 436118 274046
rect 435498 273922 435594 273978
rect 435650 273922 435718 273978
rect 435774 273922 435842 273978
rect 435898 273922 435966 273978
rect 436022 273922 436118 273978
rect 435498 256350 436118 273922
rect 435498 256294 435594 256350
rect 435650 256294 435718 256350
rect 435774 256294 435842 256350
rect 435898 256294 435966 256350
rect 436022 256294 436118 256350
rect 435498 256226 436118 256294
rect 435498 256170 435594 256226
rect 435650 256170 435718 256226
rect 435774 256170 435842 256226
rect 435898 256170 435966 256226
rect 436022 256170 436118 256226
rect 435498 256102 436118 256170
rect 435498 256046 435594 256102
rect 435650 256046 435718 256102
rect 435774 256046 435842 256102
rect 435898 256046 435966 256102
rect 436022 256046 436118 256102
rect 435498 255978 436118 256046
rect 435498 255922 435594 255978
rect 435650 255922 435718 255978
rect 435774 255922 435842 255978
rect 435898 255922 435966 255978
rect 436022 255922 436118 255978
rect 435498 238350 436118 255922
rect 435498 238294 435594 238350
rect 435650 238294 435718 238350
rect 435774 238294 435842 238350
rect 435898 238294 435966 238350
rect 436022 238294 436118 238350
rect 435498 238226 436118 238294
rect 435498 238170 435594 238226
rect 435650 238170 435718 238226
rect 435774 238170 435842 238226
rect 435898 238170 435966 238226
rect 436022 238170 436118 238226
rect 435498 238102 436118 238170
rect 435498 238046 435594 238102
rect 435650 238046 435718 238102
rect 435774 238046 435842 238102
rect 435898 238046 435966 238102
rect 436022 238046 436118 238102
rect 435498 237978 436118 238046
rect 435498 237922 435594 237978
rect 435650 237922 435718 237978
rect 435774 237922 435842 237978
rect 435898 237922 435966 237978
rect 436022 237922 436118 237978
rect 435498 220350 436118 237922
rect 435498 220294 435594 220350
rect 435650 220294 435718 220350
rect 435774 220294 435842 220350
rect 435898 220294 435966 220350
rect 436022 220294 436118 220350
rect 435498 220226 436118 220294
rect 435498 220170 435594 220226
rect 435650 220170 435718 220226
rect 435774 220170 435842 220226
rect 435898 220170 435966 220226
rect 436022 220170 436118 220226
rect 435498 220102 436118 220170
rect 435498 220046 435594 220102
rect 435650 220046 435718 220102
rect 435774 220046 435842 220102
rect 435898 220046 435966 220102
rect 436022 220046 436118 220102
rect 435498 219978 436118 220046
rect 435498 219922 435594 219978
rect 435650 219922 435718 219978
rect 435774 219922 435842 219978
rect 435898 219922 435966 219978
rect 436022 219922 436118 219978
rect 435498 202350 436118 219922
rect 435498 202294 435594 202350
rect 435650 202294 435718 202350
rect 435774 202294 435842 202350
rect 435898 202294 435966 202350
rect 436022 202294 436118 202350
rect 435498 202226 436118 202294
rect 435498 202170 435594 202226
rect 435650 202170 435718 202226
rect 435774 202170 435842 202226
rect 435898 202170 435966 202226
rect 436022 202170 436118 202226
rect 435498 202102 436118 202170
rect 435498 202046 435594 202102
rect 435650 202046 435718 202102
rect 435774 202046 435842 202102
rect 435898 202046 435966 202102
rect 436022 202046 436118 202102
rect 435498 201978 436118 202046
rect 435498 201922 435594 201978
rect 435650 201922 435718 201978
rect 435774 201922 435842 201978
rect 435898 201922 435966 201978
rect 436022 201922 436118 201978
rect 435498 184350 436118 201922
rect 435498 184294 435594 184350
rect 435650 184294 435718 184350
rect 435774 184294 435842 184350
rect 435898 184294 435966 184350
rect 436022 184294 436118 184350
rect 435498 184226 436118 184294
rect 435498 184170 435594 184226
rect 435650 184170 435718 184226
rect 435774 184170 435842 184226
rect 435898 184170 435966 184226
rect 436022 184170 436118 184226
rect 435498 184102 436118 184170
rect 435498 184046 435594 184102
rect 435650 184046 435718 184102
rect 435774 184046 435842 184102
rect 435898 184046 435966 184102
rect 436022 184046 436118 184102
rect 435498 183978 436118 184046
rect 435498 183922 435594 183978
rect 435650 183922 435718 183978
rect 435774 183922 435842 183978
rect 435898 183922 435966 183978
rect 436022 183922 436118 183978
rect 435498 166350 436118 183922
rect 435498 166294 435594 166350
rect 435650 166294 435718 166350
rect 435774 166294 435842 166350
rect 435898 166294 435966 166350
rect 436022 166294 436118 166350
rect 435498 166226 436118 166294
rect 435498 166170 435594 166226
rect 435650 166170 435718 166226
rect 435774 166170 435842 166226
rect 435898 166170 435966 166226
rect 436022 166170 436118 166226
rect 435498 166102 436118 166170
rect 435498 166046 435594 166102
rect 435650 166046 435718 166102
rect 435774 166046 435842 166102
rect 435898 166046 435966 166102
rect 436022 166046 436118 166102
rect 435498 165978 436118 166046
rect 435498 165922 435594 165978
rect 435650 165922 435718 165978
rect 435774 165922 435842 165978
rect 435898 165922 435966 165978
rect 436022 165922 436118 165978
rect 435498 148350 436118 165922
rect 435498 148294 435594 148350
rect 435650 148294 435718 148350
rect 435774 148294 435842 148350
rect 435898 148294 435966 148350
rect 436022 148294 436118 148350
rect 435498 148226 436118 148294
rect 435498 148170 435594 148226
rect 435650 148170 435718 148226
rect 435774 148170 435842 148226
rect 435898 148170 435966 148226
rect 436022 148170 436118 148226
rect 435498 148102 436118 148170
rect 435498 148046 435594 148102
rect 435650 148046 435718 148102
rect 435774 148046 435842 148102
rect 435898 148046 435966 148102
rect 436022 148046 436118 148102
rect 435498 147978 436118 148046
rect 435498 147922 435594 147978
rect 435650 147922 435718 147978
rect 435774 147922 435842 147978
rect 435898 147922 435966 147978
rect 436022 147922 436118 147978
rect 435498 130350 436118 147922
rect 435498 130294 435594 130350
rect 435650 130294 435718 130350
rect 435774 130294 435842 130350
rect 435898 130294 435966 130350
rect 436022 130294 436118 130350
rect 435498 130226 436118 130294
rect 435498 130170 435594 130226
rect 435650 130170 435718 130226
rect 435774 130170 435842 130226
rect 435898 130170 435966 130226
rect 436022 130170 436118 130226
rect 435498 130102 436118 130170
rect 435498 130046 435594 130102
rect 435650 130046 435718 130102
rect 435774 130046 435842 130102
rect 435898 130046 435966 130102
rect 436022 130046 436118 130102
rect 435498 129978 436118 130046
rect 435498 129922 435594 129978
rect 435650 129922 435718 129978
rect 435774 129922 435842 129978
rect 435898 129922 435966 129978
rect 436022 129922 436118 129978
rect 435498 112350 436118 129922
rect 435498 112294 435594 112350
rect 435650 112294 435718 112350
rect 435774 112294 435842 112350
rect 435898 112294 435966 112350
rect 436022 112294 436118 112350
rect 435498 112226 436118 112294
rect 435498 112170 435594 112226
rect 435650 112170 435718 112226
rect 435774 112170 435842 112226
rect 435898 112170 435966 112226
rect 436022 112170 436118 112226
rect 435498 112102 436118 112170
rect 435498 112046 435594 112102
rect 435650 112046 435718 112102
rect 435774 112046 435842 112102
rect 435898 112046 435966 112102
rect 436022 112046 436118 112102
rect 435498 111978 436118 112046
rect 435498 111922 435594 111978
rect 435650 111922 435718 111978
rect 435774 111922 435842 111978
rect 435898 111922 435966 111978
rect 436022 111922 436118 111978
rect 435498 94350 436118 111922
rect 435498 94294 435594 94350
rect 435650 94294 435718 94350
rect 435774 94294 435842 94350
rect 435898 94294 435966 94350
rect 436022 94294 436118 94350
rect 435498 94226 436118 94294
rect 435498 94170 435594 94226
rect 435650 94170 435718 94226
rect 435774 94170 435842 94226
rect 435898 94170 435966 94226
rect 436022 94170 436118 94226
rect 435498 94102 436118 94170
rect 435498 94046 435594 94102
rect 435650 94046 435718 94102
rect 435774 94046 435842 94102
rect 435898 94046 435966 94102
rect 436022 94046 436118 94102
rect 435498 93978 436118 94046
rect 435498 93922 435594 93978
rect 435650 93922 435718 93978
rect 435774 93922 435842 93978
rect 435898 93922 435966 93978
rect 436022 93922 436118 93978
rect 435498 76350 436118 93922
rect 435498 76294 435594 76350
rect 435650 76294 435718 76350
rect 435774 76294 435842 76350
rect 435898 76294 435966 76350
rect 436022 76294 436118 76350
rect 435498 76226 436118 76294
rect 435498 76170 435594 76226
rect 435650 76170 435718 76226
rect 435774 76170 435842 76226
rect 435898 76170 435966 76226
rect 436022 76170 436118 76226
rect 435498 76102 436118 76170
rect 435498 76046 435594 76102
rect 435650 76046 435718 76102
rect 435774 76046 435842 76102
rect 435898 76046 435966 76102
rect 436022 76046 436118 76102
rect 435498 75978 436118 76046
rect 435498 75922 435594 75978
rect 435650 75922 435718 75978
rect 435774 75922 435842 75978
rect 435898 75922 435966 75978
rect 436022 75922 436118 75978
rect 435148 72478 435204 72488
rect 408498 64294 408594 64350
rect 408650 64294 408718 64350
rect 408774 64294 408842 64350
rect 408898 64294 408966 64350
rect 409022 64294 409118 64350
rect 408498 64226 409118 64294
rect 408498 64170 408594 64226
rect 408650 64170 408718 64226
rect 408774 64170 408842 64226
rect 408898 64170 408966 64226
rect 409022 64170 409118 64226
rect 408498 64102 409118 64170
rect 408498 64046 408594 64102
rect 408650 64046 408718 64102
rect 408774 64046 408842 64102
rect 408898 64046 408966 64102
rect 409022 64046 409118 64102
rect 408498 63978 409118 64046
rect 408498 63922 408594 63978
rect 408650 63922 408718 63978
rect 408774 63922 408842 63978
rect 408898 63922 408966 63978
rect 409022 63922 409118 63978
rect 408498 46350 409118 63922
rect 408498 46294 408594 46350
rect 408650 46294 408718 46350
rect 408774 46294 408842 46350
rect 408898 46294 408966 46350
rect 409022 46294 409118 46350
rect 408498 46226 409118 46294
rect 408498 46170 408594 46226
rect 408650 46170 408718 46226
rect 408774 46170 408842 46226
rect 408898 46170 408966 46226
rect 409022 46170 409118 46226
rect 408498 46102 409118 46170
rect 408498 46046 408594 46102
rect 408650 46046 408718 46102
rect 408774 46046 408842 46102
rect 408898 46046 408966 46102
rect 409022 46046 409118 46102
rect 408498 45978 409118 46046
rect 408498 45922 408594 45978
rect 408650 45922 408718 45978
rect 408774 45922 408842 45978
rect 408898 45922 408966 45978
rect 409022 45922 409118 45978
rect 408498 28350 409118 45922
rect 431788 67438 431844 67448
rect 408498 28294 408594 28350
rect 408650 28294 408718 28350
rect 408774 28294 408842 28350
rect 408898 28294 408966 28350
rect 409022 28294 409118 28350
rect 408498 28226 409118 28294
rect 408498 28170 408594 28226
rect 408650 28170 408718 28226
rect 408774 28170 408842 28226
rect 408898 28170 408966 28226
rect 409022 28170 409118 28226
rect 408498 28102 409118 28170
rect 408498 28046 408594 28102
rect 408650 28046 408718 28102
rect 408774 28046 408842 28102
rect 408898 28046 408966 28102
rect 409022 28046 409118 28102
rect 408498 27978 409118 28046
rect 408498 27922 408594 27978
rect 408650 27922 408718 27978
rect 408774 27922 408842 27978
rect 408898 27922 408966 27978
rect 409022 27922 409118 27978
rect 408498 10350 409118 27922
rect 416668 42058 416724 42068
rect 416668 20188 416724 42002
rect 425068 35578 425124 35588
rect 420028 33958 420084 33968
rect 416668 20132 416948 20188
rect 408498 10294 408594 10350
rect 408650 10294 408718 10350
rect 408774 10294 408842 10350
rect 408898 10294 408966 10350
rect 409022 10294 409118 10350
rect 408498 10226 409118 10294
rect 408498 10170 408594 10226
rect 408650 10170 408718 10226
rect 408774 10170 408842 10226
rect 408898 10170 408966 10226
rect 409022 10170 409118 10226
rect 408498 10102 409118 10170
rect 408498 10046 408594 10102
rect 408650 10046 408718 10102
rect 408774 10046 408842 10102
rect 408898 10046 408966 10102
rect 409022 10046 409118 10102
rect 408498 9978 409118 10046
rect 408498 9922 408594 9978
rect 408650 9922 408718 9978
rect 408774 9922 408842 9978
rect 408898 9922 408966 9978
rect 409022 9922 409118 9978
rect 404778 4046 404874 4102
rect 404930 4046 404998 4102
rect 405054 4046 405122 4102
rect 405178 4046 405246 4102
rect 405302 4046 405398 4102
rect 404778 3978 405398 4046
rect 404778 3922 404874 3978
rect 404930 3922 404998 3978
rect 405054 3922 405122 3978
rect 405178 3922 405246 3978
rect 405302 3922 405398 3978
rect 404778 -160 405398 3922
rect 404778 -216 404874 -160
rect 404930 -216 404998 -160
rect 405054 -216 405122 -160
rect 405178 -216 405246 -160
rect 405302 -216 405398 -160
rect 404778 -284 405398 -216
rect 404778 -340 404874 -284
rect 404930 -340 404998 -284
rect 405054 -340 405122 -284
rect 405178 -340 405246 -284
rect 405302 -340 405398 -284
rect 404778 -408 405398 -340
rect 404778 -464 404874 -408
rect 404930 -464 404998 -408
rect 405054 -464 405122 -408
rect 405178 -464 405246 -408
rect 405302 -464 405398 -408
rect 404778 -532 405398 -464
rect 404778 -588 404874 -532
rect 404930 -588 404998 -532
rect 405054 -588 405122 -532
rect 405178 -588 405246 -532
rect 405302 -588 405398 -532
rect 404778 -1644 405398 -588
rect 408498 -1120 409118 9922
rect 409948 17038 410004 17048
rect 409276 5878 409332 5888
rect 409276 3444 409332 5822
rect 409948 4228 410004 16982
rect 409948 4162 410004 4172
rect 414988 5338 415044 5348
rect 409276 3378 409332 3388
rect 414988 3444 415044 5282
rect 416892 4228 416948 20132
rect 416892 4162 416948 4172
rect 420028 4228 420084 33902
rect 420028 4162 420084 4172
rect 422604 8758 422660 8768
rect 422604 4228 422660 8702
rect 422604 4162 422660 4172
rect 425068 4228 425124 35522
rect 425068 4162 425124 4172
rect 428428 28918 428484 28928
rect 428428 4228 428484 28862
rect 428428 4162 428484 4172
rect 431788 4228 431844 67382
rect 431788 4162 431844 4172
rect 435148 4228 435204 72422
rect 435148 4162 435204 4172
rect 435498 58350 436118 75922
rect 435498 58294 435594 58350
rect 435650 58294 435718 58350
rect 435774 58294 435842 58350
rect 435898 58294 435966 58350
rect 436022 58294 436118 58350
rect 435498 58226 436118 58294
rect 435498 58170 435594 58226
rect 435650 58170 435718 58226
rect 435774 58170 435842 58226
rect 435898 58170 435966 58226
rect 436022 58170 436118 58226
rect 435498 58102 436118 58170
rect 435498 58046 435594 58102
rect 435650 58046 435718 58102
rect 435774 58046 435842 58102
rect 435898 58046 435966 58102
rect 436022 58046 436118 58102
rect 435498 57978 436118 58046
rect 435498 57922 435594 57978
rect 435650 57922 435718 57978
rect 435774 57922 435842 57978
rect 435898 57922 435966 57978
rect 436022 57922 436118 57978
rect 435498 40350 436118 57922
rect 439218 598172 439838 598268
rect 439218 598116 439314 598172
rect 439370 598116 439438 598172
rect 439494 598116 439562 598172
rect 439618 598116 439686 598172
rect 439742 598116 439838 598172
rect 439218 598048 439838 598116
rect 439218 597992 439314 598048
rect 439370 597992 439438 598048
rect 439494 597992 439562 598048
rect 439618 597992 439686 598048
rect 439742 597992 439838 598048
rect 439218 597924 439838 597992
rect 439218 597868 439314 597924
rect 439370 597868 439438 597924
rect 439494 597868 439562 597924
rect 439618 597868 439686 597924
rect 439742 597868 439838 597924
rect 439218 597800 439838 597868
rect 439218 597744 439314 597800
rect 439370 597744 439438 597800
rect 439494 597744 439562 597800
rect 439618 597744 439686 597800
rect 439742 597744 439838 597800
rect 439218 586350 439838 597744
rect 439218 586294 439314 586350
rect 439370 586294 439438 586350
rect 439494 586294 439562 586350
rect 439618 586294 439686 586350
rect 439742 586294 439838 586350
rect 439218 586226 439838 586294
rect 439218 586170 439314 586226
rect 439370 586170 439438 586226
rect 439494 586170 439562 586226
rect 439618 586170 439686 586226
rect 439742 586170 439838 586226
rect 439218 586102 439838 586170
rect 439218 586046 439314 586102
rect 439370 586046 439438 586102
rect 439494 586046 439562 586102
rect 439618 586046 439686 586102
rect 439742 586046 439838 586102
rect 439218 585978 439838 586046
rect 439218 585922 439314 585978
rect 439370 585922 439438 585978
rect 439494 585922 439562 585978
rect 439618 585922 439686 585978
rect 439742 585922 439838 585978
rect 439218 568350 439838 585922
rect 439218 568294 439314 568350
rect 439370 568294 439438 568350
rect 439494 568294 439562 568350
rect 439618 568294 439686 568350
rect 439742 568294 439838 568350
rect 439218 568226 439838 568294
rect 439218 568170 439314 568226
rect 439370 568170 439438 568226
rect 439494 568170 439562 568226
rect 439618 568170 439686 568226
rect 439742 568170 439838 568226
rect 439218 568102 439838 568170
rect 439218 568046 439314 568102
rect 439370 568046 439438 568102
rect 439494 568046 439562 568102
rect 439618 568046 439686 568102
rect 439742 568046 439838 568102
rect 439218 567978 439838 568046
rect 439218 567922 439314 567978
rect 439370 567922 439438 567978
rect 439494 567922 439562 567978
rect 439618 567922 439686 567978
rect 439742 567922 439838 567978
rect 439218 550350 439838 567922
rect 439218 550294 439314 550350
rect 439370 550294 439438 550350
rect 439494 550294 439562 550350
rect 439618 550294 439686 550350
rect 439742 550294 439838 550350
rect 439218 550226 439838 550294
rect 439218 550170 439314 550226
rect 439370 550170 439438 550226
rect 439494 550170 439562 550226
rect 439618 550170 439686 550226
rect 439742 550170 439838 550226
rect 439218 550102 439838 550170
rect 439218 550046 439314 550102
rect 439370 550046 439438 550102
rect 439494 550046 439562 550102
rect 439618 550046 439686 550102
rect 439742 550046 439838 550102
rect 439218 549978 439838 550046
rect 439218 549922 439314 549978
rect 439370 549922 439438 549978
rect 439494 549922 439562 549978
rect 439618 549922 439686 549978
rect 439742 549922 439838 549978
rect 439218 532350 439838 549922
rect 439218 532294 439314 532350
rect 439370 532294 439438 532350
rect 439494 532294 439562 532350
rect 439618 532294 439686 532350
rect 439742 532294 439838 532350
rect 439218 532226 439838 532294
rect 439218 532170 439314 532226
rect 439370 532170 439438 532226
rect 439494 532170 439562 532226
rect 439618 532170 439686 532226
rect 439742 532170 439838 532226
rect 439218 532102 439838 532170
rect 439218 532046 439314 532102
rect 439370 532046 439438 532102
rect 439494 532046 439562 532102
rect 439618 532046 439686 532102
rect 439742 532046 439838 532102
rect 439218 531978 439838 532046
rect 439218 531922 439314 531978
rect 439370 531922 439438 531978
rect 439494 531922 439562 531978
rect 439618 531922 439686 531978
rect 439742 531922 439838 531978
rect 439218 514350 439838 531922
rect 439218 514294 439314 514350
rect 439370 514294 439438 514350
rect 439494 514294 439562 514350
rect 439618 514294 439686 514350
rect 439742 514294 439838 514350
rect 439218 514226 439838 514294
rect 439218 514170 439314 514226
rect 439370 514170 439438 514226
rect 439494 514170 439562 514226
rect 439618 514170 439686 514226
rect 439742 514170 439838 514226
rect 439218 514102 439838 514170
rect 439218 514046 439314 514102
rect 439370 514046 439438 514102
rect 439494 514046 439562 514102
rect 439618 514046 439686 514102
rect 439742 514046 439838 514102
rect 439218 513978 439838 514046
rect 439218 513922 439314 513978
rect 439370 513922 439438 513978
rect 439494 513922 439562 513978
rect 439618 513922 439686 513978
rect 439742 513922 439838 513978
rect 439218 496350 439838 513922
rect 439218 496294 439314 496350
rect 439370 496294 439438 496350
rect 439494 496294 439562 496350
rect 439618 496294 439686 496350
rect 439742 496294 439838 496350
rect 439218 496226 439838 496294
rect 439218 496170 439314 496226
rect 439370 496170 439438 496226
rect 439494 496170 439562 496226
rect 439618 496170 439686 496226
rect 439742 496170 439838 496226
rect 439218 496102 439838 496170
rect 439218 496046 439314 496102
rect 439370 496046 439438 496102
rect 439494 496046 439562 496102
rect 439618 496046 439686 496102
rect 439742 496046 439838 496102
rect 439218 495978 439838 496046
rect 439218 495922 439314 495978
rect 439370 495922 439438 495978
rect 439494 495922 439562 495978
rect 439618 495922 439686 495978
rect 439742 495922 439838 495978
rect 439218 478350 439838 495922
rect 439218 478294 439314 478350
rect 439370 478294 439438 478350
rect 439494 478294 439562 478350
rect 439618 478294 439686 478350
rect 439742 478294 439838 478350
rect 439218 478226 439838 478294
rect 439218 478170 439314 478226
rect 439370 478170 439438 478226
rect 439494 478170 439562 478226
rect 439618 478170 439686 478226
rect 439742 478170 439838 478226
rect 439218 478102 439838 478170
rect 439218 478046 439314 478102
rect 439370 478046 439438 478102
rect 439494 478046 439562 478102
rect 439618 478046 439686 478102
rect 439742 478046 439838 478102
rect 439218 477978 439838 478046
rect 439218 477922 439314 477978
rect 439370 477922 439438 477978
rect 439494 477922 439562 477978
rect 439618 477922 439686 477978
rect 439742 477922 439838 477978
rect 439218 460350 439838 477922
rect 439218 460294 439314 460350
rect 439370 460294 439438 460350
rect 439494 460294 439562 460350
rect 439618 460294 439686 460350
rect 439742 460294 439838 460350
rect 439218 460226 439838 460294
rect 439218 460170 439314 460226
rect 439370 460170 439438 460226
rect 439494 460170 439562 460226
rect 439618 460170 439686 460226
rect 439742 460170 439838 460226
rect 439218 460102 439838 460170
rect 439218 460046 439314 460102
rect 439370 460046 439438 460102
rect 439494 460046 439562 460102
rect 439618 460046 439686 460102
rect 439742 460046 439838 460102
rect 439218 459978 439838 460046
rect 439218 459922 439314 459978
rect 439370 459922 439438 459978
rect 439494 459922 439562 459978
rect 439618 459922 439686 459978
rect 439742 459922 439838 459978
rect 439218 442350 439838 459922
rect 439218 442294 439314 442350
rect 439370 442294 439438 442350
rect 439494 442294 439562 442350
rect 439618 442294 439686 442350
rect 439742 442294 439838 442350
rect 439218 442226 439838 442294
rect 439218 442170 439314 442226
rect 439370 442170 439438 442226
rect 439494 442170 439562 442226
rect 439618 442170 439686 442226
rect 439742 442170 439838 442226
rect 439218 442102 439838 442170
rect 439218 442046 439314 442102
rect 439370 442046 439438 442102
rect 439494 442046 439562 442102
rect 439618 442046 439686 442102
rect 439742 442046 439838 442102
rect 439218 441978 439838 442046
rect 439218 441922 439314 441978
rect 439370 441922 439438 441978
rect 439494 441922 439562 441978
rect 439618 441922 439686 441978
rect 439742 441922 439838 441978
rect 439218 424350 439838 441922
rect 439218 424294 439314 424350
rect 439370 424294 439438 424350
rect 439494 424294 439562 424350
rect 439618 424294 439686 424350
rect 439742 424294 439838 424350
rect 439218 424226 439838 424294
rect 439218 424170 439314 424226
rect 439370 424170 439438 424226
rect 439494 424170 439562 424226
rect 439618 424170 439686 424226
rect 439742 424170 439838 424226
rect 439218 424102 439838 424170
rect 439218 424046 439314 424102
rect 439370 424046 439438 424102
rect 439494 424046 439562 424102
rect 439618 424046 439686 424102
rect 439742 424046 439838 424102
rect 439218 423978 439838 424046
rect 439218 423922 439314 423978
rect 439370 423922 439438 423978
rect 439494 423922 439562 423978
rect 439618 423922 439686 423978
rect 439742 423922 439838 423978
rect 439218 406350 439838 423922
rect 439218 406294 439314 406350
rect 439370 406294 439438 406350
rect 439494 406294 439562 406350
rect 439618 406294 439686 406350
rect 439742 406294 439838 406350
rect 439218 406226 439838 406294
rect 439218 406170 439314 406226
rect 439370 406170 439438 406226
rect 439494 406170 439562 406226
rect 439618 406170 439686 406226
rect 439742 406170 439838 406226
rect 439218 406102 439838 406170
rect 439218 406046 439314 406102
rect 439370 406046 439438 406102
rect 439494 406046 439562 406102
rect 439618 406046 439686 406102
rect 439742 406046 439838 406102
rect 439218 405978 439838 406046
rect 439218 405922 439314 405978
rect 439370 405922 439438 405978
rect 439494 405922 439562 405978
rect 439618 405922 439686 405978
rect 439742 405922 439838 405978
rect 439218 388350 439838 405922
rect 439218 388294 439314 388350
rect 439370 388294 439438 388350
rect 439494 388294 439562 388350
rect 439618 388294 439686 388350
rect 439742 388294 439838 388350
rect 439218 388226 439838 388294
rect 439218 388170 439314 388226
rect 439370 388170 439438 388226
rect 439494 388170 439562 388226
rect 439618 388170 439686 388226
rect 439742 388170 439838 388226
rect 439218 388102 439838 388170
rect 439218 388046 439314 388102
rect 439370 388046 439438 388102
rect 439494 388046 439562 388102
rect 439618 388046 439686 388102
rect 439742 388046 439838 388102
rect 439218 387978 439838 388046
rect 439218 387922 439314 387978
rect 439370 387922 439438 387978
rect 439494 387922 439562 387978
rect 439618 387922 439686 387978
rect 439742 387922 439838 387978
rect 439218 370350 439838 387922
rect 439218 370294 439314 370350
rect 439370 370294 439438 370350
rect 439494 370294 439562 370350
rect 439618 370294 439686 370350
rect 439742 370294 439838 370350
rect 439218 370226 439838 370294
rect 439218 370170 439314 370226
rect 439370 370170 439438 370226
rect 439494 370170 439562 370226
rect 439618 370170 439686 370226
rect 439742 370170 439838 370226
rect 439218 370102 439838 370170
rect 439218 370046 439314 370102
rect 439370 370046 439438 370102
rect 439494 370046 439562 370102
rect 439618 370046 439686 370102
rect 439742 370046 439838 370102
rect 439218 369978 439838 370046
rect 439218 369922 439314 369978
rect 439370 369922 439438 369978
rect 439494 369922 439562 369978
rect 439618 369922 439686 369978
rect 439742 369922 439838 369978
rect 439218 352350 439838 369922
rect 439218 352294 439314 352350
rect 439370 352294 439438 352350
rect 439494 352294 439562 352350
rect 439618 352294 439686 352350
rect 439742 352294 439838 352350
rect 439218 352226 439838 352294
rect 439218 352170 439314 352226
rect 439370 352170 439438 352226
rect 439494 352170 439562 352226
rect 439618 352170 439686 352226
rect 439742 352170 439838 352226
rect 439218 352102 439838 352170
rect 439218 352046 439314 352102
rect 439370 352046 439438 352102
rect 439494 352046 439562 352102
rect 439618 352046 439686 352102
rect 439742 352046 439838 352102
rect 439218 351978 439838 352046
rect 439218 351922 439314 351978
rect 439370 351922 439438 351978
rect 439494 351922 439562 351978
rect 439618 351922 439686 351978
rect 439742 351922 439838 351978
rect 439218 334350 439838 351922
rect 439218 334294 439314 334350
rect 439370 334294 439438 334350
rect 439494 334294 439562 334350
rect 439618 334294 439686 334350
rect 439742 334294 439838 334350
rect 439218 334226 439838 334294
rect 439218 334170 439314 334226
rect 439370 334170 439438 334226
rect 439494 334170 439562 334226
rect 439618 334170 439686 334226
rect 439742 334170 439838 334226
rect 439218 334102 439838 334170
rect 439218 334046 439314 334102
rect 439370 334046 439438 334102
rect 439494 334046 439562 334102
rect 439618 334046 439686 334102
rect 439742 334046 439838 334102
rect 439218 333978 439838 334046
rect 439218 333922 439314 333978
rect 439370 333922 439438 333978
rect 439494 333922 439562 333978
rect 439618 333922 439686 333978
rect 439742 333922 439838 333978
rect 439218 316350 439838 333922
rect 439218 316294 439314 316350
rect 439370 316294 439438 316350
rect 439494 316294 439562 316350
rect 439618 316294 439686 316350
rect 439742 316294 439838 316350
rect 439218 316226 439838 316294
rect 439218 316170 439314 316226
rect 439370 316170 439438 316226
rect 439494 316170 439562 316226
rect 439618 316170 439686 316226
rect 439742 316170 439838 316226
rect 439218 316102 439838 316170
rect 439218 316046 439314 316102
rect 439370 316046 439438 316102
rect 439494 316046 439562 316102
rect 439618 316046 439686 316102
rect 439742 316046 439838 316102
rect 439218 315978 439838 316046
rect 439218 315922 439314 315978
rect 439370 315922 439438 315978
rect 439494 315922 439562 315978
rect 439618 315922 439686 315978
rect 439742 315922 439838 315978
rect 439218 298350 439838 315922
rect 439218 298294 439314 298350
rect 439370 298294 439438 298350
rect 439494 298294 439562 298350
rect 439618 298294 439686 298350
rect 439742 298294 439838 298350
rect 439218 298226 439838 298294
rect 439218 298170 439314 298226
rect 439370 298170 439438 298226
rect 439494 298170 439562 298226
rect 439618 298170 439686 298226
rect 439742 298170 439838 298226
rect 439218 298102 439838 298170
rect 439218 298046 439314 298102
rect 439370 298046 439438 298102
rect 439494 298046 439562 298102
rect 439618 298046 439686 298102
rect 439742 298046 439838 298102
rect 439218 297978 439838 298046
rect 439218 297922 439314 297978
rect 439370 297922 439438 297978
rect 439494 297922 439562 297978
rect 439618 297922 439686 297978
rect 439742 297922 439838 297978
rect 439218 280350 439838 297922
rect 439218 280294 439314 280350
rect 439370 280294 439438 280350
rect 439494 280294 439562 280350
rect 439618 280294 439686 280350
rect 439742 280294 439838 280350
rect 439218 280226 439838 280294
rect 439218 280170 439314 280226
rect 439370 280170 439438 280226
rect 439494 280170 439562 280226
rect 439618 280170 439686 280226
rect 439742 280170 439838 280226
rect 439218 280102 439838 280170
rect 439218 280046 439314 280102
rect 439370 280046 439438 280102
rect 439494 280046 439562 280102
rect 439618 280046 439686 280102
rect 439742 280046 439838 280102
rect 439218 279978 439838 280046
rect 439218 279922 439314 279978
rect 439370 279922 439438 279978
rect 439494 279922 439562 279978
rect 439618 279922 439686 279978
rect 439742 279922 439838 279978
rect 439218 262350 439838 279922
rect 439218 262294 439314 262350
rect 439370 262294 439438 262350
rect 439494 262294 439562 262350
rect 439618 262294 439686 262350
rect 439742 262294 439838 262350
rect 439218 262226 439838 262294
rect 439218 262170 439314 262226
rect 439370 262170 439438 262226
rect 439494 262170 439562 262226
rect 439618 262170 439686 262226
rect 439742 262170 439838 262226
rect 439218 262102 439838 262170
rect 439218 262046 439314 262102
rect 439370 262046 439438 262102
rect 439494 262046 439562 262102
rect 439618 262046 439686 262102
rect 439742 262046 439838 262102
rect 439218 261978 439838 262046
rect 439218 261922 439314 261978
rect 439370 261922 439438 261978
rect 439494 261922 439562 261978
rect 439618 261922 439686 261978
rect 439742 261922 439838 261978
rect 439218 244350 439838 261922
rect 439218 244294 439314 244350
rect 439370 244294 439438 244350
rect 439494 244294 439562 244350
rect 439618 244294 439686 244350
rect 439742 244294 439838 244350
rect 439218 244226 439838 244294
rect 439218 244170 439314 244226
rect 439370 244170 439438 244226
rect 439494 244170 439562 244226
rect 439618 244170 439686 244226
rect 439742 244170 439838 244226
rect 439218 244102 439838 244170
rect 439218 244046 439314 244102
rect 439370 244046 439438 244102
rect 439494 244046 439562 244102
rect 439618 244046 439686 244102
rect 439742 244046 439838 244102
rect 439218 243978 439838 244046
rect 439218 243922 439314 243978
rect 439370 243922 439438 243978
rect 439494 243922 439562 243978
rect 439618 243922 439686 243978
rect 439742 243922 439838 243978
rect 439218 226350 439838 243922
rect 439218 226294 439314 226350
rect 439370 226294 439438 226350
rect 439494 226294 439562 226350
rect 439618 226294 439686 226350
rect 439742 226294 439838 226350
rect 439218 226226 439838 226294
rect 439218 226170 439314 226226
rect 439370 226170 439438 226226
rect 439494 226170 439562 226226
rect 439618 226170 439686 226226
rect 439742 226170 439838 226226
rect 439218 226102 439838 226170
rect 439218 226046 439314 226102
rect 439370 226046 439438 226102
rect 439494 226046 439562 226102
rect 439618 226046 439686 226102
rect 439742 226046 439838 226102
rect 439218 225978 439838 226046
rect 439218 225922 439314 225978
rect 439370 225922 439438 225978
rect 439494 225922 439562 225978
rect 439618 225922 439686 225978
rect 439742 225922 439838 225978
rect 439218 208350 439838 225922
rect 439218 208294 439314 208350
rect 439370 208294 439438 208350
rect 439494 208294 439562 208350
rect 439618 208294 439686 208350
rect 439742 208294 439838 208350
rect 439218 208226 439838 208294
rect 439218 208170 439314 208226
rect 439370 208170 439438 208226
rect 439494 208170 439562 208226
rect 439618 208170 439686 208226
rect 439742 208170 439838 208226
rect 439218 208102 439838 208170
rect 439218 208046 439314 208102
rect 439370 208046 439438 208102
rect 439494 208046 439562 208102
rect 439618 208046 439686 208102
rect 439742 208046 439838 208102
rect 439218 207978 439838 208046
rect 439218 207922 439314 207978
rect 439370 207922 439438 207978
rect 439494 207922 439562 207978
rect 439618 207922 439686 207978
rect 439742 207922 439838 207978
rect 439218 190350 439838 207922
rect 439218 190294 439314 190350
rect 439370 190294 439438 190350
rect 439494 190294 439562 190350
rect 439618 190294 439686 190350
rect 439742 190294 439838 190350
rect 439218 190226 439838 190294
rect 439218 190170 439314 190226
rect 439370 190170 439438 190226
rect 439494 190170 439562 190226
rect 439618 190170 439686 190226
rect 439742 190170 439838 190226
rect 439218 190102 439838 190170
rect 439218 190046 439314 190102
rect 439370 190046 439438 190102
rect 439494 190046 439562 190102
rect 439618 190046 439686 190102
rect 439742 190046 439838 190102
rect 439218 189978 439838 190046
rect 439218 189922 439314 189978
rect 439370 189922 439438 189978
rect 439494 189922 439562 189978
rect 439618 189922 439686 189978
rect 439742 189922 439838 189978
rect 439218 172350 439838 189922
rect 439218 172294 439314 172350
rect 439370 172294 439438 172350
rect 439494 172294 439562 172350
rect 439618 172294 439686 172350
rect 439742 172294 439838 172350
rect 439218 172226 439838 172294
rect 439218 172170 439314 172226
rect 439370 172170 439438 172226
rect 439494 172170 439562 172226
rect 439618 172170 439686 172226
rect 439742 172170 439838 172226
rect 439218 172102 439838 172170
rect 439218 172046 439314 172102
rect 439370 172046 439438 172102
rect 439494 172046 439562 172102
rect 439618 172046 439686 172102
rect 439742 172046 439838 172102
rect 439218 171978 439838 172046
rect 439218 171922 439314 171978
rect 439370 171922 439438 171978
rect 439494 171922 439562 171978
rect 439618 171922 439686 171978
rect 439742 171922 439838 171978
rect 439218 154350 439838 171922
rect 439218 154294 439314 154350
rect 439370 154294 439438 154350
rect 439494 154294 439562 154350
rect 439618 154294 439686 154350
rect 439742 154294 439838 154350
rect 439218 154226 439838 154294
rect 439218 154170 439314 154226
rect 439370 154170 439438 154226
rect 439494 154170 439562 154226
rect 439618 154170 439686 154226
rect 439742 154170 439838 154226
rect 439218 154102 439838 154170
rect 439218 154046 439314 154102
rect 439370 154046 439438 154102
rect 439494 154046 439562 154102
rect 439618 154046 439686 154102
rect 439742 154046 439838 154102
rect 439218 153978 439838 154046
rect 439218 153922 439314 153978
rect 439370 153922 439438 153978
rect 439494 153922 439562 153978
rect 439618 153922 439686 153978
rect 439742 153922 439838 153978
rect 439218 136350 439838 153922
rect 439218 136294 439314 136350
rect 439370 136294 439438 136350
rect 439494 136294 439562 136350
rect 439618 136294 439686 136350
rect 439742 136294 439838 136350
rect 439218 136226 439838 136294
rect 439218 136170 439314 136226
rect 439370 136170 439438 136226
rect 439494 136170 439562 136226
rect 439618 136170 439686 136226
rect 439742 136170 439838 136226
rect 439218 136102 439838 136170
rect 439218 136046 439314 136102
rect 439370 136046 439438 136102
rect 439494 136046 439562 136102
rect 439618 136046 439686 136102
rect 439742 136046 439838 136102
rect 439218 135978 439838 136046
rect 439218 135922 439314 135978
rect 439370 135922 439438 135978
rect 439494 135922 439562 135978
rect 439618 135922 439686 135978
rect 439742 135922 439838 135978
rect 439218 118350 439838 135922
rect 439218 118294 439314 118350
rect 439370 118294 439438 118350
rect 439494 118294 439562 118350
rect 439618 118294 439686 118350
rect 439742 118294 439838 118350
rect 439218 118226 439838 118294
rect 439218 118170 439314 118226
rect 439370 118170 439438 118226
rect 439494 118170 439562 118226
rect 439618 118170 439686 118226
rect 439742 118170 439838 118226
rect 439218 118102 439838 118170
rect 439218 118046 439314 118102
rect 439370 118046 439438 118102
rect 439494 118046 439562 118102
rect 439618 118046 439686 118102
rect 439742 118046 439838 118102
rect 439218 117978 439838 118046
rect 439218 117922 439314 117978
rect 439370 117922 439438 117978
rect 439494 117922 439562 117978
rect 439618 117922 439686 117978
rect 439742 117922 439838 117978
rect 439218 100350 439838 117922
rect 439218 100294 439314 100350
rect 439370 100294 439438 100350
rect 439494 100294 439562 100350
rect 439618 100294 439686 100350
rect 439742 100294 439838 100350
rect 439218 100226 439838 100294
rect 439218 100170 439314 100226
rect 439370 100170 439438 100226
rect 439494 100170 439562 100226
rect 439618 100170 439686 100226
rect 439742 100170 439838 100226
rect 439218 100102 439838 100170
rect 439218 100046 439314 100102
rect 439370 100046 439438 100102
rect 439494 100046 439562 100102
rect 439618 100046 439686 100102
rect 439742 100046 439838 100102
rect 439218 99978 439838 100046
rect 439218 99922 439314 99978
rect 439370 99922 439438 99978
rect 439494 99922 439562 99978
rect 439618 99922 439686 99978
rect 439742 99922 439838 99978
rect 439218 82350 439838 99922
rect 439218 82294 439314 82350
rect 439370 82294 439438 82350
rect 439494 82294 439562 82350
rect 439618 82294 439686 82350
rect 439742 82294 439838 82350
rect 439218 82226 439838 82294
rect 439218 82170 439314 82226
rect 439370 82170 439438 82226
rect 439494 82170 439562 82226
rect 439618 82170 439686 82226
rect 439742 82170 439838 82226
rect 439218 82102 439838 82170
rect 439218 82046 439314 82102
rect 439370 82046 439438 82102
rect 439494 82046 439562 82102
rect 439618 82046 439686 82102
rect 439742 82046 439838 82102
rect 439218 81978 439838 82046
rect 439218 81922 439314 81978
rect 439370 81922 439438 81978
rect 439494 81922 439562 81978
rect 439618 81922 439686 81978
rect 439742 81922 439838 81978
rect 439218 64350 439838 81922
rect 466218 597212 466838 598268
rect 466218 597156 466314 597212
rect 466370 597156 466438 597212
rect 466494 597156 466562 597212
rect 466618 597156 466686 597212
rect 466742 597156 466838 597212
rect 466218 597088 466838 597156
rect 466218 597032 466314 597088
rect 466370 597032 466438 597088
rect 466494 597032 466562 597088
rect 466618 597032 466686 597088
rect 466742 597032 466838 597088
rect 466218 596964 466838 597032
rect 466218 596908 466314 596964
rect 466370 596908 466438 596964
rect 466494 596908 466562 596964
rect 466618 596908 466686 596964
rect 466742 596908 466838 596964
rect 466218 596840 466838 596908
rect 466218 596784 466314 596840
rect 466370 596784 466438 596840
rect 466494 596784 466562 596840
rect 466618 596784 466686 596840
rect 466742 596784 466838 596840
rect 466218 580350 466838 596784
rect 466218 580294 466314 580350
rect 466370 580294 466438 580350
rect 466494 580294 466562 580350
rect 466618 580294 466686 580350
rect 466742 580294 466838 580350
rect 466218 580226 466838 580294
rect 466218 580170 466314 580226
rect 466370 580170 466438 580226
rect 466494 580170 466562 580226
rect 466618 580170 466686 580226
rect 466742 580170 466838 580226
rect 466218 580102 466838 580170
rect 466218 580046 466314 580102
rect 466370 580046 466438 580102
rect 466494 580046 466562 580102
rect 466618 580046 466686 580102
rect 466742 580046 466838 580102
rect 466218 579978 466838 580046
rect 466218 579922 466314 579978
rect 466370 579922 466438 579978
rect 466494 579922 466562 579978
rect 466618 579922 466686 579978
rect 466742 579922 466838 579978
rect 466218 562350 466838 579922
rect 466218 562294 466314 562350
rect 466370 562294 466438 562350
rect 466494 562294 466562 562350
rect 466618 562294 466686 562350
rect 466742 562294 466838 562350
rect 466218 562226 466838 562294
rect 466218 562170 466314 562226
rect 466370 562170 466438 562226
rect 466494 562170 466562 562226
rect 466618 562170 466686 562226
rect 466742 562170 466838 562226
rect 466218 562102 466838 562170
rect 466218 562046 466314 562102
rect 466370 562046 466438 562102
rect 466494 562046 466562 562102
rect 466618 562046 466686 562102
rect 466742 562046 466838 562102
rect 466218 561978 466838 562046
rect 466218 561922 466314 561978
rect 466370 561922 466438 561978
rect 466494 561922 466562 561978
rect 466618 561922 466686 561978
rect 466742 561922 466838 561978
rect 466218 544350 466838 561922
rect 466218 544294 466314 544350
rect 466370 544294 466438 544350
rect 466494 544294 466562 544350
rect 466618 544294 466686 544350
rect 466742 544294 466838 544350
rect 466218 544226 466838 544294
rect 466218 544170 466314 544226
rect 466370 544170 466438 544226
rect 466494 544170 466562 544226
rect 466618 544170 466686 544226
rect 466742 544170 466838 544226
rect 466218 544102 466838 544170
rect 466218 544046 466314 544102
rect 466370 544046 466438 544102
rect 466494 544046 466562 544102
rect 466618 544046 466686 544102
rect 466742 544046 466838 544102
rect 466218 543978 466838 544046
rect 466218 543922 466314 543978
rect 466370 543922 466438 543978
rect 466494 543922 466562 543978
rect 466618 543922 466686 543978
rect 466742 543922 466838 543978
rect 466218 526350 466838 543922
rect 466218 526294 466314 526350
rect 466370 526294 466438 526350
rect 466494 526294 466562 526350
rect 466618 526294 466686 526350
rect 466742 526294 466838 526350
rect 466218 526226 466838 526294
rect 466218 526170 466314 526226
rect 466370 526170 466438 526226
rect 466494 526170 466562 526226
rect 466618 526170 466686 526226
rect 466742 526170 466838 526226
rect 466218 526102 466838 526170
rect 466218 526046 466314 526102
rect 466370 526046 466438 526102
rect 466494 526046 466562 526102
rect 466618 526046 466686 526102
rect 466742 526046 466838 526102
rect 466218 525978 466838 526046
rect 466218 525922 466314 525978
rect 466370 525922 466438 525978
rect 466494 525922 466562 525978
rect 466618 525922 466686 525978
rect 466742 525922 466838 525978
rect 466218 508350 466838 525922
rect 466218 508294 466314 508350
rect 466370 508294 466438 508350
rect 466494 508294 466562 508350
rect 466618 508294 466686 508350
rect 466742 508294 466838 508350
rect 466218 508226 466838 508294
rect 466218 508170 466314 508226
rect 466370 508170 466438 508226
rect 466494 508170 466562 508226
rect 466618 508170 466686 508226
rect 466742 508170 466838 508226
rect 466218 508102 466838 508170
rect 466218 508046 466314 508102
rect 466370 508046 466438 508102
rect 466494 508046 466562 508102
rect 466618 508046 466686 508102
rect 466742 508046 466838 508102
rect 466218 507978 466838 508046
rect 466218 507922 466314 507978
rect 466370 507922 466438 507978
rect 466494 507922 466562 507978
rect 466618 507922 466686 507978
rect 466742 507922 466838 507978
rect 466218 490350 466838 507922
rect 466218 490294 466314 490350
rect 466370 490294 466438 490350
rect 466494 490294 466562 490350
rect 466618 490294 466686 490350
rect 466742 490294 466838 490350
rect 466218 490226 466838 490294
rect 466218 490170 466314 490226
rect 466370 490170 466438 490226
rect 466494 490170 466562 490226
rect 466618 490170 466686 490226
rect 466742 490170 466838 490226
rect 466218 490102 466838 490170
rect 466218 490046 466314 490102
rect 466370 490046 466438 490102
rect 466494 490046 466562 490102
rect 466618 490046 466686 490102
rect 466742 490046 466838 490102
rect 466218 489978 466838 490046
rect 466218 489922 466314 489978
rect 466370 489922 466438 489978
rect 466494 489922 466562 489978
rect 466618 489922 466686 489978
rect 466742 489922 466838 489978
rect 466218 472350 466838 489922
rect 466218 472294 466314 472350
rect 466370 472294 466438 472350
rect 466494 472294 466562 472350
rect 466618 472294 466686 472350
rect 466742 472294 466838 472350
rect 466218 472226 466838 472294
rect 466218 472170 466314 472226
rect 466370 472170 466438 472226
rect 466494 472170 466562 472226
rect 466618 472170 466686 472226
rect 466742 472170 466838 472226
rect 466218 472102 466838 472170
rect 466218 472046 466314 472102
rect 466370 472046 466438 472102
rect 466494 472046 466562 472102
rect 466618 472046 466686 472102
rect 466742 472046 466838 472102
rect 466218 471978 466838 472046
rect 466218 471922 466314 471978
rect 466370 471922 466438 471978
rect 466494 471922 466562 471978
rect 466618 471922 466686 471978
rect 466742 471922 466838 471978
rect 466218 454350 466838 471922
rect 466218 454294 466314 454350
rect 466370 454294 466438 454350
rect 466494 454294 466562 454350
rect 466618 454294 466686 454350
rect 466742 454294 466838 454350
rect 466218 454226 466838 454294
rect 466218 454170 466314 454226
rect 466370 454170 466438 454226
rect 466494 454170 466562 454226
rect 466618 454170 466686 454226
rect 466742 454170 466838 454226
rect 466218 454102 466838 454170
rect 466218 454046 466314 454102
rect 466370 454046 466438 454102
rect 466494 454046 466562 454102
rect 466618 454046 466686 454102
rect 466742 454046 466838 454102
rect 466218 453978 466838 454046
rect 466218 453922 466314 453978
rect 466370 453922 466438 453978
rect 466494 453922 466562 453978
rect 466618 453922 466686 453978
rect 466742 453922 466838 453978
rect 466218 436350 466838 453922
rect 466218 436294 466314 436350
rect 466370 436294 466438 436350
rect 466494 436294 466562 436350
rect 466618 436294 466686 436350
rect 466742 436294 466838 436350
rect 466218 436226 466838 436294
rect 466218 436170 466314 436226
rect 466370 436170 466438 436226
rect 466494 436170 466562 436226
rect 466618 436170 466686 436226
rect 466742 436170 466838 436226
rect 466218 436102 466838 436170
rect 466218 436046 466314 436102
rect 466370 436046 466438 436102
rect 466494 436046 466562 436102
rect 466618 436046 466686 436102
rect 466742 436046 466838 436102
rect 466218 435978 466838 436046
rect 466218 435922 466314 435978
rect 466370 435922 466438 435978
rect 466494 435922 466562 435978
rect 466618 435922 466686 435978
rect 466742 435922 466838 435978
rect 466218 418350 466838 435922
rect 466218 418294 466314 418350
rect 466370 418294 466438 418350
rect 466494 418294 466562 418350
rect 466618 418294 466686 418350
rect 466742 418294 466838 418350
rect 466218 418226 466838 418294
rect 466218 418170 466314 418226
rect 466370 418170 466438 418226
rect 466494 418170 466562 418226
rect 466618 418170 466686 418226
rect 466742 418170 466838 418226
rect 466218 418102 466838 418170
rect 466218 418046 466314 418102
rect 466370 418046 466438 418102
rect 466494 418046 466562 418102
rect 466618 418046 466686 418102
rect 466742 418046 466838 418102
rect 466218 417978 466838 418046
rect 466218 417922 466314 417978
rect 466370 417922 466438 417978
rect 466494 417922 466562 417978
rect 466618 417922 466686 417978
rect 466742 417922 466838 417978
rect 466218 400350 466838 417922
rect 466218 400294 466314 400350
rect 466370 400294 466438 400350
rect 466494 400294 466562 400350
rect 466618 400294 466686 400350
rect 466742 400294 466838 400350
rect 466218 400226 466838 400294
rect 466218 400170 466314 400226
rect 466370 400170 466438 400226
rect 466494 400170 466562 400226
rect 466618 400170 466686 400226
rect 466742 400170 466838 400226
rect 466218 400102 466838 400170
rect 466218 400046 466314 400102
rect 466370 400046 466438 400102
rect 466494 400046 466562 400102
rect 466618 400046 466686 400102
rect 466742 400046 466838 400102
rect 466218 399978 466838 400046
rect 466218 399922 466314 399978
rect 466370 399922 466438 399978
rect 466494 399922 466562 399978
rect 466618 399922 466686 399978
rect 466742 399922 466838 399978
rect 466218 382350 466838 399922
rect 466218 382294 466314 382350
rect 466370 382294 466438 382350
rect 466494 382294 466562 382350
rect 466618 382294 466686 382350
rect 466742 382294 466838 382350
rect 466218 382226 466838 382294
rect 466218 382170 466314 382226
rect 466370 382170 466438 382226
rect 466494 382170 466562 382226
rect 466618 382170 466686 382226
rect 466742 382170 466838 382226
rect 466218 382102 466838 382170
rect 466218 382046 466314 382102
rect 466370 382046 466438 382102
rect 466494 382046 466562 382102
rect 466618 382046 466686 382102
rect 466742 382046 466838 382102
rect 466218 381978 466838 382046
rect 466218 381922 466314 381978
rect 466370 381922 466438 381978
rect 466494 381922 466562 381978
rect 466618 381922 466686 381978
rect 466742 381922 466838 381978
rect 466218 364350 466838 381922
rect 466218 364294 466314 364350
rect 466370 364294 466438 364350
rect 466494 364294 466562 364350
rect 466618 364294 466686 364350
rect 466742 364294 466838 364350
rect 466218 364226 466838 364294
rect 466218 364170 466314 364226
rect 466370 364170 466438 364226
rect 466494 364170 466562 364226
rect 466618 364170 466686 364226
rect 466742 364170 466838 364226
rect 466218 364102 466838 364170
rect 466218 364046 466314 364102
rect 466370 364046 466438 364102
rect 466494 364046 466562 364102
rect 466618 364046 466686 364102
rect 466742 364046 466838 364102
rect 466218 363978 466838 364046
rect 466218 363922 466314 363978
rect 466370 363922 466438 363978
rect 466494 363922 466562 363978
rect 466618 363922 466686 363978
rect 466742 363922 466838 363978
rect 466218 346350 466838 363922
rect 466218 346294 466314 346350
rect 466370 346294 466438 346350
rect 466494 346294 466562 346350
rect 466618 346294 466686 346350
rect 466742 346294 466838 346350
rect 466218 346226 466838 346294
rect 466218 346170 466314 346226
rect 466370 346170 466438 346226
rect 466494 346170 466562 346226
rect 466618 346170 466686 346226
rect 466742 346170 466838 346226
rect 466218 346102 466838 346170
rect 466218 346046 466314 346102
rect 466370 346046 466438 346102
rect 466494 346046 466562 346102
rect 466618 346046 466686 346102
rect 466742 346046 466838 346102
rect 466218 345978 466838 346046
rect 466218 345922 466314 345978
rect 466370 345922 466438 345978
rect 466494 345922 466562 345978
rect 466618 345922 466686 345978
rect 466742 345922 466838 345978
rect 466218 328350 466838 345922
rect 466218 328294 466314 328350
rect 466370 328294 466438 328350
rect 466494 328294 466562 328350
rect 466618 328294 466686 328350
rect 466742 328294 466838 328350
rect 466218 328226 466838 328294
rect 466218 328170 466314 328226
rect 466370 328170 466438 328226
rect 466494 328170 466562 328226
rect 466618 328170 466686 328226
rect 466742 328170 466838 328226
rect 466218 328102 466838 328170
rect 466218 328046 466314 328102
rect 466370 328046 466438 328102
rect 466494 328046 466562 328102
rect 466618 328046 466686 328102
rect 466742 328046 466838 328102
rect 466218 327978 466838 328046
rect 466218 327922 466314 327978
rect 466370 327922 466438 327978
rect 466494 327922 466562 327978
rect 466618 327922 466686 327978
rect 466742 327922 466838 327978
rect 466218 310350 466838 327922
rect 466218 310294 466314 310350
rect 466370 310294 466438 310350
rect 466494 310294 466562 310350
rect 466618 310294 466686 310350
rect 466742 310294 466838 310350
rect 466218 310226 466838 310294
rect 466218 310170 466314 310226
rect 466370 310170 466438 310226
rect 466494 310170 466562 310226
rect 466618 310170 466686 310226
rect 466742 310170 466838 310226
rect 466218 310102 466838 310170
rect 466218 310046 466314 310102
rect 466370 310046 466438 310102
rect 466494 310046 466562 310102
rect 466618 310046 466686 310102
rect 466742 310046 466838 310102
rect 466218 309978 466838 310046
rect 466218 309922 466314 309978
rect 466370 309922 466438 309978
rect 466494 309922 466562 309978
rect 466618 309922 466686 309978
rect 466742 309922 466838 309978
rect 466218 292350 466838 309922
rect 466218 292294 466314 292350
rect 466370 292294 466438 292350
rect 466494 292294 466562 292350
rect 466618 292294 466686 292350
rect 466742 292294 466838 292350
rect 466218 292226 466838 292294
rect 466218 292170 466314 292226
rect 466370 292170 466438 292226
rect 466494 292170 466562 292226
rect 466618 292170 466686 292226
rect 466742 292170 466838 292226
rect 466218 292102 466838 292170
rect 466218 292046 466314 292102
rect 466370 292046 466438 292102
rect 466494 292046 466562 292102
rect 466618 292046 466686 292102
rect 466742 292046 466838 292102
rect 466218 291978 466838 292046
rect 466218 291922 466314 291978
rect 466370 291922 466438 291978
rect 466494 291922 466562 291978
rect 466618 291922 466686 291978
rect 466742 291922 466838 291978
rect 466218 274350 466838 291922
rect 466218 274294 466314 274350
rect 466370 274294 466438 274350
rect 466494 274294 466562 274350
rect 466618 274294 466686 274350
rect 466742 274294 466838 274350
rect 466218 274226 466838 274294
rect 466218 274170 466314 274226
rect 466370 274170 466438 274226
rect 466494 274170 466562 274226
rect 466618 274170 466686 274226
rect 466742 274170 466838 274226
rect 466218 274102 466838 274170
rect 466218 274046 466314 274102
rect 466370 274046 466438 274102
rect 466494 274046 466562 274102
rect 466618 274046 466686 274102
rect 466742 274046 466838 274102
rect 466218 273978 466838 274046
rect 466218 273922 466314 273978
rect 466370 273922 466438 273978
rect 466494 273922 466562 273978
rect 466618 273922 466686 273978
rect 466742 273922 466838 273978
rect 466218 256350 466838 273922
rect 466218 256294 466314 256350
rect 466370 256294 466438 256350
rect 466494 256294 466562 256350
rect 466618 256294 466686 256350
rect 466742 256294 466838 256350
rect 466218 256226 466838 256294
rect 466218 256170 466314 256226
rect 466370 256170 466438 256226
rect 466494 256170 466562 256226
rect 466618 256170 466686 256226
rect 466742 256170 466838 256226
rect 466218 256102 466838 256170
rect 466218 256046 466314 256102
rect 466370 256046 466438 256102
rect 466494 256046 466562 256102
rect 466618 256046 466686 256102
rect 466742 256046 466838 256102
rect 466218 255978 466838 256046
rect 466218 255922 466314 255978
rect 466370 255922 466438 255978
rect 466494 255922 466562 255978
rect 466618 255922 466686 255978
rect 466742 255922 466838 255978
rect 466218 238350 466838 255922
rect 466218 238294 466314 238350
rect 466370 238294 466438 238350
rect 466494 238294 466562 238350
rect 466618 238294 466686 238350
rect 466742 238294 466838 238350
rect 466218 238226 466838 238294
rect 466218 238170 466314 238226
rect 466370 238170 466438 238226
rect 466494 238170 466562 238226
rect 466618 238170 466686 238226
rect 466742 238170 466838 238226
rect 466218 238102 466838 238170
rect 466218 238046 466314 238102
rect 466370 238046 466438 238102
rect 466494 238046 466562 238102
rect 466618 238046 466686 238102
rect 466742 238046 466838 238102
rect 466218 237978 466838 238046
rect 466218 237922 466314 237978
rect 466370 237922 466438 237978
rect 466494 237922 466562 237978
rect 466618 237922 466686 237978
rect 466742 237922 466838 237978
rect 466218 220350 466838 237922
rect 466218 220294 466314 220350
rect 466370 220294 466438 220350
rect 466494 220294 466562 220350
rect 466618 220294 466686 220350
rect 466742 220294 466838 220350
rect 466218 220226 466838 220294
rect 466218 220170 466314 220226
rect 466370 220170 466438 220226
rect 466494 220170 466562 220226
rect 466618 220170 466686 220226
rect 466742 220170 466838 220226
rect 466218 220102 466838 220170
rect 466218 220046 466314 220102
rect 466370 220046 466438 220102
rect 466494 220046 466562 220102
rect 466618 220046 466686 220102
rect 466742 220046 466838 220102
rect 466218 219978 466838 220046
rect 466218 219922 466314 219978
rect 466370 219922 466438 219978
rect 466494 219922 466562 219978
rect 466618 219922 466686 219978
rect 466742 219922 466838 219978
rect 466218 202350 466838 219922
rect 466218 202294 466314 202350
rect 466370 202294 466438 202350
rect 466494 202294 466562 202350
rect 466618 202294 466686 202350
rect 466742 202294 466838 202350
rect 466218 202226 466838 202294
rect 466218 202170 466314 202226
rect 466370 202170 466438 202226
rect 466494 202170 466562 202226
rect 466618 202170 466686 202226
rect 466742 202170 466838 202226
rect 466218 202102 466838 202170
rect 466218 202046 466314 202102
rect 466370 202046 466438 202102
rect 466494 202046 466562 202102
rect 466618 202046 466686 202102
rect 466742 202046 466838 202102
rect 466218 201978 466838 202046
rect 466218 201922 466314 201978
rect 466370 201922 466438 201978
rect 466494 201922 466562 201978
rect 466618 201922 466686 201978
rect 466742 201922 466838 201978
rect 466218 184350 466838 201922
rect 466218 184294 466314 184350
rect 466370 184294 466438 184350
rect 466494 184294 466562 184350
rect 466618 184294 466686 184350
rect 466742 184294 466838 184350
rect 466218 184226 466838 184294
rect 466218 184170 466314 184226
rect 466370 184170 466438 184226
rect 466494 184170 466562 184226
rect 466618 184170 466686 184226
rect 466742 184170 466838 184226
rect 466218 184102 466838 184170
rect 466218 184046 466314 184102
rect 466370 184046 466438 184102
rect 466494 184046 466562 184102
rect 466618 184046 466686 184102
rect 466742 184046 466838 184102
rect 466218 183978 466838 184046
rect 466218 183922 466314 183978
rect 466370 183922 466438 183978
rect 466494 183922 466562 183978
rect 466618 183922 466686 183978
rect 466742 183922 466838 183978
rect 466218 166350 466838 183922
rect 466218 166294 466314 166350
rect 466370 166294 466438 166350
rect 466494 166294 466562 166350
rect 466618 166294 466686 166350
rect 466742 166294 466838 166350
rect 466218 166226 466838 166294
rect 466218 166170 466314 166226
rect 466370 166170 466438 166226
rect 466494 166170 466562 166226
rect 466618 166170 466686 166226
rect 466742 166170 466838 166226
rect 466218 166102 466838 166170
rect 466218 166046 466314 166102
rect 466370 166046 466438 166102
rect 466494 166046 466562 166102
rect 466618 166046 466686 166102
rect 466742 166046 466838 166102
rect 466218 165978 466838 166046
rect 466218 165922 466314 165978
rect 466370 165922 466438 165978
rect 466494 165922 466562 165978
rect 466618 165922 466686 165978
rect 466742 165922 466838 165978
rect 466218 148350 466838 165922
rect 466218 148294 466314 148350
rect 466370 148294 466438 148350
rect 466494 148294 466562 148350
rect 466618 148294 466686 148350
rect 466742 148294 466838 148350
rect 466218 148226 466838 148294
rect 466218 148170 466314 148226
rect 466370 148170 466438 148226
rect 466494 148170 466562 148226
rect 466618 148170 466686 148226
rect 466742 148170 466838 148226
rect 466218 148102 466838 148170
rect 466218 148046 466314 148102
rect 466370 148046 466438 148102
rect 466494 148046 466562 148102
rect 466618 148046 466686 148102
rect 466742 148046 466838 148102
rect 466218 147978 466838 148046
rect 466218 147922 466314 147978
rect 466370 147922 466438 147978
rect 466494 147922 466562 147978
rect 466618 147922 466686 147978
rect 466742 147922 466838 147978
rect 466218 130350 466838 147922
rect 466218 130294 466314 130350
rect 466370 130294 466438 130350
rect 466494 130294 466562 130350
rect 466618 130294 466686 130350
rect 466742 130294 466838 130350
rect 466218 130226 466838 130294
rect 466218 130170 466314 130226
rect 466370 130170 466438 130226
rect 466494 130170 466562 130226
rect 466618 130170 466686 130226
rect 466742 130170 466838 130226
rect 466218 130102 466838 130170
rect 466218 130046 466314 130102
rect 466370 130046 466438 130102
rect 466494 130046 466562 130102
rect 466618 130046 466686 130102
rect 466742 130046 466838 130102
rect 466218 129978 466838 130046
rect 466218 129922 466314 129978
rect 466370 129922 466438 129978
rect 466494 129922 466562 129978
rect 466618 129922 466686 129978
rect 466742 129922 466838 129978
rect 466218 112350 466838 129922
rect 466218 112294 466314 112350
rect 466370 112294 466438 112350
rect 466494 112294 466562 112350
rect 466618 112294 466686 112350
rect 466742 112294 466838 112350
rect 466218 112226 466838 112294
rect 466218 112170 466314 112226
rect 466370 112170 466438 112226
rect 466494 112170 466562 112226
rect 466618 112170 466686 112226
rect 466742 112170 466838 112226
rect 466218 112102 466838 112170
rect 466218 112046 466314 112102
rect 466370 112046 466438 112102
rect 466494 112046 466562 112102
rect 466618 112046 466686 112102
rect 466742 112046 466838 112102
rect 466218 111978 466838 112046
rect 466218 111922 466314 111978
rect 466370 111922 466438 111978
rect 466494 111922 466562 111978
rect 466618 111922 466686 111978
rect 466742 111922 466838 111978
rect 466218 94350 466838 111922
rect 466218 94294 466314 94350
rect 466370 94294 466438 94350
rect 466494 94294 466562 94350
rect 466618 94294 466686 94350
rect 466742 94294 466838 94350
rect 466218 94226 466838 94294
rect 466218 94170 466314 94226
rect 466370 94170 466438 94226
rect 466494 94170 466562 94226
rect 466618 94170 466686 94226
rect 466742 94170 466838 94226
rect 466218 94102 466838 94170
rect 466218 94046 466314 94102
rect 466370 94046 466438 94102
rect 466494 94046 466562 94102
rect 466618 94046 466686 94102
rect 466742 94046 466838 94102
rect 466218 93978 466838 94046
rect 466218 93922 466314 93978
rect 466370 93922 466438 93978
rect 466494 93922 466562 93978
rect 466618 93922 466686 93978
rect 466742 93922 466838 93978
rect 439218 64294 439314 64350
rect 439370 64294 439438 64350
rect 439494 64294 439562 64350
rect 439618 64294 439686 64350
rect 439742 64294 439838 64350
rect 439218 64226 439838 64294
rect 439218 64170 439314 64226
rect 439370 64170 439438 64226
rect 439494 64170 439562 64226
rect 439618 64170 439686 64226
rect 439742 64170 439838 64226
rect 439218 64102 439838 64170
rect 439218 64046 439314 64102
rect 439370 64046 439438 64102
rect 439494 64046 439562 64102
rect 439618 64046 439686 64102
rect 439742 64046 439838 64102
rect 439218 63978 439838 64046
rect 439218 63922 439314 63978
rect 439370 63922 439438 63978
rect 439494 63922 439562 63978
rect 439618 63922 439686 63978
rect 439742 63922 439838 63978
rect 435498 40294 435594 40350
rect 435650 40294 435718 40350
rect 435774 40294 435842 40350
rect 435898 40294 435966 40350
rect 436022 40294 436118 40350
rect 435498 40226 436118 40294
rect 435498 40170 435594 40226
rect 435650 40170 435718 40226
rect 435774 40170 435842 40226
rect 435898 40170 435966 40226
rect 436022 40170 436118 40226
rect 435498 40102 436118 40170
rect 435498 40046 435594 40102
rect 435650 40046 435718 40102
rect 435774 40046 435842 40102
rect 435898 40046 435966 40102
rect 436022 40046 436118 40102
rect 435498 39978 436118 40046
rect 435498 39922 435594 39978
rect 435650 39922 435718 39978
rect 435774 39922 435842 39978
rect 435898 39922 435966 39978
rect 436022 39922 436118 39978
rect 435498 22350 436118 39922
rect 435498 22294 435594 22350
rect 435650 22294 435718 22350
rect 435774 22294 435842 22350
rect 435898 22294 435966 22350
rect 436022 22294 436118 22350
rect 435498 22226 436118 22294
rect 435498 22170 435594 22226
rect 435650 22170 435718 22226
rect 435774 22170 435842 22226
rect 435898 22170 435966 22226
rect 436022 22170 436118 22226
rect 435498 22102 436118 22170
rect 435498 22046 435594 22102
rect 435650 22046 435718 22102
rect 435774 22046 435842 22102
rect 435898 22046 435966 22102
rect 436022 22046 436118 22102
rect 435498 21978 436118 22046
rect 435498 21922 435594 21978
rect 435650 21922 435718 21978
rect 435774 21922 435842 21978
rect 435898 21922 435966 21978
rect 436022 21922 436118 21978
rect 435498 4350 436118 21922
rect 435498 4294 435594 4350
rect 435650 4294 435718 4350
rect 435774 4294 435842 4350
rect 435898 4294 435966 4350
rect 436022 4294 436118 4350
rect 435498 4226 436118 4294
rect 435498 4170 435594 4226
rect 435650 4170 435718 4226
rect 435774 4170 435842 4226
rect 435898 4170 435966 4226
rect 436022 4170 436118 4226
rect 414988 3378 415044 3388
rect 435498 4102 436118 4170
rect 436828 51058 436884 51068
rect 436828 4228 436884 51002
rect 439218 46350 439838 63922
rect 446908 79318 446964 79328
rect 439218 46294 439314 46350
rect 439370 46294 439438 46350
rect 439494 46294 439562 46350
rect 439618 46294 439686 46350
rect 439742 46294 439838 46350
rect 439218 46226 439838 46294
rect 439218 46170 439314 46226
rect 439370 46170 439438 46226
rect 439494 46170 439562 46226
rect 439618 46170 439686 46226
rect 439742 46170 439838 46226
rect 439218 46102 439838 46170
rect 439218 46046 439314 46102
rect 439370 46046 439438 46102
rect 439494 46046 439562 46102
rect 439618 46046 439686 46102
rect 439742 46046 439838 46102
rect 439218 45978 439838 46046
rect 439218 45922 439314 45978
rect 439370 45922 439438 45978
rect 439494 45922 439562 45978
rect 439618 45922 439686 45978
rect 439742 45922 439838 45978
rect 439218 28350 439838 45922
rect 439218 28294 439314 28350
rect 439370 28294 439438 28350
rect 439494 28294 439562 28350
rect 439618 28294 439686 28350
rect 439742 28294 439838 28350
rect 439218 28226 439838 28294
rect 439218 28170 439314 28226
rect 439370 28170 439438 28226
rect 439494 28170 439562 28226
rect 439618 28170 439686 28226
rect 439742 28170 439838 28226
rect 439218 28102 439838 28170
rect 439218 28046 439314 28102
rect 439370 28046 439438 28102
rect 439494 28046 439562 28102
rect 439618 28046 439686 28102
rect 439742 28046 439838 28102
rect 439218 27978 439838 28046
rect 439218 27922 439314 27978
rect 439370 27922 439438 27978
rect 439494 27922 439562 27978
rect 439618 27922 439686 27978
rect 439742 27922 439838 27978
rect 436828 4162 436884 4172
rect 438508 11998 438564 12008
rect 438508 4228 438564 11942
rect 438508 4162 438564 4172
rect 439218 10350 439838 27922
rect 439218 10294 439314 10350
rect 439370 10294 439438 10350
rect 439494 10294 439562 10350
rect 439618 10294 439686 10350
rect 439742 10294 439838 10350
rect 439218 10226 439838 10294
rect 439218 10170 439314 10226
rect 439370 10170 439438 10226
rect 439494 10170 439562 10226
rect 439618 10170 439686 10226
rect 439742 10170 439838 10226
rect 439218 10102 439838 10170
rect 439218 10046 439314 10102
rect 439370 10046 439438 10102
rect 439494 10046 439562 10102
rect 439618 10046 439686 10102
rect 439742 10046 439838 10102
rect 439218 9978 439838 10046
rect 439218 9922 439314 9978
rect 439370 9922 439438 9978
rect 439494 9922 439562 9978
rect 439618 9922 439686 9978
rect 439742 9922 439838 9978
rect 435498 4046 435594 4102
rect 435650 4046 435718 4102
rect 435774 4046 435842 4102
rect 435898 4046 435966 4102
rect 436022 4046 436118 4102
rect 435498 3978 436118 4046
rect 435498 3922 435594 3978
rect 435650 3922 435718 3978
rect 435774 3922 435842 3978
rect 435898 3922 435966 3978
rect 436022 3922 436118 3978
rect 408498 -1176 408594 -1120
rect 408650 -1176 408718 -1120
rect 408774 -1176 408842 -1120
rect 408898 -1176 408966 -1120
rect 409022 -1176 409118 -1120
rect 408498 -1244 409118 -1176
rect 408498 -1300 408594 -1244
rect 408650 -1300 408718 -1244
rect 408774 -1300 408842 -1244
rect 408898 -1300 408966 -1244
rect 409022 -1300 409118 -1244
rect 408498 -1368 409118 -1300
rect 408498 -1424 408594 -1368
rect 408650 -1424 408718 -1368
rect 408774 -1424 408842 -1368
rect 408898 -1424 408966 -1368
rect 409022 -1424 409118 -1368
rect 408498 -1492 409118 -1424
rect 408498 -1548 408594 -1492
rect 408650 -1548 408718 -1492
rect 408774 -1548 408842 -1492
rect 408898 -1548 408966 -1492
rect 409022 -1548 409118 -1492
rect 408498 -1644 409118 -1548
rect 435498 -160 436118 3922
rect 435498 -216 435594 -160
rect 435650 -216 435718 -160
rect 435774 -216 435842 -160
rect 435898 -216 435966 -160
rect 436022 -216 436118 -160
rect 435498 -284 436118 -216
rect 435498 -340 435594 -284
rect 435650 -340 435718 -284
rect 435774 -340 435842 -284
rect 435898 -340 435966 -284
rect 436022 -340 436118 -284
rect 435498 -408 436118 -340
rect 435498 -464 435594 -408
rect 435650 -464 435718 -408
rect 435774 -464 435842 -408
rect 435898 -464 435966 -408
rect 436022 -464 436118 -408
rect 435498 -532 436118 -464
rect 435498 -588 435594 -532
rect 435650 -588 435718 -532
rect 435774 -588 435842 -532
rect 435898 -588 435966 -532
rect 436022 -588 436118 -532
rect 435498 -1644 436118 -588
rect 439218 -1120 439838 9922
rect 443548 49078 443604 49088
rect 443548 4228 443604 49022
rect 443548 4162 443604 4172
rect 446908 4228 446964 79262
rect 466218 76350 466838 93922
rect 466218 76294 466314 76350
rect 466370 76294 466438 76350
rect 466494 76294 466562 76350
rect 466618 76294 466686 76350
rect 466742 76294 466838 76350
rect 466218 76226 466838 76294
rect 466218 76170 466314 76226
rect 466370 76170 466438 76226
rect 466494 76170 466562 76226
rect 466618 76170 466686 76226
rect 466742 76170 466838 76226
rect 466218 76102 466838 76170
rect 466218 76046 466314 76102
rect 466370 76046 466438 76102
rect 466494 76046 466562 76102
rect 466618 76046 466686 76102
rect 466742 76046 466838 76102
rect 466218 75978 466838 76046
rect 466218 75922 466314 75978
rect 466370 75922 466438 75978
rect 466494 75922 466562 75978
rect 466618 75922 466686 75978
rect 466742 75922 466838 75978
rect 451948 74098 452004 74108
rect 446908 4162 446964 4172
rect 448588 47458 448644 47468
rect 448588 4228 448644 47402
rect 448588 4162 448644 4172
rect 450268 22618 450324 22628
rect 450268 4228 450324 22562
rect 450268 4162 450324 4172
rect 451948 4228 452004 74042
rect 458668 59338 458724 59348
rect 451948 4162 452004 4172
rect 453628 54478 453684 54488
rect 453628 4228 453684 54422
rect 458668 20188 458724 59282
rect 466218 58350 466838 75922
rect 469938 598172 470558 598268
rect 469938 598116 470034 598172
rect 470090 598116 470158 598172
rect 470214 598116 470282 598172
rect 470338 598116 470406 598172
rect 470462 598116 470558 598172
rect 469938 598048 470558 598116
rect 469938 597992 470034 598048
rect 470090 597992 470158 598048
rect 470214 597992 470282 598048
rect 470338 597992 470406 598048
rect 470462 597992 470558 598048
rect 469938 597924 470558 597992
rect 469938 597868 470034 597924
rect 470090 597868 470158 597924
rect 470214 597868 470282 597924
rect 470338 597868 470406 597924
rect 470462 597868 470558 597924
rect 469938 597800 470558 597868
rect 469938 597744 470034 597800
rect 470090 597744 470158 597800
rect 470214 597744 470282 597800
rect 470338 597744 470406 597800
rect 470462 597744 470558 597800
rect 469938 586350 470558 597744
rect 469938 586294 470034 586350
rect 470090 586294 470158 586350
rect 470214 586294 470282 586350
rect 470338 586294 470406 586350
rect 470462 586294 470558 586350
rect 469938 586226 470558 586294
rect 469938 586170 470034 586226
rect 470090 586170 470158 586226
rect 470214 586170 470282 586226
rect 470338 586170 470406 586226
rect 470462 586170 470558 586226
rect 469938 586102 470558 586170
rect 469938 586046 470034 586102
rect 470090 586046 470158 586102
rect 470214 586046 470282 586102
rect 470338 586046 470406 586102
rect 470462 586046 470558 586102
rect 469938 585978 470558 586046
rect 469938 585922 470034 585978
rect 470090 585922 470158 585978
rect 470214 585922 470282 585978
rect 470338 585922 470406 585978
rect 470462 585922 470558 585978
rect 469938 568350 470558 585922
rect 469938 568294 470034 568350
rect 470090 568294 470158 568350
rect 470214 568294 470282 568350
rect 470338 568294 470406 568350
rect 470462 568294 470558 568350
rect 469938 568226 470558 568294
rect 469938 568170 470034 568226
rect 470090 568170 470158 568226
rect 470214 568170 470282 568226
rect 470338 568170 470406 568226
rect 470462 568170 470558 568226
rect 469938 568102 470558 568170
rect 469938 568046 470034 568102
rect 470090 568046 470158 568102
rect 470214 568046 470282 568102
rect 470338 568046 470406 568102
rect 470462 568046 470558 568102
rect 469938 567978 470558 568046
rect 469938 567922 470034 567978
rect 470090 567922 470158 567978
rect 470214 567922 470282 567978
rect 470338 567922 470406 567978
rect 470462 567922 470558 567978
rect 469938 550350 470558 567922
rect 469938 550294 470034 550350
rect 470090 550294 470158 550350
rect 470214 550294 470282 550350
rect 470338 550294 470406 550350
rect 470462 550294 470558 550350
rect 469938 550226 470558 550294
rect 469938 550170 470034 550226
rect 470090 550170 470158 550226
rect 470214 550170 470282 550226
rect 470338 550170 470406 550226
rect 470462 550170 470558 550226
rect 469938 550102 470558 550170
rect 469938 550046 470034 550102
rect 470090 550046 470158 550102
rect 470214 550046 470282 550102
rect 470338 550046 470406 550102
rect 470462 550046 470558 550102
rect 469938 549978 470558 550046
rect 469938 549922 470034 549978
rect 470090 549922 470158 549978
rect 470214 549922 470282 549978
rect 470338 549922 470406 549978
rect 470462 549922 470558 549978
rect 469938 532350 470558 549922
rect 469938 532294 470034 532350
rect 470090 532294 470158 532350
rect 470214 532294 470282 532350
rect 470338 532294 470406 532350
rect 470462 532294 470558 532350
rect 469938 532226 470558 532294
rect 469938 532170 470034 532226
rect 470090 532170 470158 532226
rect 470214 532170 470282 532226
rect 470338 532170 470406 532226
rect 470462 532170 470558 532226
rect 469938 532102 470558 532170
rect 469938 532046 470034 532102
rect 470090 532046 470158 532102
rect 470214 532046 470282 532102
rect 470338 532046 470406 532102
rect 470462 532046 470558 532102
rect 469938 531978 470558 532046
rect 469938 531922 470034 531978
rect 470090 531922 470158 531978
rect 470214 531922 470282 531978
rect 470338 531922 470406 531978
rect 470462 531922 470558 531978
rect 469938 514350 470558 531922
rect 469938 514294 470034 514350
rect 470090 514294 470158 514350
rect 470214 514294 470282 514350
rect 470338 514294 470406 514350
rect 470462 514294 470558 514350
rect 469938 514226 470558 514294
rect 469938 514170 470034 514226
rect 470090 514170 470158 514226
rect 470214 514170 470282 514226
rect 470338 514170 470406 514226
rect 470462 514170 470558 514226
rect 469938 514102 470558 514170
rect 469938 514046 470034 514102
rect 470090 514046 470158 514102
rect 470214 514046 470282 514102
rect 470338 514046 470406 514102
rect 470462 514046 470558 514102
rect 469938 513978 470558 514046
rect 469938 513922 470034 513978
rect 470090 513922 470158 513978
rect 470214 513922 470282 513978
rect 470338 513922 470406 513978
rect 470462 513922 470558 513978
rect 469938 496350 470558 513922
rect 469938 496294 470034 496350
rect 470090 496294 470158 496350
rect 470214 496294 470282 496350
rect 470338 496294 470406 496350
rect 470462 496294 470558 496350
rect 469938 496226 470558 496294
rect 469938 496170 470034 496226
rect 470090 496170 470158 496226
rect 470214 496170 470282 496226
rect 470338 496170 470406 496226
rect 470462 496170 470558 496226
rect 469938 496102 470558 496170
rect 469938 496046 470034 496102
rect 470090 496046 470158 496102
rect 470214 496046 470282 496102
rect 470338 496046 470406 496102
rect 470462 496046 470558 496102
rect 469938 495978 470558 496046
rect 469938 495922 470034 495978
rect 470090 495922 470158 495978
rect 470214 495922 470282 495978
rect 470338 495922 470406 495978
rect 470462 495922 470558 495978
rect 469938 478350 470558 495922
rect 469938 478294 470034 478350
rect 470090 478294 470158 478350
rect 470214 478294 470282 478350
rect 470338 478294 470406 478350
rect 470462 478294 470558 478350
rect 469938 478226 470558 478294
rect 469938 478170 470034 478226
rect 470090 478170 470158 478226
rect 470214 478170 470282 478226
rect 470338 478170 470406 478226
rect 470462 478170 470558 478226
rect 469938 478102 470558 478170
rect 469938 478046 470034 478102
rect 470090 478046 470158 478102
rect 470214 478046 470282 478102
rect 470338 478046 470406 478102
rect 470462 478046 470558 478102
rect 469938 477978 470558 478046
rect 469938 477922 470034 477978
rect 470090 477922 470158 477978
rect 470214 477922 470282 477978
rect 470338 477922 470406 477978
rect 470462 477922 470558 477978
rect 469938 460350 470558 477922
rect 469938 460294 470034 460350
rect 470090 460294 470158 460350
rect 470214 460294 470282 460350
rect 470338 460294 470406 460350
rect 470462 460294 470558 460350
rect 469938 460226 470558 460294
rect 469938 460170 470034 460226
rect 470090 460170 470158 460226
rect 470214 460170 470282 460226
rect 470338 460170 470406 460226
rect 470462 460170 470558 460226
rect 469938 460102 470558 460170
rect 469938 460046 470034 460102
rect 470090 460046 470158 460102
rect 470214 460046 470282 460102
rect 470338 460046 470406 460102
rect 470462 460046 470558 460102
rect 469938 459978 470558 460046
rect 469938 459922 470034 459978
rect 470090 459922 470158 459978
rect 470214 459922 470282 459978
rect 470338 459922 470406 459978
rect 470462 459922 470558 459978
rect 469938 442350 470558 459922
rect 469938 442294 470034 442350
rect 470090 442294 470158 442350
rect 470214 442294 470282 442350
rect 470338 442294 470406 442350
rect 470462 442294 470558 442350
rect 469938 442226 470558 442294
rect 469938 442170 470034 442226
rect 470090 442170 470158 442226
rect 470214 442170 470282 442226
rect 470338 442170 470406 442226
rect 470462 442170 470558 442226
rect 469938 442102 470558 442170
rect 469938 442046 470034 442102
rect 470090 442046 470158 442102
rect 470214 442046 470282 442102
rect 470338 442046 470406 442102
rect 470462 442046 470558 442102
rect 469938 441978 470558 442046
rect 469938 441922 470034 441978
rect 470090 441922 470158 441978
rect 470214 441922 470282 441978
rect 470338 441922 470406 441978
rect 470462 441922 470558 441978
rect 469938 424350 470558 441922
rect 469938 424294 470034 424350
rect 470090 424294 470158 424350
rect 470214 424294 470282 424350
rect 470338 424294 470406 424350
rect 470462 424294 470558 424350
rect 469938 424226 470558 424294
rect 469938 424170 470034 424226
rect 470090 424170 470158 424226
rect 470214 424170 470282 424226
rect 470338 424170 470406 424226
rect 470462 424170 470558 424226
rect 469938 424102 470558 424170
rect 469938 424046 470034 424102
rect 470090 424046 470158 424102
rect 470214 424046 470282 424102
rect 470338 424046 470406 424102
rect 470462 424046 470558 424102
rect 469938 423978 470558 424046
rect 469938 423922 470034 423978
rect 470090 423922 470158 423978
rect 470214 423922 470282 423978
rect 470338 423922 470406 423978
rect 470462 423922 470558 423978
rect 469938 406350 470558 423922
rect 469938 406294 470034 406350
rect 470090 406294 470158 406350
rect 470214 406294 470282 406350
rect 470338 406294 470406 406350
rect 470462 406294 470558 406350
rect 469938 406226 470558 406294
rect 469938 406170 470034 406226
rect 470090 406170 470158 406226
rect 470214 406170 470282 406226
rect 470338 406170 470406 406226
rect 470462 406170 470558 406226
rect 469938 406102 470558 406170
rect 469938 406046 470034 406102
rect 470090 406046 470158 406102
rect 470214 406046 470282 406102
rect 470338 406046 470406 406102
rect 470462 406046 470558 406102
rect 469938 405978 470558 406046
rect 469938 405922 470034 405978
rect 470090 405922 470158 405978
rect 470214 405922 470282 405978
rect 470338 405922 470406 405978
rect 470462 405922 470558 405978
rect 469938 388350 470558 405922
rect 469938 388294 470034 388350
rect 470090 388294 470158 388350
rect 470214 388294 470282 388350
rect 470338 388294 470406 388350
rect 470462 388294 470558 388350
rect 469938 388226 470558 388294
rect 469938 388170 470034 388226
rect 470090 388170 470158 388226
rect 470214 388170 470282 388226
rect 470338 388170 470406 388226
rect 470462 388170 470558 388226
rect 469938 388102 470558 388170
rect 469938 388046 470034 388102
rect 470090 388046 470158 388102
rect 470214 388046 470282 388102
rect 470338 388046 470406 388102
rect 470462 388046 470558 388102
rect 469938 387978 470558 388046
rect 469938 387922 470034 387978
rect 470090 387922 470158 387978
rect 470214 387922 470282 387978
rect 470338 387922 470406 387978
rect 470462 387922 470558 387978
rect 469938 370350 470558 387922
rect 469938 370294 470034 370350
rect 470090 370294 470158 370350
rect 470214 370294 470282 370350
rect 470338 370294 470406 370350
rect 470462 370294 470558 370350
rect 469938 370226 470558 370294
rect 469938 370170 470034 370226
rect 470090 370170 470158 370226
rect 470214 370170 470282 370226
rect 470338 370170 470406 370226
rect 470462 370170 470558 370226
rect 469938 370102 470558 370170
rect 469938 370046 470034 370102
rect 470090 370046 470158 370102
rect 470214 370046 470282 370102
rect 470338 370046 470406 370102
rect 470462 370046 470558 370102
rect 469938 369978 470558 370046
rect 469938 369922 470034 369978
rect 470090 369922 470158 369978
rect 470214 369922 470282 369978
rect 470338 369922 470406 369978
rect 470462 369922 470558 369978
rect 469938 352350 470558 369922
rect 469938 352294 470034 352350
rect 470090 352294 470158 352350
rect 470214 352294 470282 352350
rect 470338 352294 470406 352350
rect 470462 352294 470558 352350
rect 469938 352226 470558 352294
rect 469938 352170 470034 352226
rect 470090 352170 470158 352226
rect 470214 352170 470282 352226
rect 470338 352170 470406 352226
rect 470462 352170 470558 352226
rect 469938 352102 470558 352170
rect 469938 352046 470034 352102
rect 470090 352046 470158 352102
rect 470214 352046 470282 352102
rect 470338 352046 470406 352102
rect 470462 352046 470558 352102
rect 469938 351978 470558 352046
rect 469938 351922 470034 351978
rect 470090 351922 470158 351978
rect 470214 351922 470282 351978
rect 470338 351922 470406 351978
rect 470462 351922 470558 351978
rect 469938 334350 470558 351922
rect 469938 334294 470034 334350
rect 470090 334294 470158 334350
rect 470214 334294 470282 334350
rect 470338 334294 470406 334350
rect 470462 334294 470558 334350
rect 469938 334226 470558 334294
rect 469938 334170 470034 334226
rect 470090 334170 470158 334226
rect 470214 334170 470282 334226
rect 470338 334170 470406 334226
rect 470462 334170 470558 334226
rect 469938 334102 470558 334170
rect 469938 334046 470034 334102
rect 470090 334046 470158 334102
rect 470214 334046 470282 334102
rect 470338 334046 470406 334102
rect 470462 334046 470558 334102
rect 469938 333978 470558 334046
rect 469938 333922 470034 333978
rect 470090 333922 470158 333978
rect 470214 333922 470282 333978
rect 470338 333922 470406 333978
rect 470462 333922 470558 333978
rect 469938 316350 470558 333922
rect 469938 316294 470034 316350
rect 470090 316294 470158 316350
rect 470214 316294 470282 316350
rect 470338 316294 470406 316350
rect 470462 316294 470558 316350
rect 469938 316226 470558 316294
rect 469938 316170 470034 316226
rect 470090 316170 470158 316226
rect 470214 316170 470282 316226
rect 470338 316170 470406 316226
rect 470462 316170 470558 316226
rect 469938 316102 470558 316170
rect 469938 316046 470034 316102
rect 470090 316046 470158 316102
rect 470214 316046 470282 316102
rect 470338 316046 470406 316102
rect 470462 316046 470558 316102
rect 469938 315978 470558 316046
rect 469938 315922 470034 315978
rect 470090 315922 470158 315978
rect 470214 315922 470282 315978
rect 470338 315922 470406 315978
rect 470462 315922 470558 315978
rect 469938 298350 470558 315922
rect 469938 298294 470034 298350
rect 470090 298294 470158 298350
rect 470214 298294 470282 298350
rect 470338 298294 470406 298350
rect 470462 298294 470558 298350
rect 469938 298226 470558 298294
rect 469938 298170 470034 298226
rect 470090 298170 470158 298226
rect 470214 298170 470282 298226
rect 470338 298170 470406 298226
rect 470462 298170 470558 298226
rect 469938 298102 470558 298170
rect 469938 298046 470034 298102
rect 470090 298046 470158 298102
rect 470214 298046 470282 298102
rect 470338 298046 470406 298102
rect 470462 298046 470558 298102
rect 469938 297978 470558 298046
rect 469938 297922 470034 297978
rect 470090 297922 470158 297978
rect 470214 297922 470282 297978
rect 470338 297922 470406 297978
rect 470462 297922 470558 297978
rect 469938 280350 470558 297922
rect 469938 280294 470034 280350
rect 470090 280294 470158 280350
rect 470214 280294 470282 280350
rect 470338 280294 470406 280350
rect 470462 280294 470558 280350
rect 469938 280226 470558 280294
rect 469938 280170 470034 280226
rect 470090 280170 470158 280226
rect 470214 280170 470282 280226
rect 470338 280170 470406 280226
rect 470462 280170 470558 280226
rect 469938 280102 470558 280170
rect 469938 280046 470034 280102
rect 470090 280046 470158 280102
rect 470214 280046 470282 280102
rect 470338 280046 470406 280102
rect 470462 280046 470558 280102
rect 469938 279978 470558 280046
rect 469938 279922 470034 279978
rect 470090 279922 470158 279978
rect 470214 279922 470282 279978
rect 470338 279922 470406 279978
rect 470462 279922 470558 279978
rect 469938 262350 470558 279922
rect 469938 262294 470034 262350
rect 470090 262294 470158 262350
rect 470214 262294 470282 262350
rect 470338 262294 470406 262350
rect 470462 262294 470558 262350
rect 469938 262226 470558 262294
rect 469938 262170 470034 262226
rect 470090 262170 470158 262226
rect 470214 262170 470282 262226
rect 470338 262170 470406 262226
rect 470462 262170 470558 262226
rect 469938 262102 470558 262170
rect 469938 262046 470034 262102
rect 470090 262046 470158 262102
rect 470214 262046 470282 262102
rect 470338 262046 470406 262102
rect 470462 262046 470558 262102
rect 469938 261978 470558 262046
rect 469938 261922 470034 261978
rect 470090 261922 470158 261978
rect 470214 261922 470282 261978
rect 470338 261922 470406 261978
rect 470462 261922 470558 261978
rect 469938 244350 470558 261922
rect 469938 244294 470034 244350
rect 470090 244294 470158 244350
rect 470214 244294 470282 244350
rect 470338 244294 470406 244350
rect 470462 244294 470558 244350
rect 469938 244226 470558 244294
rect 469938 244170 470034 244226
rect 470090 244170 470158 244226
rect 470214 244170 470282 244226
rect 470338 244170 470406 244226
rect 470462 244170 470558 244226
rect 469938 244102 470558 244170
rect 469938 244046 470034 244102
rect 470090 244046 470158 244102
rect 470214 244046 470282 244102
rect 470338 244046 470406 244102
rect 470462 244046 470558 244102
rect 469938 243978 470558 244046
rect 469938 243922 470034 243978
rect 470090 243922 470158 243978
rect 470214 243922 470282 243978
rect 470338 243922 470406 243978
rect 470462 243922 470558 243978
rect 469938 226350 470558 243922
rect 469938 226294 470034 226350
rect 470090 226294 470158 226350
rect 470214 226294 470282 226350
rect 470338 226294 470406 226350
rect 470462 226294 470558 226350
rect 469938 226226 470558 226294
rect 469938 226170 470034 226226
rect 470090 226170 470158 226226
rect 470214 226170 470282 226226
rect 470338 226170 470406 226226
rect 470462 226170 470558 226226
rect 469938 226102 470558 226170
rect 469938 226046 470034 226102
rect 470090 226046 470158 226102
rect 470214 226046 470282 226102
rect 470338 226046 470406 226102
rect 470462 226046 470558 226102
rect 469938 225978 470558 226046
rect 469938 225922 470034 225978
rect 470090 225922 470158 225978
rect 470214 225922 470282 225978
rect 470338 225922 470406 225978
rect 470462 225922 470558 225978
rect 469938 208350 470558 225922
rect 469938 208294 470034 208350
rect 470090 208294 470158 208350
rect 470214 208294 470282 208350
rect 470338 208294 470406 208350
rect 470462 208294 470558 208350
rect 469938 208226 470558 208294
rect 469938 208170 470034 208226
rect 470090 208170 470158 208226
rect 470214 208170 470282 208226
rect 470338 208170 470406 208226
rect 470462 208170 470558 208226
rect 469938 208102 470558 208170
rect 469938 208046 470034 208102
rect 470090 208046 470158 208102
rect 470214 208046 470282 208102
rect 470338 208046 470406 208102
rect 470462 208046 470558 208102
rect 469938 207978 470558 208046
rect 469938 207922 470034 207978
rect 470090 207922 470158 207978
rect 470214 207922 470282 207978
rect 470338 207922 470406 207978
rect 470462 207922 470558 207978
rect 469938 190350 470558 207922
rect 469938 190294 470034 190350
rect 470090 190294 470158 190350
rect 470214 190294 470282 190350
rect 470338 190294 470406 190350
rect 470462 190294 470558 190350
rect 469938 190226 470558 190294
rect 469938 190170 470034 190226
rect 470090 190170 470158 190226
rect 470214 190170 470282 190226
rect 470338 190170 470406 190226
rect 470462 190170 470558 190226
rect 469938 190102 470558 190170
rect 469938 190046 470034 190102
rect 470090 190046 470158 190102
rect 470214 190046 470282 190102
rect 470338 190046 470406 190102
rect 470462 190046 470558 190102
rect 469938 189978 470558 190046
rect 469938 189922 470034 189978
rect 470090 189922 470158 189978
rect 470214 189922 470282 189978
rect 470338 189922 470406 189978
rect 470462 189922 470558 189978
rect 469938 172350 470558 189922
rect 469938 172294 470034 172350
rect 470090 172294 470158 172350
rect 470214 172294 470282 172350
rect 470338 172294 470406 172350
rect 470462 172294 470558 172350
rect 469938 172226 470558 172294
rect 469938 172170 470034 172226
rect 470090 172170 470158 172226
rect 470214 172170 470282 172226
rect 470338 172170 470406 172226
rect 470462 172170 470558 172226
rect 469938 172102 470558 172170
rect 469938 172046 470034 172102
rect 470090 172046 470158 172102
rect 470214 172046 470282 172102
rect 470338 172046 470406 172102
rect 470462 172046 470558 172102
rect 469938 171978 470558 172046
rect 469938 171922 470034 171978
rect 470090 171922 470158 171978
rect 470214 171922 470282 171978
rect 470338 171922 470406 171978
rect 470462 171922 470558 171978
rect 469938 154350 470558 171922
rect 469938 154294 470034 154350
rect 470090 154294 470158 154350
rect 470214 154294 470282 154350
rect 470338 154294 470406 154350
rect 470462 154294 470558 154350
rect 469938 154226 470558 154294
rect 469938 154170 470034 154226
rect 470090 154170 470158 154226
rect 470214 154170 470282 154226
rect 470338 154170 470406 154226
rect 470462 154170 470558 154226
rect 469938 154102 470558 154170
rect 469938 154046 470034 154102
rect 470090 154046 470158 154102
rect 470214 154046 470282 154102
rect 470338 154046 470406 154102
rect 470462 154046 470558 154102
rect 469938 153978 470558 154046
rect 469938 153922 470034 153978
rect 470090 153922 470158 153978
rect 470214 153922 470282 153978
rect 470338 153922 470406 153978
rect 470462 153922 470558 153978
rect 469938 136350 470558 153922
rect 469938 136294 470034 136350
rect 470090 136294 470158 136350
rect 470214 136294 470282 136350
rect 470338 136294 470406 136350
rect 470462 136294 470558 136350
rect 469938 136226 470558 136294
rect 469938 136170 470034 136226
rect 470090 136170 470158 136226
rect 470214 136170 470282 136226
rect 470338 136170 470406 136226
rect 470462 136170 470558 136226
rect 469938 136102 470558 136170
rect 469938 136046 470034 136102
rect 470090 136046 470158 136102
rect 470214 136046 470282 136102
rect 470338 136046 470406 136102
rect 470462 136046 470558 136102
rect 469938 135978 470558 136046
rect 469938 135922 470034 135978
rect 470090 135922 470158 135978
rect 470214 135922 470282 135978
rect 470338 135922 470406 135978
rect 470462 135922 470558 135978
rect 469938 118350 470558 135922
rect 469938 118294 470034 118350
rect 470090 118294 470158 118350
rect 470214 118294 470282 118350
rect 470338 118294 470406 118350
rect 470462 118294 470558 118350
rect 469938 118226 470558 118294
rect 469938 118170 470034 118226
rect 470090 118170 470158 118226
rect 470214 118170 470282 118226
rect 470338 118170 470406 118226
rect 470462 118170 470558 118226
rect 469938 118102 470558 118170
rect 469938 118046 470034 118102
rect 470090 118046 470158 118102
rect 470214 118046 470282 118102
rect 470338 118046 470406 118102
rect 470462 118046 470558 118102
rect 469938 117978 470558 118046
rect 469938 117922 470034 117978
rect 470090 117922 470158 117978
rect 470214 117922 470282 117978
rect 470338 117922 470406 117978
rect 470462 117922 470558 117978
rect 469938 100350 470558 117922
rect 469938 100294 470034 100350
rect 470090 100294 470158 100350
rect 470214 100294 470282 100350
rect 470338 100294 470406 100350
rect 470462 100294 470558 100350
rect 469938 100226 470558 100294
rect 469938 100170 470034 100226
rect 470090 100170 470158 100226
rect 470214 100170 470282 100226
rect 470338 100170 470406 100226
rect 470462 100170 470558 100226
rect 469938 100102 470558 100170
rect 469938 100046 470034 100102
rect 470090 100046 470158 100102
rect 470214 100046 470282 100102
rect 470338 100046 470406 100102
rect 470462 100046 470558 100102
rect 469938 99978 470558 100046
rect 469938 99922 470034 99978
rect 470090 99922 470158 99978
rect 470214 99922 470282 99978
rect 470338 99922 470406 99978
rect 470462 99922 470558 99978
rect 469938 82350 470558 99922
rect 496938 597212 497558 598268
rect 496938 597156 497034 597212
rect 497090 597156 497158 597212
rect 497214 597156 497282 597212
rect 497338 597156 497406 597212
rect 497462 597156 497558 597212
rect 496938 597088 497558 597156
rect 496938 597032 497034 597088
rect 497090 597032 497158 597088
rect 497214 597032 497282 597088
rect 497338 597032 497406 597088
rect 497462 597032 497558 597088
rect 496938 596964 497558 597032
rect 496938 596908 497034 596964
rect 497090 596908 497158 596964
rect 497214 596908 497282 596964
rect 497338 596908 497406 596964
rect 497462 596908 497558 596964
rect 496938 596840 497558 596908
rect 496938 596784 497034 596840
rect 497090 596784 497158 596840
rect 497214 596784 497282 596840
rect 497338 596784 497406 596840
rect 497462 596784 497558 596840
rect 496938 580350 497558 596784
rect 496938 580294 497034 580350
rect 497090 580294 497158 580350
rect 497214 580294 497282 580350
rect 497338 580294 497406 580350
rect 497462 580294 497558 580350
rect 496938 580226 497558 580294
rect 496938 580170 497034 580226
rect 497090 580170 497158 580226
rect 497214 580170 497282 580226
rect 497338 580170 497406 580226
rect 497462 580170 497558 580226
rect 496938 580102 497558 580170
rect 496938 580046 497034 580102
rect 497090 580046 497158 580102
rect 497214 580046 497282 580102
rect 497338 580046 497406 580102
rect 497462 580046 497558 580102
rect 496938 579978 497558 580046
rect 496938 579922 497034 579978
rect 497090 579922 497158 579978
rect 497214 579922 497282 579978
rect 497338 579922 497406 579978
rect 497462 579922 497558 579978
rect 496938 562350 497558 579922
rect 496938 562294 497034 562350
rect 497090 562294 497158 562350
rect 497214 562294 497282 562350
rect 497338 562294 497406 562350
rect 497462 562294 497558 562350
rect 496938 562226 497558 562294
rect 496938 562170 497034 562226
rect 497090 562170 497158 562226
rect 497214 562170 497282 562226
rect 497338 562170 497406 562226
rect 497462 562170 497558 562226
rect 496938 562102 497558 562170
rect 496938 562046 497034 562102
rect 497090 562046 497158 562102
rect 497214 562046 497282 562102
rect 497338 562046 497406 562102
rect 497462 562046 497558 562102
rect 496938 561978 497558 562046
rect 496938 561922 497034 561978
rect 497090 561922 497158 561978
rect 497214 561922 497282 561978
rect 497338 561922 497406 561978
rect 497462 561922 497558 561978
rect 496938 544350 497558 561922
rect 496938 544294 497034 544350
rect 497090 544294 497158 544350
rect 497214 544294 497282 544350
rect 497338 544294 497406 544350
rect 497462 544294 497558 544350
rect 496938 544226 497558 544294
rect 496938 544170 497034 544226
rect 497090 544170 497158 544226
rect 497214 544170 497282 544226
rect 497338 544170 497406 544226
rect 497462 544170 497558 544226
rect 496938 544102 497558 544170
rect 496938 544046 497034 544102
rect 497090 544046 497158 544102
rect 497214 544046 497282 544102
rect 497338 544046 497406 544102
rect 497462 544046 497558 544102
rect 496938 543978 497558 544046
rect 496938 543922 497034 543978
rect 497090 543922 497158 543978
rect 497214 543922 497282 543978
rect 497338 543922 497406 543978
rect 497462 543922 497558 543978
rect 496938 526350 497558 543922
rect 496938 526294 497034 526350
rect 497090 526294 497158 526350
rect 497214 526294 497282 526350
rect 497338 526294 497406 526350
rect 497462 526294 497558 526350
rect 496938 526226 497558 526294
rect 496938 526170 497034 526226
rect 497090 526170 497158 526226
rect 497214 526170 497282 526226
rect 497338 526170 497406 526226
rect 497462 526170 497558 526226
rect 496938 526102 497558 526170
rect 496938 526046 497034 526102
rect 497090 526046 497158 526102
rect 497214 526046 497282 526102
rect 497338 526046 497406 526102
rect 497462 526046 497558 526102
rect 496938 525978 497558 526046
rect 496938 525922 497034 525978
rect 497090 525922 497158 525978
rect 497214 525922 497282 525978
rect 497338 525922 497406 525978
rect 497462 525922 497558 525978
rect 496938 508350 497558 525922
rect 496938 508294 497034 508350
rect 497090 508294 497158 508350
rect 497214 508294 497282 508350
rect 497338 508294 497406 508350
rect 497462 508294 497558 508350
rect 496938 508226 497558 508294
rect 496938 508170 497034 508226
rect 497090 508170 497158 508226
rect 497214 508170 497282 508226
rect 497338 508170 497406 508226
rect 497462 508170 497558 508226
rect 496938 508102 497558 508170
rect 496938 508046 497034 508102
rect 497090 508046 497158 508102
rect 497214 508046 497282 508102
rect 497338 508046 497406 508102
rect 497462 508046 497558 508102
rect 496938 507978 497558 508046
rect 496938 507922 497034 507978
rect 497090 507922 497158 507978
rect 497214 507922 497282 507978
rect 497338 507922 497406 507978
rect 497462 507922 497558 507978
rect 496938 490350 497558 507922
rect 496938 490294 497034 490350
rect 497090 490294 497158 490350
rect 497214 490294 497282 490350
rect 497338 490294 497406 490350
rect 497462 490294 497558 490350
rect 496938 490226 497558 490294
rect 496938 490170 497034 490226
rect 497090 490170 497158 490226
rect 497214 490170 497282 490226
rect 497338 490170 497406 490226
rect 497462 490170 497558 490226
rect 496938 490102 497558 490170
rect 496938 490046 497034 490102
rect 497090 490046 497158 490102
rect 497214 490046 497282 490102
rect 497338 490046 497406 490102
rect 497462 490046 497558 490102
rect 496938 489978 497558 490046
rect 496938 489922 497034 489978
rect 497090 489922 497158 489978
rect 497214 489922 497282 489978
rect 497338 489922 497406 489978
rect 497462 489922 497558 489978
rect 496938 472350 497558 489922
rect 496938 472294 497034 472350
rect 497090 472294 497158 472350
rect 497214 472294 497282 472350
rect 497338 472294 497406 472350
rect 497462 472294 497558 472350
rect 496938 472226 497558 472294
rect 496938 472170 497034 472226
rect 497090 472170 497158 472226
rect 497214 472170 497282 472226
rect 497338 472170 497406 472226
rect 497462 472170 497558 472226
rect 496938 472102 497558 472170
rect 496938 472046 497034 472102
rect 497090 472046 497158 472102
rect 497214 472046 497282 472102
rect 497338 472046 497406 472102
rect 497462 472046 497558 472102
rect 496938 471978 497558 472046
rect 496938 471922 497034 471978
rect 497090 471922 497158 471978
rect 497214 471922 497282 471978
rect 497338 471922 497406 471978
rect 497462 471922 497558 471978
rect 496938 454350 497558 471922
rect 496938 454294 497034 454350
rect 497090 454294 497158 454350
rect 497214 454294 497282 454350
rect 497338 454294 497406 454350
rect 497462 454294 497558 454350
rect 496938 454226 497558 454294
rect 496938 454170 497034 454226
rect 497090 454170 497158 454226
rect 497214 454170 497282 454226
rect 497338 454170 497406 454226
rect 497462 454170 497558 454226
rect 496938 454102 497558 454170
rect 496938 454046 497034 454102
rect 497090 454046 497158 454102
rect 497214 454046 497282 454102
rect 497338 454046 497406 454102
rect 497462 454046 497558 454102
rect 496938 453978 497558 454046
rect 496938 453922 497034 453978
rect 497090 453922 497158 453978
rect 497214 453922 497282 453978
rect 497338 453922 497406 453978
rect 497462 453922 497558 453978
rect 496938 436350 497558 453922
rect 496938 436294 497034 436350
rect 497090 436294 497158 436350
rect 497214 436294 497282 436350
rect 497338 436294 497406 436350
rect 497462 436294 497558 436350
rect 496938 436226 497558 436294
rect 496938 436170 497034 436226
rect 497090 436170 497158 436226
rect 497214 436170 497282 436226
rect 497338 436170 497406 436226
rect 497462 436170 497558 436226
rect 496938 436102 497558 436170
rect 496938 436046 497034 436102
rect 497090 436046 497158 436102
rect 497214 436046 497282 436102
rect 497338 436046 497406 436102
rect 497462 436046 497558 436102
rect 496938 435978 497558 436046
rect 496938 435922 497034 435978
rect 497090 435922 497158 435978
rect 497214 435922 497282 435978
rect 497338 435922 497406 435978
rect 497462 435922 497558 435978
rect 496938 418350 497558 435922
rect 496938 418294 497034 418350
rect 497090 418294 497158 418350
rect 497214 418294 497282 418350
rect 497338 418294 497406 418350
rect 497462 418294 497558 418350
rect 496938 418226 497558 418294
rect 496938 418170 497034 418226
rect 497090 418170 497158 418226
rect 497214 418170 497282 418226
rect 497338 418170 497406 418226
rect 497462 418170 497558 418226
rect 496938 418102 497558 418170
rect 496938 418046 497034 418102
rect 497090 418046 497158 418102
rect 497214 418046 497282 418102
rect 497338 418046 497406 418102
rect 497462 418046 497558 418102
rect 496938 417978 497558 418046
rect 496938 417922 497034 417978
rect 497090 417922 497158 417978
rect 497214 417922 497282 417978
rect 497338 417922 497406 417978
rect 497462 417922 497558 417978
rect 496938 400350 497558 417922
rect 496938 400294 497034 400350
rect 497090 400294 497158 400350
rect 497214 400294 497282 400350
rect 497338 400294 497406 400350
rect 497462 400294 497558 400350
rect 496938 400226 497558 400294
rect 496938 400170 497034 400226
rect 497090 400170 497158 400226
rect 497214 400170 497282 400226
rect 497338 400170 497406 400226
rect 497462 400170 497558 400226
rect 496938 400102 497558 400170
rect 496938 400046 497034 400102
rect 497090 400046 497158 400102
rect 497214 400046 497282 400102
rect 497338 400046 497406 400102
rect 497462 400046 497558 400102
rect 496938 399978 497558 400046
rect 496938 399922 497034 399978
rect 497090 399922 497158 399978
rect 497214 399922 497282 399978
rect 497338 399922 497406 399978
rect 497462 399922 497558 399978
rect 496938 382350 497558 399922
rect 496938 382294 497034 382350
rect 497090 382294 497158 382350
rect 497214 382294 497282 382350
rect 497338 382294 497406 382350
rect 497462 382294 497558 382350
rect 496938 382226 497558 382294
rect 496938 382170 497034 382226
rect 497090 382170 497158 382226
rect 497214 382170 497282 382226
rect 497338 382170 497406 382226
rect 497462 382170 497558 382226
rect 496938 382102 497558 382170
rect 496938 382046 497034 382102
rect 497090 382046 497158 382102
rect 497214 382046 497282 382102
rect 497338 382046 497406 382102
rect 497462 382046 497558 382102
rect 496938 381978 497558 382046
rect 496938 381922 497034 381978
rect 497090 381922 497158 381978
rect 497214 381922 497282 381978
rect 497338 381922 497406 381978
rect 497462 381922 497558 381978
rect 496938 364350 497558 381922
rect 496938 364294 497034 364350
rect 497090 364294 497158 364350
rect 497214 364294 497282 364350
rect 497338 364294 497406 364350
rect 497462 364294 497558 364350
rect 496938 364226 497558 364294
rect 496938 364170 497034 364226
rect 497090 364170 497158 364226
rect 497214 364170 497282 364226
rect 497338 364170 497406 364226
rect 497462 364170 497558 364226
rect 496938 364102 497558 364170
rect 496938 364046 497034 364102
rect 497090 364046 497158 364102
rect 497214 364046 497282 364102
rect 497338 364046 497406 364102
rect 497462 364046 497558 364102
rect 496938 363978 497558 364046
rect 496938 363922 497034 363978
rect 497090 363922 497158 363978
rect 497214 363922 497282 363978
rect 497338 363922 497406 363978
rect 497462 363922 497558 363978
rect 496938 346350 497558 363922
rect 496938 346294 497034 346350
rect 497090 346294 497158 346350
rect 497214 346294 497282 346350
rect 497338 346294 497406 346350
rect 497462 346294 497558 346350
rect 496938 346226 497558 346294
rect 496938 346170 497034 346226
rect 497090 346170 497158 346226
rect 497214 346170 497282 346226
rect 497338 346170 497406 346226
rect 497462 346170 497558 346226
rect 496938 346102 497558 346170
rect 496938 346046 497034 346102
rect 497090 346046 497158 346102
rect 497214 346046 497282 346102
rect 497338 346046 497406 346102
rect 497462 346046 497558 346102
rect 496938 345978 497558 346046
rect 496938 345922 497034 345978
rect 497090 345922 497158 345978
rect 497214 345922 497282 345978
rect 497338 345922 497406 345978
rect 497462 345922 497558 345978
rect 496938 328350 497558 345922
rect 496938 328294 497034 328350
rect 497090 328294 497158 328350
rect 497214 328294 497282 328350
rect 497338 328294 497406 328350
rect 497462 328294 497558 328350
rect 496938 328226 497558 328294
rect 496938 328170 497034 328226
rect 497090 328170 497158 328226
rect 497214 328170 497282 328226
rect 497338 328170 497406 328226
rect 497462 328170 497558 328226
rect 496938 328102 497558 328170
rect 496938 328046 497034 328102
rect 497090 328046 497158 328102
rect 497214 328046 497282 328102
rect 497338 328046 497406 328102
rect 497462 328046 497558 328102
rect 496938 327978 497558 328046
rect 496938 327922 497034 327978
rect 497090 327922 497158 327978
rect 497214 327922 497282 327978
rect 497338 327922 497406 327978
rect 497462 327922 497558 327978
rect 496938 310350 497558 327922
rect 496938 310294 497034 310350
rect 497090 310294 497158 310350
rect 497214 310294 497282 310350
rect 497338 310294 497406 310350
rect 497462 310294 497558 310350
rect 496938 310226 497558 310294
rect 496938 310170 497034 310226
rect 497090 310170 497158 310226
rect 497214 310170 497282 310226
rect 497338 310170 497406 310226
rect 497462 310170 497558 310226
rect 496938 310102 497558 310170
rect 496938 310046 497034 310102
rect 497090 310046 497158 310102
rect 497214 310046 497282 310102
rect 497338 310046 497406 310102
rect 497462 310046 497558 310102
rect 496938 309978 497558 310046
rect 496938 309922 497034 309978
rect 497090 309922 497158 309978
rect 497214 309922 497282 309978
rect 497338 309922 497406 309978
rect 497462 309922 497558 309978
rect 496938 292350 497558 309922
rect 496938 292294 497034 292350
rect 497090 292294 497158 292350
rect 497214 292294 497282 292350
rect 497338 292294 497406 292350
rect 497462 292294 497558 292350
rect 496938 292226 497558 292294
rect 496938 292170 497034 292226
rect 497090 292170 497158 292226
rect 497214 292170 497282 292226
rect 497338 292170 497406 292226
rect 497462 292170 497558 292226
rect 496938 292102 497558 292170
rect 496938 292046 497034 292102
rect 497090 292046 497158 292102
rect 497214 292046 497282 292102
rect 497338 292046 497406 292102
rect 497462 292046 497558 292102
rect 496938 291978 497558 292046
rect 496938 291922 497034 291978
rect 497090 291922 497158 291978
rect 497214 291922 497282 291978
rect 497338 291922 497406 291978
rect 497462 291922 497558 291978
rect 496938 274350 497558 291922
rect 496938 274294 497034 274350
rect 497090 274294 497158 274350
rect 497214 274294 497282 274350
rect 497338 274294 497406 274350
rect 497462 274294 497558 274350
rect 496938 274226 497558 274294
rect 496938 274170 497034 274226
rect 497090 274170 497158 274226
rect 497214 274170 497282 274226
rect 497338 274170 497406 274226
rect 497462 274170 497558 274226
rect 496938 274102 497558 274170
rect 496938 274046 497034 274102
rect 497090 274046 497158 274102
rect 497214 274046 497282 274102
rect 497338 274046 497406 274102
rect 497462 274046 497558 274102
rect 496938 273978 497558 274046
rect 496938 273922 497034 273978
rect 497090 273922 497158 273978
rect 497214 273922 497282 273978
rect 497338 273922 497406 273978
rect 497462 273922 497558 273978
rect 496938 256350 497558 273922
rect 496938 256294 497034 256350
rect 497090 256294 497158 256350
rect 497214 256294 497282 256350
rect 497338 256294 497406 256350
rect 497462 256294 497558 256350
rect 496938 256226 497558 256294
rect 496938 256170 497034 256226
rect 497090 256170 497158 256226
rect 497214 256170 497282 256226
rect 497338 256170 497406 256226
rect 497462 256170 497558 256226
rect 496938 256102 497558 256170
rect 496938 256046 497034 256102
rect 497090 256046 497158 256102
rect 497214 256046 497282 256102
rect 497338 256046 497406 256102
rect 497462 256046 497558 256102
rect 496938 255978 497558 256046
rect 496938 255922 497034 255978
rect 497090 255922 497158 255978
rect 497214 255922 497282 255978
rect 497338 255922 497406 255978
rect 497462 255922 497558 255978
rect 496938 238350 497558 255922
rect 496938 238294 497034 238350
rect 497090 238294 497158 238350
rect 497214 238294 497282 238350
rect 497338 238294 497406 238350
rect 497462 238294 497558 238350
rect 496938 238226 497558 238294
rect 496938 238170 497034 238226
rect 497090 238170 497158 238226
rect 497214 238170 497282 238226
rect 497338 238170 497406 238226
rect 497462 238170 497558 238226
rect 496938 238102 497558 238170
rect 496938 238046 497034 238102
rect 497090 238046 497158 238102
rect 497214 238046 497282 238102
rect 497338 238046 497406 238102
rect 497462 238046 497558 238102
rect 496938 237978 497558 238046
rect 496938 237922 497034 237978
rect 497090 237922 497158 237978
rect 497214 237922 497282 237978
rect 497338 237922 497406 237978
rect 497462 237922 497558 237978
rect 496938 220350 497558 237922
rect 496938 220294 497034 220350
rect 497090 220294 497158 220350
rect 497214 220294 497282 220350
rect 497338 220294 497406 220350
rect 497462 220294 497558 220350
rect 496938 220226 497558 220294
rect 496938 220170 497034 220226
rect 497090 220170 497158 220226
rect 497214 220170 497282 220226
rect 497338 220170 497406 220226
rect 497462 220170 497558 220226
rect 496938 220102 497558 220170
rect 496938 220046 497034 220102
rect 497090 220046 497158 220102
rect 497214 220046 497282 220102
rect 497338 220046 497406 220102
rect 497462 220046 497558 220102
rect 496938 219978 497558 220046
rect 496938 219922 497034 219978
rect 497090 219922 497158 219978
rect 497214 219922 497282 219978
rect 497338 219922 497406 219978
rect 497462 219922 497558 219978
rect 496938 202350 497558 219922
rect 496938 202294 497034 202350
rect 497090 202294 497158 202350
rect 497214 202294 497282 202350
rect 497338 202294 497406 202350
rect 497462 202294 497558 202350
rect 496938 202226 497558 202294
rect 496938 202170 497034 202226
rect 497090 202170 497158 202226
rect 497214 202170 497282 202226
rect 497338 202170 497406 202226
rect 497462 202170 497558 202226
rect 496938 202102 497558 202170
rect 496938 202046 497034 202102
rect 497090 202046 497158 202102
rect 497214 202046 497282 202102
rect 497338 202046 497406 202102
rect 497462 202046 497558 202102
rect 496938 201978 497558 202046
rect 496938 201922 497034 201978
rect 497090 201922 497158 201978
rect 497214 201922 497282 201978
rect 497338 201922 497406 201978
rect 497462 201922 497558 201978
rect 496938 184350 497558 201922
rect 496938 184294 497034 184350
rect 497090 184294 497158 184350
rect 497214 184294 497282 184350
rect 497338 184294 497406 184350
rect 497462 184294 497558 184350
rect 496938 184226 497558 184294
rect 496938 184170 497034 184226
rect 497090 184170 497158 184226
rect 497214 184170 497282 184226
rect 497338 184170 497406 184226
rect 497462 184170 497558 184226
rect 496938 184102 497558 184170
rect 496938 184046 497034 184102
rect 497090 184046 497158 184102
rect 497214 184046 497282 184102
rect 497338 184046 497406 184102
rect 497462 184046 497558 184102
rect 496938 183978 497558 184046
rect 496938 183922 497034 183978
rect 497090 183922 497158 183978
rect 497214 183922 497282 183978
rect 497338 183922 497406 183978
rect 497462 183922 497558 183978
rect 496938 166350 497558 183922
rect 496938 166294 497034 166350
rect 497090 166294 497158 166350
rect 497214 166294 497282 166350
rect 497338 166294 497406 166350
rect 497462 166294 497558 166350
rect 496938 166226 497558 166294
rect 496938 166170 497034 166226
rect 497090 166170 497158 166226
rect 497214 166170 497282 166226
rect 497338 166170 497406 166226
rect 497462 166170 497558 166226
rect 496938 166102 497558 166170
rect 496938 166046 497034 166102
rect 497090 166046 497158 166102
rect 497214 166046 497282 166102
rect 497338 166046 497406 166102
rect 497462 166046 497558 166102
rect 496938 165978 497558 166046
rect 496938 165922 497034 165978
rect 497090 165922 497158 165978
rect 497214 165922 497282 165978
rect 497338 165922 497406 165978
rect 497462 165922 497558 165978
rect 496938 148350 497558 165922
rect 496938 148294 497034 148350
rect 497090 148294 497158 148350
rect 497214 148294 497282 148350
rect 497338 148294 497406 148350
rect 497462 148294 497558 148350
rect 496938 148226 497558 148294
rect 496938 148170 497034 148226
rect 497090 148170 497158 148226
rect 497214 148170 497282 148226
rect 497338 148170 497406 148226
rect 497462 148170 497558 148226
rect 496938 148102 497558 148170
rect 496938 148046 497034 148102
rect 497090 148046 497158 148102
rect 497214 148046 497282 148102
rect 497338 148046 497406 148102
rect 497462 148046 497558 148102
rect 496938 147978 497558 148046
rect 496938 147922 497034 147978
rect 497090 147922 497158 147978
rect 497214 147922 497282 147978
rect 497338 147922 497406 147978
rect 497462 147922 497558 147978
rect 496938 130350 497558 147922
rect 496938 130294 497034 130350
rect 497090 130294 497158 130350
rect 497214 130294 497282 130350
rect 497338 130294 497406 130350
rect 497462 130294 497558 130350
rect 496938 130226 497558 130294
rect 496938 130170 497034 130226
rect 497090 130170 497158 130226
rect 497214 130170 497282 130226
rect 497338 130170 497406 130226
rect 497462 130170 497558 130226
rect 496938 130102 497558 130170
rect 496938 130046 497034 130102
rect 497090 130046 497158 130102
rect 497214 130046 497282 130102
rect 497338 130046 497406 130102
rect 497462 130046 497558 130102
rect 496938 129978 497558 130046
rect 496938 129922 497034 129978
rect 497090 129922 497158 129978
rect 497214 129922 497282 129978
rect 497338 129922 497406 129978
rect 497462 129922 497558 129978
rect 496938 112350 497558 129922
rect 496938 112294 497034 112350
rect 497090 112294 497158 112350
rect 497214 112294 497282 112350
rect 497338 112294 497406 112350
rect 497462 112294 497558 112350
rect 496938 112226 497558 112294
rect 496938 112170 497034 112226
rect 497090 112170 497158 112226
rect 497214 112170 497282 112226
rect 497338 112170 497406 112226
rect 497462 112170 497558 112226
rect 496938 112102 497558 112170
rect 496938 112046 497034 112102
rect 497090 112046 497158 112102
rect 497214 112046 497282 112102
rect 497338 112046 497406 112102
rect 497462 112046 497558 112102
rect 496938 111978 497558 112046
rect 496938 111922 497034 111978
rect 497090 111922 497158 111978
rect 497214 111922 497282 111978
rect 497338 111922 497406 111978
rect 497462 111922 497558 111978
rect 469938 82294 470034 82350
rect 470090 82294 470158 82350
rect 470214 82294 470282 82350
rect 470338 82294 470406 82350
rect 470462 82294 470558 82350
rect 469938 82226 470558 82294
rect 469938 82170 470034 82226
rect 470090 82170 470158 82226
rect 470214 82170 470282 82226
rect 470338 82170 470406 82226
rect 470462 82170 470558 82226
rect 469938 82102 470558 82170
rect 469938 82046 470034 82102
rect 470090 82046 470158 82102
rect 470214 82046 470282 82102
rect 470338 82046 470406 82102
rect 470462 82046 470558 82102
rect 469938 81978 470558 82046
rect 469938 81922 470034 81978
rect 470090 81922 470158 81978
rect 470214 81922 470282 81978
rect 470338 81922 470406 81978
rect 470462 81922 470558 81978
rect 466218 58294 466314 58350
rect 466370 58294 466438 58350
rect 466494 58294 466562 58350
rect 466618 58294 466686 58350
rect 466742 58294 466838 58350
rect 466218 58226 466838 58294
rect 466218 58170 466314 58226
rect 466370 58170 466438 58226
rect 466494 58170 466562 58226
rect 466618 58170 466686 58226
rect 466742 58170 466838 58226
rect 466218 58102 466838 58170
rect 466218 58046 466314 58102
rect 466370 58046 466438 58102
rect 466494 58046 466562 58102
rect 466618 58046 466686 58102
rect 466742 58046 466838 58102
rect 466218 57978 466838 58046
rect 466218 57922 466314 57978
rect 466370 57922 466438 57978
rect 466494 57922 466562 57978
rect 466618 57922 466686 57978
rect 466742 57922 466838 57978
rect 465388 52498 465444 52508
rect 460348 25498 460404 25508
rect 458668 20132 458836 20188
rect 453628 4162 453684 4172
rect 456988 8578 457044 8588
rect 456988 4228 457044 8522
rect 456988 4162 457044 4172
rect 458780 4228 458836 20132
rect 458780 4162 458836 4172
rect 460348 4228 460404 25442
rect 460348 4162 460404 4172
rect 462588 5158 462644 5168
rect 462588 3444 462644 5102
rect 465388 4228 465444 52442
rect 465388 4162 465444 4172
rect 466218 40350 466838 57922
rect 466218 40294 466314 40350
rect 466370 40294 466438 40350
rect 466494 40294 466562 40350
rect 466618 40294 466686 40350
rect 466742 40294 466838 40350
rect 466218 40226 466838 40294
rect 466218 40170 466314 40226
rect 466370 40170 466438 40226
rect 466494 40170 466562 40226
rect 466618 40170 466686 40226
rect 466742 40170 466838 40226
rect 466218 40102 466838 40170
rect 466218 40046 466314 40102
rect 466370 40046 466438 40102
rect 466494 40046 466562 40102
rect 466618 40046 466686 40102
rect 466742 40046 466838 40102
rect 466218 39978 466838 40046
rect 466218 39922 466314 39978
rect 466370 39922 466438 39978
rect 466494 39922 466562 39978
rect 466618 39922 466686 39978
rect 466742 39922 466838 39978
rect 466218 22350 466838 39922
rect 466218 22294 466314 22350
rect 466370 22294 466438 22350
rect 466494 22294 466562 22350
rect 466618 22294 466686 22350
rect 466742 22294 466838 22350
rect 466218 22226 466838 22294
rect 466218 22170 466314 22226
rect 466370 22170 466438 22226
rect 466494 22170 466562 22226
rect 466618 22170 466686 22226
rect 466742 22170 466838 22226
rect 466218 22102 466838 22170
rect 466218 22046 466314 22102
rect 466370 22046 466438 22102
rect 466494 22046 466562 22102
rect 466618 22046 466686 22102
rect 466742 22046 466838 22102
rect 466218 21978 466838 22046
rect 466218 21922 466314 21978
rect 466370 21922 466438 21978
rect 466494 21922 466562 21978
rect 466618 21922 466686 21978
rect 466742 21922 466838 21978
rect 466218 4350 466838 21922
rect 468748 72298 468804 72308
rect 466218 4294 466314 4350
rect 466370 4294 466438 4350
rect 466494 4294 466562 4350
rect 466618 4294 466686 4350
rect 466742 4294 466838 4350
rect 466218 4226 466838 4294
rect 466218 4170 466314 4226
rect 466370 4170 466438 4226
rect 466494 4170 466562 4226
rect 466618 4170 466686 4226
rect 466742 4170 466838 4226
rect 462588 3378 462644 3388
rect 466218 4102 466838 4170
rect 466218 4046 466314 4102
rect 466370 4046 466438 4102
rect 466494 4046 466562 4102
rect 466618 4046 466686 4102
rect 466742 4046 466838 4102
rect 466218 3978 466838 4046
rect 466218 3922 466314 3978
rect 466370 3922 466438 3978
rect 466494 3922 466562 3978
rect 466618 3922 466686 3978
rect 466742 3922 466838 3978
rect 439218 -1176 439314 -1120
rect 439370 -1176 439438 -1120
rect 439494 -1176 439562 -1120
rect 439618 -1176 439686 -1120
rect 439742 -1176 439838 -1120
rect 439218 -1244 439838 -1176
rect 439218 -1300 439314 -1244
rect 439370 -1300 439438 -1244
rect 439494 -1300 439562 -1244
rect 439618 -1300 439686 -1244
rect 439742 -1300 439838 -1244
rect 439218 -1368 439838 -1300
rect 439218 -1424 439314 -1368
rect 439370 -1424 439438 -1368
rect 439494 -1424 439562 -1368
rect 439618 -1424 439686 -1368
rect 439742 -1424 439838 -1368
rect 439218 -1492 439838 -1424
rect 439218 -1548 439314 -1492
rect 439370 -1548 439438 -1492
rect 439494 -1548 439562 -1492
rect 439618 -1548 439686 -1492
rect 439742 -1548 439838 -1492
rect 439218 -1644 439838 -1548
rect 466218 -160 466838 3922
rect 468300 6958 468356 6968
rect 468300 3556 468356 6902
rect 468748 4228 468804 72242
rect 468748 4162 468804 4172
rect 469938 64350 470558 81922
rect 469938 64294 470034 64350
rect 470090 64294 470158 64350
rect 470214 64294 470282 64350
rect 470338 64294 470406 64350
rect 470462 64294 470558 64350
rect 469938 64226 470558 64294
rect 469938 64170 470034 64226
rect 470090 64170 470158 64226
rect 470214 64170 470282 64226
rect 470338 64170 470406 64226
rect 470462 64170 470558 64226
rect 469938 64102 470558 64170
rect 469938 64046 470034 64102
rect 470090 64046 470158 64102
rect 470214 64046 470282 64102
rect 470338 64046 470406 64102
rect 470462 64046 470558 64102
rect 469938 63978 470558 64046
rect 469938 63922 470034 63978
rect 470090 63922 470158 63978
rect 470214 63922 470282 63978
rect 470338 63922 470406 63978
rect 470462 63922 470558 63978
rect 469938 46350 470558 63922
rect 474572 98308 474628 98318
rect 469938 46294 470034 46350
rect 470090 46294 470158 46350
rect 470214 46294 470282 46350
rect 470338 46294 470406 46350
rect 470462 46294 470558 46350
rect 469938 46226 470558 46294
rect 469938 46170 470034 46226
rect 470090 46170 470158 46226
rect 470214 46170 470282 46226
rect 470338 46170 470406 46226
rect 470462 46170 470558 46226
rect 469938 46102 470558 46170
rect 469938 46046 470034 46102
rect 470090 46046 470158 46102
rect 470214 46046 470282 46102
rect 470338 46046 470406 46102
rect 470462 46046 470558 46102
rect 469938 45978 470558 46046
rect 469938 45922 470034 45978
rect 470090 45922 470158 45978
rect 470214 45922 470282 45978
rect 470338 45922 470406 45978
rect 470462 45922 470558 45978
rect 469938 28350 470558 45922
rect 469938 28294 470034 28350
rect 470090 28294 470158 28350
rect 470214 28294 470282 28350
rect 470338 28294 470406 28350
rect 470462 28294 470558 28350
rect 469938 28226 470558 28294
rect 469938 28170 470034 28226
rect 470090 28170 470158 28226
rect 470214 28170 470282 28226
rect 470338 28170 470406 28226
rect 470462 28170 470558 28226
rect 469938 28102 470558 28170
rect 469938 28046 470034 28102
rect 470090 28046 470158 28102
rect 470214 28046 470282 28102
rect 470338 28046 470406 28102
rect 470462 28046 470558 28102
rect 469938 27978 470558 28046
rect 469938 27922 470034 27978
rect 470090 27922 470158 27978
rect 470214 27922 470282 27978
rect 470338 27922 470406 27978
rect 470462 27922 470558 27978
rect 469938 10350 470558 27922
rect 469938 10294 470034 10350
rect 470090 10294 470158 10350
rect 470214 10294 470282 10350
rect 470338 10294 470406 10350
rect 470462 10294 470558 10350
rect 469938 10226 470558 10294
rect 469938 10170 470034 10226
rect 470090 10170 470158 10226
rect 470214 10170 470282 10226
rect 470338 10170 470406 10226
rect 470462 10170 470558 10226
rect 469938 10102 470558 10170
rect 469938 10046 470034 10102
rect 470090 10046 470158 10102
rect 470214 10046 470282 10102
rect 470338 10046 470406 10102
rect 470462 10046 470558 10102
rect 469938 9978 470558 10046
rect 469938 9922 470034 9978
rect 470090 9922 470158 9978
rect 470214 9922 470282 9978
rect 470338 9922 470406 9978
rect 470462 9922 470558 9978
rect 468300 3490 468356 3500
rect 466218 -216 466314 -160
rect 466370 -216 466438 -160
rect 466494 -216 466562 -160
rect 466618 -216 466686 -160
rect 466742 -216 466838 -160
rect 466218 -284 466838 -216
rect 466218 -340 466314 -284
rect 466370 -340 466438 -284
rect 466494 -340 466562 -284
rect 466618 -340 466686 -284
rect 466742 -340 466838 -284
rect 466218 -408 466838 -340
rect 466218 -464 466314 -408
rect 466370 -464 466438 -408
rect 466494 -464 466562 -408
rect 466618 -464 466686 -408
rect 466742 -464 466838 -408
rect 466218 -532 466838 -464
rect 466218 -588 466314 -532
rect 466370 -588 466438 -532
rect 466494 -588 466562 -532
rect 466618 -588 466686 -532
rect 466742 -588 466838 -532
rect 466218 -1644 466838 -588
rect 469938 -1120 470558 9922
rect 472108 62398 472164 62408
rect 472108 4228 472164 62342
rect 474572 25956 474628 98252
rect 496938 94350 497558 111922
rect 496938 94294 497034 94350
rect 497090 94294 497158 94350
rect 497214 94294 497282 94350
rect 497338 94294 497406 94350
rect 497462 94294 497558 94350
rect 496938 94226 497558 94294
rect 496938 94170 497034 94226
rect 497090 94170 497158 94226
rect 497214 94170 497282 94226
rect 497338 94170 497406 94226
rect 497462 94170 497558 94226
rect 496938 94102 497558 94170
rect 496938 94046 497034 94102
rect 497090 94046 497158 94102
rect 497214 94046 497282 94102
rect 497338 94046 497406 94102
rect 497462 94046 497558 94102
rect 496938 93978 497558 94046
rect 496938 93922 497034 93978
rect 497090 93922 497158 93978
rect 497214 93922 497282 93978
rect 497338 93922 497406 93978
rect 497462 93922 497558 93978
rect 480508 79138 480564 79148
rect 477148 59158 477204 59168
rect 474572 25890 474628 25900
rect 475468 50878 475524 50888
rect 472108 4162 472164 4172
rect 474012 13618 474068 13628
rect 474012 4228 474068 13562
rect 474012 4162 474068 4172
rect 475468 4228 475524 50822
rect 475468 4162 475524 4172
rect 477148 4228 477204 59102
rect 477148 4162 477204 4172
rect 478828 15418 478884 15428
rect 478828 4228 478884 15362
rect 478828 4162 478884 4172
rect 480508 4228 480564 79082
rect 496938 76350 497558 93922
rect 500658 598172 501278 598268
rect 500658 598116 500754 598172
rect 500810 598116 500878 598172
rect 500934 598116 501002 598172
rect 501058 598116 501126 598172
rect 501182 598116 501278 598172
rect 500658 598048 501278 598116
rect 500658 597992 500754 598048
rect 500810 597992 500878 598048
rect 500934 597992 501002 598048
rect 501058 597992 501126 598048
rect 501182 597992 501278 598048
rect 500658 597924 501278 597992
rect 500658 597868 500754 597924
rect 500810 597868 500878 597924
rect 500934 597868 501002 597924
rect 501058 597868 501126 597924
rect 501182 597868 501278 597924
rect 500658 597800 501278 597868
rect 500658 597744 500754 597800
rect 500810 597744 500878 597800
rect 500934 597744 501002 597800
rect 501058 597744 501126 597800
rect 501182 597744 501278 597800
rect 500658 586350 501278 597744
rect 500658 586294 500754 586350
rect 500810 586294 500878 586350
rect 500934 586294 501002 586350
rect 501058 586294 501126 586350
rect 501182 586294 501278 586350
rect 500658 586226 501278 586294
rect 500658 586170 500754 586226
rect 500810 586170 500878 586226
rect 500934 586170 501002 586226
rect 501058 586170 501126 586226
rect 501182 586170 501278 586226
rect 500658 586102 501278 586170
rect 500658 586046 500754 586102
rect 500810 586046 500878 586102
rect 500934 586046 501002 586102
rect 501058 586046 501126 586102
rect 501182 586046 501278 586102
rect 500658 585978 501278 586046
rect 500658 585922 500754 585978
rect 500810 585922 500878 585978
rect 500934 585922 501002 585978
rect 501058 585922 501126 585978
rect 501182 585922 501278 585978
rect 500658 568350 501278 585922
rect 500658 568294 500754 568350
rect 500810 568294 500878 568350
rect 500934 568294 501002 568350
rect 501058 568294 501126 568350
rect 501182 568294 501278 568350
rect 500658 568226 501278 568294
rect 500658 568170 500754 568226
rect 500810 568170 500878 568226
rect 500934 568170 501002 568226
rect 501058 568170 501126 568226
rect 501182 568170 501278 568226
rect 500658 568102 501278 568170
rect 500658 568046 500754 568102
rect 500810 568046 500878 568102
rect 500934 568046 501002 568102
rect 501058 568046 501126 568102
rect 501182 568046 501278 568102
rect 500658 567978 501278 568046
rect 500658 567922 500754 567978
rect 500810 567922 500878 567978
rect 500934 567922 501002 567978
rect 501058 567922 501126 567978
rect 501182 567922 501278 567978
rect 500658 550350 501278 567922
rect 500658 550294 500754 550350
rect 500810 550294 500878 550350
rect 500934 550294 501002 550350
rect 501058 550294 501126 550350
rect 501182 550294 501278 550350
rect 500658 550226 501278 550294
rect 500658 550170 500754 550226
rect 500810 550170 500878 550226
rect 500934 550170 501002 550226
rect 501058 550170 501126 550226
rect 501182 550170 501278 550226
rect 500658 550102 501278 550170
rect 500658 550046 500754 550102
rect 500810 550046 500878 550102
rect 500934 550046 501002 550102
rect 501058 550046 501126 550102
rect 501182 550046 501278 550102
rect 500658 549978 501278 550046
rect 500658 549922 500754 549978
rect 500810 549922 500878 549978
rect 500934 549922 501002 549978
rect 501058 549922 501126 549978
rect 501182 549922 501278 549978
rect 500658 532350 501278 549922
rect 500658 532294 500754 532350
rect 500810 532294 500878 532350
rect 500934 532294 501002 532350
rect 501058 532294 501126 532350
rect 501182 532294 501278 532350
rect 500658 532226 501278 532294
rect 500658 532170 500754 532226
rect 500810 532170 500878 532226
rect 500934 532170 501002 532226
rect 501058 532170 501126 532226
rect 501182 532170 501278 532226
rect 500658 532102 501278 532170
rect 500658 532046 500754 532102
rect 500810 532046 500878 532102
rect 500934 532046 501002 532102
rect 501058 532046 501126 532102
rect 501182 532046 501278 532102
rect 500658 531978 501278 532046
rect 500658 531922 500754 531978
rect 500810 531922 500878 531978
rect 500934 531922 501002 531978
rect 501058 531922 501126 531978
rect 501182 531922 501278 531978
rect 500658 514350 501278 531922
rect 500658 514294 500754 514350
rect 500810 514294 500878 514350
rect 500934 514294 501002 514350
rect 501058 514294 501126 514350
rect 501182 514294 501278 514350
rect 500658 514226 501278 514294
rect 500658 514170 500754 514226
rect 500810 514170 500878 514226
rect 500934 514170 501002 514226
rect 501058 514170 501126 514226
rect 501182 514170 501278 514226
rect 500658 514102 501278 514170
rect 500658 514046 500754 514102
rect 500810 514046 500878 514102
rect 500934 514046 501002 514102
rect 501058 514046 501126 514102
rect 501182 514046 501278 514102
rect 500658 513978 501278 514046
rect 500658 513922 500754 513978
rect 500810 513922 500878 513978
rect 500934 513922 501002 513978
rect 501058 513922 501126 513978
rect 501182 513922 501278 513978
rect 500658 496350 501278 513922
rect 500658 496294 500754 496350
rect 500810 496294 500878 496350
rect 500934 496294 501002 496350
rect 501058 496294 501126 496350
rect 501182 496294 501278 496350
rect 500658 496226 501278 496294
rect 500658 496170 500754 496226
rect 500810 496170 500878 496226
rect 500934 496170 501002 496226
rect 501058 496170 501126 496226
rect 501182 496170 501278 496226
rect 500658 496102 501278 496170
rect 500658 496046 500754 496102
rect 500810 496046 500878 496102
rect 500934 496046 501002 496102
rect 501058 496046 501126 496102
rect 501182 496046 501278 496102
rect 500658 495978 501278 496046
rect 500658 495922 500754 495978
rect 500810 495922 500878 495978
rect 500934 495922 501002 495978
rect 501058 495922 501126 495978
rect 501182 495922 501278 495978
rect 500658 478350 501278 495922
rect 500658 478294 500754 478350
rect 500810 478294 500878 478350
rect 500934 478294 501002 478350
rect 501058 478294 501126 478350
rect 501182 478294 501278 478350
rect 500658 478226 501278 478294
rect 500658 478170 500754 478226
rect 500810 478170 500878 478226
rect 500934 478170 501002 478226
rect 501058 478170 501126 478226
rect 501182 478170 501278 478226
rect 500658 478102 501278 478170
rect 500658 478046 500754 478102
rect 500810 478046 500878 478102
rect 500934 478046 501002 478102
rect 501058 478046 501126 478102
rect 501182 478046 501278 478102
rect 500658 477978 501278 478046
rect 500658 477922 500754 477978
rect 500810 477922 500878 477978
rect 500934 477922 501002 477978
rect 501058 477922 501126 477978
rect 501182 477922 501278 477978
rect 500658 460350 501278 477922
rect 500658 460294 500754 460350
rect 500810 460294 500878 460350
rect 500934 460294 501002 460350
rect 501058 460294 501126 460350
rect 501182 460294 501278 460350
rect 500658 460226 501278 460294
rect 500658 460170 500754 460226
rect 500810 460170 500878 460226
rect 500934 460170 501002 460226
rect 501058 460170 501126 460226
rect 501182 460170 501278 460226
rect 500658 460102 501278 460170
rect 500658 460046 500754 460102
rect 500810 460046 500878 460102
rect 500934 460046 501002 460102
rect 501058 460046 501126 460102
rect 501182 460046 501278 460102
rect 500658 459978 501278 460046
rect 500658 459922 500754 459978
rect 500810 459922 500878 459978
rect 500934 459922 501002 459978
rect 501058 459922 501126 459978
rect 501182 459922 501278 459978
rect 500658 442350 501278 459922
rect 500658 442294 500754 442350
rect 500810 442294 500878 442350
rect 500934 442294 501002 442350
rect 501058 442294 501126 442350
rect 501182 442294 501278 442350
rect 500658 442226 501278 442294
rect 500658 442170 500754 442226
rect 500810 442170 500878 442226
rect 500934 442170 501002 442226
rect 501058 442170 501126 442226
rect 501182 442170 501278 442226
rect 500658 442102 501278 442170
rect 500658 442046 500754 442102
rect 500810 442046 500878 442102
rect 500934 442046 501002 442102
rect 501058 442046 501126 442102
rect 501182 442046 501278 442102
rect 500658 441978 501278 442046
rect 500658 441922 500754 441978
rect 500810 441922 500878 441978
rect 500934 441922 501002 441978
rect 501058 441922 501126 441978
rect 501182 441922 501278 441978
rect 500658 424350 501278 441922
rect 500658 424294 500754 424350
rect 500810 424294 500878 424350
rect 500934 424294 501002 424350
rect 501058 424294 501126 424350
rect 501182 424294 501278 424350
rect 500658 424226 501278 424294
rect 500658 424170 500754 424226
rect 500810 424170 500878 424226
rect 500934 424170 501002 424226
rect 501058 424170 501126 424226
rect 501182 424170 501278 424226
rect 500658 424102 501278 424170
rect 500658 424046 500754 424102
rect 500810 424046 500878 424102
rect 500934 424046 501002 424102
rect 501058 424046 501126 424102
rect 501182 424046 501278 424102
rect 500658 423978 501278 424046
rect 500658 423922 500754 423978
rect 500810 423922 500878 423978
rect 500934 423922 501002 423978
rect 501058 423922 501126 423978
rect 501182 423922 501278 423978
rect 500658 406350 501278 423922
rect 500658 406294 500754 406350
rect 500810 406294 500878 406350
rect 500934 406294 501002 406350
rect 501058 406294 501126 406350
rect 501182 406294 501278 406350
rect 500658 406226 501278 406294
rect 500658 406170 500754 406226
rect 500810 406170 500878 406226
rect 500934 406170 501002 406226
rect 501058 406170 501126 406226
rect 501182 406170 501278 406226
rect 500658 406102 501278 406170
rect 500658 406046 500754 406102
rect 500810 406046 500878 406102
rect 500934 406046 501002 406102
rect 501058 406046 501126 406102
rect 501182 406046 501278 406102
rect 500658 405978 501278 406046
rect 500658 405922 500754 405978
rect 500810 405922 500878 405978
rect 500934 405922 501002 405978
rect 501058 405922 501126 405978
rect 501182 405922 501278 405978
rect 500658 388350 501278 405922
rect 500658 388294 500754 388350
rect 500810 388294 500878 388350
rect 500934 388294 501002 388350
rect 501058 388294 501126 388350
rect 501182 388294 501278 388350
rect 500658 388226 501278 388294
rect 500658 388170 500754 388226
rect 500810 388170 500878 388226
rect 500934 388170 501002 388226
rect 501058 388170 501126 388226
rect 501182 388170 501278 388226
rect 500658 388102 501278 388170
rect 500658 388046 500754 388102
rect 500810 388046 500878 388102
rect 500934 388046 501002 388102
rect 501058 388046 501126 388102
rect 501182 388046 501278 388102
rect 500658 387978 501278 388046
rect 500658 387922 500754 387978
rect 500810 387922 500878 387978
rect 500934 387922 501002 387978
rect 501058 387922 501126 387978
rect 501182 387922 501278 387978
rect 500658 370350 501278 387922
rect 500658 370294 500754 370350
rect 500810 370294 500878 370350
rect 500934 370294 501002 370350
rect 501058 370294 501126 370350
rect 501182 370294 501278 370350
rect 500658 370226 501278 370294
rect 500658 370170 500754 370226
rect 500810 370170 500878 370226
rect 500934 370170 501002 370226
rect 501058 370170 501126 370226
rect 501182 370170 501278 370226
rect 500658 370102 501278 370170
rect 500658 370046 500754 370102
rect 500810 370046 500878 370102
rect 500934 370046 501002 370102
rect 501058 370046 501126 370102
rect 501182 370046 501278 370102
rect 500658 369978 501278 370046
rect 500658 369922 500754 369978
rect 500810 369922 500878 369978
rect 500934 369922 501002 369978
rect 501058 369922 501126 369978
rect 501182 369922 501278 369978
rect 500658 352350 501278 369922
rect 500658 352294 500754 352350
rect 500810 352294 500878 352350
rect 500934 352294 501002 352350
rect 501058 352294 501126 352350
rect 501182 352294 501278 352350
rect 500658 352226 501278 352294
rect 500658 352170 500754 352226
rect 500810 352170 500878 352226
rect 500934 352170 501002 352226
rect 501058 352170 501126 352226
rect 501182 352170 501278 352226
rect 500658 352102 501278 352170
rect 500658 352046 500754 352102
rect 500810 352046 500878 352102
rect 500934 352046 501002 352102
rect 501058 352046 501126 352102
rect 501182 352046 501278 352102
rect 500658 351978 501278 352046
rect 500658 351922 500754 351978
rect 500810 351922 500878 351978
rect 500934 351922 501002 351978
rect 501058 351922 501126 351978
rect 501182 351922 501278 351978
rect 500658 334350 501278 351922
rect 500658 334294 500754 334350
rect 500810 334294 500878 334350
rect 500934 334294 501002 334350
rect 501058 334294 501126 334350
rect 501182 334294 501278 334350
rect 500658 334226 501278 334294
rect 500658 334170 500754 334226
rect 500810 334170 500878 334226
rect 500934 334170 501002 334226
rect 501058 334170 501126 334226
rect 501182 334170 501278 334226
rect 500658 334102 501278 334170
rect 500658 334046 500754 334102
rect 500810 334046 500878 334102
rect 500934 334046 501002 334102
rect 501058 334046 501126 334102
rect 501182 334046 501278 334102
rect 500658 333978 501278 334046
rect 500658 333922 500754 333978
rect 500810 333922 500878 333978
rect 500934 333922 501002 333978
rect 501058 333922 501126 333978
rect 501182 333922 501278 333978
rect 500658 316350 501278 333922
rect 500658 316294 500754 316350
rect 500810 316294 500878 316350
rect 500934 316294 501002 316350
rect 501058 316294 501126 316350
rect 501182 316294 501278 316350
rect 500658 316226 501278 316294
rect 500658 316170 500754 316226
rect 500810 316170 500878 316226
rect 500934 316170 501002 316226
rect 501058 316170 501126 316226
rect 501182 316170 501278 316226
rect 500658 316102 501278 316170
rect 500658 316046 500754 316102
rect 500810 316046 500878 316102
rect 500934 316046 501002 316102
rect 501058 316046 501126 316102
rect 501182 316046 501278 316102
rect 500658 315978 501278 316046
rect 500658 315922 500754 315978
rect 500810 315922 500878 315978
rect 500934 315922 501002 315978
rect 501058 315922 501126 315978
rect 501182 315922 501278 315978
rect 500658 298350 501278 315922
rect 500658 298294 500754 298350
rect 500810 298294 500878 298350
rect 500934 298294 501002 298350
rect 501058 298294 501126 298350
rect 501182 298294 501278 298350
rect 500658 298226 501278 298294
rect 500658 298170 500754 298226
rect 500810 298170 500878 298226
rect 500934 298170 501002 298226
rect 501058 298170 501126 298226
rect 501182 298170 501278 298226
rect 500658 298102 501278 298170
rect 500658 298046 500754 298102
rect 500810 298046 500878 298102
rect 500934 298046 501002 298102
rect 501058 298046 501126 298102
rect 501182 298046 501278 298102
rect 500658 297978 501278 298046
rect 500658 297922 500754 297978
rect 500810 297922 500878 297978
rect 500934 297922 501002 297978
rect 501058 297922 501126 297978
rect 501182 297922 501278 297978
rect 500658 280350 501278 297922
rect 500658 280294 500754 280350
rect 500810 280294 500878 280350
rect 500934 280294 501002 280350
rect 501058 280294 501126 280350
rect 501182 280294 501278 280350
rect 500658 280226 501278 280294
rect 500658 280170 500754 280226
rect 500810 280170 500878 280226
rect 500934 280170 501002 280226
rect 501058 280170 501126 280226
rect 501182 280170 501278 280226
rect 500658 280102 501278 280170
rect 500658 280046 500754 280102
rect 500810 280046 500878 280102
rect 500934 280046 501002 280102
rect 501058 280046 501126 280102
rect 501182 280046 501278 280102
rect 500658 279978 501278 280046
rect 500658 279922 500754 279978
rect 500810 279922 500878 279978
rect 500934 279922 501002 279978
rect 501058 279922 501126 279978
rect 501182 279922 501278 279978
rect 500658 262350 501278 279922
rect 500658 262294 500754 262350
rect 500810 262294 500878 262350
rect 500934 262294 501002 262350
rect 501058 262294 501126 262350
rect 501182 262294 501278 262350
rect 500658 262226 501278 262294
rect 500658 262170 500754 262226
rect 500810 262170 500878 262226
rect 500934 262170 501002 262226
rect 501058 262170 501126 262226
rect 501182 262170 501278 262226
rect 500658 262102 501278 262170
rect 500658 262046 500754 262102
rect 500810 262046 500878 262102
rect 500934 262046 501002 262102
rect 501058 262046 501126 262102
rect 501182 262046 501278 262102
rect 500658 261978 501278 262046
rect 500658 261922 500754 261978
rect 500810 261922 500878 261978
rect 500934 261922 501002 261978
rect 501058 261922 501126 261978
rect 501182 261922 501278 261978
rect 500658 244350 501278 261922
rect 500658 244294 500754 244350
rect 500810 244294 500878 244350
rect 500934 244294 501002 244350
rect 501058 244294 501126 244350
rect 501182 244294 501278 244350
rect 500658 244226 501278 244294
rect 500658 244170 500754 244226
rect 500810 244170 500878 244226
rect 500934 244170 501002 244226
rect 501058 244170 501126 244226
rect 501182 244170 501278 244226
rect 500658 244102 501278 244170
rect 500658 244046 500754 244102
rect 500810 244046 500878 244102
rect 500934 244046 501002 244102
rect 501058 244046 501126 244102
rect 501182 244046 501278 244102
rect 500658 243978 501278 244046
rect 500658 243922 500754 243978
rect 500810 243922 500878 243978
rect 500934 243922 501002 243978
rect 501058 243922 501126 243978
rect 501182 243922 501278 243978
rect 500658 226350 501278 243922
rect 500658 226294 500754 226350
rect 500810 226294 500878 226350
rect 500934 226294 501002 226350
rect 501058 226294 501126 226350
rect 501182 226294 501278 226350
rect 500658 226226 501278 226294
rect 500658 226170 500754 226226
rect 500810 226170 500878 226226
rect 500934 226170 501002 226226
rect 501058 226170 501126 226226
rect 501182 226170 501278 226226
rect 500658 226102 501278 226170
rect 500658 226046 500754 226102
rect 500810 226046 500878 226102
rect 500934 226046 501002 226102
rect 501058 226046 501126 226102
rect 501182 226046 501278 226102
rect 500658 225978 501278 226046
rect 500658 225922 500754 225978
rect 500810 225922 500878 225978
rect 500934 225922 501002 225978
rect 501058 225922 501126 225978
rect 501182 225922 501278 225978
rect 500658 208350 501278 225922
rect 500658 208294 500754 208350
rect 500810 208294 500878 208350
rect 500934 208294 501002 208350
rect 501058 208294 501126 208350
rect 501182 208294 501278 208350
rect 500658 208226 501278 208294
rect 500658 208170 500754 208226
rect 500810 208170 500878 208226
rect 500934 208170 501002 208226
rect 501058 208170 501126 208226
rect 501182 208170 501278 208226
rect 500658 208102 501278 208170
rect 500658 208046 500754 208102
rect 500810 208046 500878 208102
rect 500934 208046 501002 208102
rect 501058 208046 501126 208102
rect 501182 208046 501278 208102
rect 500658 207978 501278 208046
rect 500658 207922 500754 207978
rect 500810 207922 500878 207978
rect 500934 207922 501002 207978
rect 501058 207922 501126 207978
rect 501182 207922 501278 207978
rect 500658 190350 501278 207922
rect 500658 190294 500754 190350
rect 500810 190294 500878 190350
rect 500934 190294 501002 190350
rect 501058 190294 501126 190350
rect 501182 190294 501278 190350
rect 500658 190226 501278 190294
rect 500658 190170 500754 190226
rect 500810 190170 500878 190226
rect 500934 190170 501002 190226
rect 501058 190170 501126 190226
rect 501182 190170 501278 190226
rect 500658 190102 501278 190170
rect 500658 190046 500754 190102
rect 500810 190046 500878 190102
rect 500934 190046 501002 190102
rect 501058 190046 501126 190102
rect 501182 190046 501278 190102
rect 500658 189978 501278 190046
rect 500658 189922 500754 189978
rect 500810 189922 500878 189978
rect 500934 189922 501002 189978
rect 501058 189922 501126 189978
rect 501182 189922 501278 189978
rect 500658 172350 501278 189922
rect 500658 172294 500754 172350
rect 500810 172294 500878 172350
rect 500934 172294 501002 172350
rect 501058 172294 501126 172350
rect 501182 172294 501278 172350
rect 500658 172226 501278 172294
rect 500658 172170 500754 172226
rect 500810 172170 500878 172226
rect 500934 172170 501002 172226
rect 501058 172170 501126 172226
rect 501182 172170 501278 172226
rect 500658 172102 501278 172170
rect 500658 172046 500754 172102
rect 500810 172046 500878 172102
rect 500934 172046 501002 172102
rect 501058 172046 501126 172102
rect 501182 172046 501278 172102
rect 500658 171978 501278 172046
rect 500658 171922 500754 171978
rect 500810 171922 500878 171978
rect 500934 171922 501002 171978
rect 501058 171922 501126 171978
rect 501182 171922 501278 171978
rect 500658 154350 501278 171922
rect 500658 154294 500754 154350
rect 500810 154294 500878 154350
rect 500934 154294 501002 154350
rect 501058 154294 501126 154350
rect 501182 154294 501278 154350
rect 500658 154226 501278 154294
rect 500658 154170 500754 154226
rect 500810 154170 500878 154226
rect 500934 154170 501002 154226
rect 501058 154170 501126 154226
rect 501182 154170 501278 154226
rect 500658 154102 501278 154170
rect 500658 154046 500754 154102
rect 500810 154046 500878 154102
rect 500934 154046 501002 154102
rect 501058 154046 501126 154102
rect 501182 154046 501278 154102
rect 500658 153978 501278 154046
rect 500658 153922 500754 153978
rect 500810 153922 500878 153978
rect 500934 153922 501002 153978
rect 501058 153922 501126 153978
rect 501182 153922 501278 153978
rect 500658 136350 501278 153922
rect 500658 136294 500754 136350
rect 500810 136294 500878 136350
rect 500934 136294 501002 136350
rect 501058 136294 501126 136350
rect 501182 136294 501278 136350
rect 500658 136226 501278 136294
rect 500658 136170 500754 136226
rect 500810 136170 500878 136226
rect 500934 136170 501002 136226
rect 501058 136170 501126 136226
rect 501182 136170 501278 136226
rect 500658 136102 501278 136170
rect 500658 136046 500754 136102
rect 500810 136046 500878 136102
rect 500934 136046 501002 136102
rect 501058 136046 501126 136102
rect 501182 136046 501278 136102
rect 500658 135978 501278 136046
rect 500658 135922 500754 135978
rect 500810 135922 500878 135978
rect 500934 135922 501002 135978
rect 501058 135922 501126 135978
rect 501182 135922 501278 135978
rect 500658 118350 501278 135922
rect 500658 118294 500754 118350
rect 500810 118294 500878 118350
rect 500934 118294 501002 118350
rect 501058 118294 501126 118350
rect 501182 118294 501278 118350
rect 500658 118226 501278 118294
rect 500658 118170 500754 118226
rect 500810 118170 500878 118226
rect 500934 118170 501002 118226
rect 501058 118170 501126 118226
rect 501182 118170 501278 118226
rect 500658 118102 501278 118170
rect 500658 118046 500754 118102
rect 500810 118046 500878 118102
rect 500934 118046 501002 118102
rect 501058 118046 501126 118102
rect 501182 118046 501278 118102
rect 500658 117978 501278 118046
rect 500658 117922 500754 117978
rect 500810 117922 500878 117978
rect 500934 117922 501002 117978
rect 501058 117922 501126 117978
rect 501182 117922 501278 117978
rect 500658 100350 501278 117922
rect 500658 100294 500754 100350
rect 500810 100294 500878 100350
rect 500934 100294 501002 100350
rect 501058 100294 501126 100350
rect 501182 100294 501278 100350
rect 500658 100226 501278 100294
rect 500658 100170 500754 100226
rect 500810 100170 500878 100226
rect 500934 100170 501002 100226
rect 501058 100170 501126 100226
rect 501182 100170 501278 100226
rect 500658 100102 501278 100170
rect 500658 100046 500754 100102
rect 500810 100046 500878 100102
rect 500934 100046 501002 100102
rect 501058 100046 501126 100102
rect 501182 100046 501278 100102
rect 500658 99978 501278 100046
rect 500658 99922 500754 99978
rect 500810 99922 500878 99978
rect 500934 99922 501002 99978
rect 501058 99922 501126 99978
rect 501182 99922 501278 99978
rect 500658 82350 501278 99922
rect 527658 597212 528278 598268
rect 527658 597156 527754 597212
rect 527810 597156 527878 597212
rect 527934 597156 528002 597212
rect 528058 597156 528126 597212
rect 528182 597156 528278 597212
rect 527658 597088 528278 597156
rect 527658 597032 527754 597088
rect 527810 597032 527878 597088
rect 527934 597032 528002 597088
rect 528058 597032 528126 597088
rect 528182 597032 528278 597088
rect 527658 596964 528278 597032
rect 527658 596908 527754 596964
rect 527810 596908 527878 596964
rect 527934 596908 528002 596964
rect 528058 596908 528126 596964
rect 528182 596908 528278 596964
rect 527658 596840 528278 596908
rect 527658 596784 527754 596840
rect 527810 596784 527878 596840
rect 527934 596784 528002 596840
rect 528058 596784 528126 596840
rect 528182 596784 528278 596840
rect 527658 580350 528278 596784
rect 527658 580294 527754 580350
rect 527810 580294 527878 580350
rect 527934 580294 528002 580350
rect 528058 580294 528126 580350
rect 528182 580294 528278 580350
rect 527658 580226 528278 580294
rect 527658 580170 527754 580226
rect 527810 580170 527878 580226
rect 527934 580170 528002 580226
rect 528058 580170 528126 580226
rect 528182 580170 528278 580226
rect 527658 580102 528278 580170
rect 527658 580046 527754 580102
rect 527810 580046 527878 580102
rect 527934 580046 528002 580102
rect 528058 580046 528126 580102
rect 528182 580046 528278 580102
rect 527658 579978 528278 580046
rect 527658 579922 527754 579978
rect 527810 579922 527878 579978
rect 527934 579922 528002 579978
rect 528058 579922 528126 579978
rect 528182 579922 528278 579978
rect 527658 562350 528278 579922
rect 527658 562294 527754 562350
rect 527810 562294 527878 562350
rect 527934 562294 528002 562350
rect 528058 562294 528126 562350
rect 528182 562294 528278 562350
rect 527658 562226 528278 562294
rect 527658 562170 527754 562226
rect 527810 562170 527878 562226
rect 527934 562170 528002 562226
rect 528058 562170 528126 562226
rect 528182 562170 528278 562226
rect 527658 562102 528278 562170
rect 527658 562046 527754 562102
rect 527810 562046 527878 562102
rect 527934 562046 528002 562102
rect 528058 562046 528126 562102
rect 528182 562046 528278 562102
rect 527658 561978 528278 562046
rect 527658 561922 527754 561978
rect 527810 561922 527878 561978
rect 527934 561922 528002 561978
rect 528058 561922 528126 561978
rect 528182 561922 528278 561978
rect 527658 544350 528278 561922
rect 527658 544294 527754 544350
rect 527810 544294 527878 544350
rect 527934 544294 528002 544350
rect 528058 544294 528126 544350
rect 528182 544294 528278 544350
rect 527658 544226 528278 544294
rect 527658 544170 527754 544226
rect 527810 544170 527878 544226
rect 527934 544170 528002 544226
rect 528058 544170 528126 544226
rect 528182 544170 528278 544226
rect 527658 544102 528278 544170
rect 527658 544046 527754 544102
rect 527810 544046 527878 544102
rect 527934 544046 528002 544102
rect 528058 544046 528126 544102
rect 528182 544046 528278 544102
rect 527658 543978 528278 544046
rect 527658 543922 527754 543978
rect 527810 543922 527878 543978
rect 527934 543922 528002 543978
rect 528058 543922 528126 543978
rect 528182 543922 528278 543978
rect 527658 526350 528278 543922
rect 527658 526294 527754 526350
rect 527810 526294 527878 526350
rect 527934 526294 528002 526350
rect 528058 526294 528126 526350
rect 528182 526294 528278 526350
rect 527658 526226 528278 526294
rect 527658 526170 527754 526226
rect 527810 526170 527878 526226
rect 527934 526170 528002 526226
rect 528058 526170 528126 526226
rect 528182 526170 528278 526226
rect 527658 526102 528278 526170
rect 527658 526046 527754 526102
rect 527810 526046 527878 526102
rect 527934 526046 528002 526102
rect 528058 526046 528126 526102
rect 528182 526046 528278 526102
rect 527658 525978 528278 526046
rect 527658 525922 527754 525978
rect 527810 525922 527878 525978
rect 527934 525922 528002 525978
rect 528058 525922 528126 525978
rect 528182 525922 528278 525978
rect 527658 508350 528278 525922
rect 527658 508294 527754 508350
rect 527810 508294 527878 508350
rect 527934 508294 528002 508350
rect 528058 508294 528126 508350
rect 528182 508294 528278 508350
rect 527658 508226 528278 508294
rect 527658 508170 527754 508226
rect 527810 508170 527878 508226
rect 527934 508170 528002 508226
rect 528058 508170 528126 508226
rect 528182 508170 528278 508226
rect 527658 508102 528278 508170
rect 527658 508046 527754 508102
rect 527810 508046 527878 508102
rect 527934 508046 528002 508102
rect 528058 508046 528126 508102
rect 528182 508046 528278 508102
rect 527658 507978 528278 508046
rect 527658 507922 527754 507978
rect 527810 507922 527878 507978
rect 527934 507922 528002 507978
rect 528058 507922 528126 507978
rect 528182 507922 528278 507978
rect 527658 490350 528278 507922
rect 527658 490294 527754 490350
rect 527810 490294 527878 490350
rect 527934 490294 528002 490350
rect 528058 490294 528126 490350
rect 528182 490294 528278 490350
rect 527658 490226 528278 490294
rect 527658 490170 527754 490226
rect 527810 490170 527878 490226
rect 527934 490170 528002 490226
rect 528058 490170 528126 490226
rect 528182 490170 528278 490226
rect 527658 490102 528278 490170
rect 527658 490046 527754 490102
rect 527810 490046 527878 490102
rect 527934 490046 528002 490102
rect 528058 490046 528126 490102
rect 528182 490046 528278 490102
rect 527658 489978 528278 490046
rect 527658 489922 527754 489978
rect 527810 489922 527878 489978
rect 527934 489922 528002 489978
rect 528058 489922 528126 489978
rect 528182 489922 528278 489978
rect 527658 472350 528278 489922
rect 527658 472294 527754 472350
rect 527810 472294 527878 472350
rect 527934 472294 528002 472350
rect 528058 472294 528126 472350
rect 528182 472294 528278 472350
rect 527658 472226 528278 472294
rect 527658 472170 527754 472226
rect 527810 472170 527878 472226
rect 527934 472170 528002 472226
rect 528058 472170 528126 472226
rect 528182 472170 528278 472226
rect 527658 472102 528278 472170
rect 527658 472046 527754 472102
rect 527810 472046 527878 472102
rect 527934 472046 528002 472102
rect 528058 472046 528126 472102
rect 528182 472046 528278 472102
rect 527658 471978 528278 472046
rect 527658 471922 527754 471978
rect 527810 471922 527878 471978
rect 527934 471922 528002 471978
rect 528058 471922 528126 471978
rect 528182 471922 528278 471978
rect 527658 454350 528278 471922
rect 527658 454294 527754 454350
rect 527810 454294 527878 454350
rect 527934 454294 528002 454350
rect 528058 454294 528126 454350
rect 528182 454294 528278 454350
rect 527658 454226 528278 454294
rect 527658 454170 527754 454226
rect 527810 454170 527878 454226
rect 527934 454170 528002 454226
rect 528058 454170 528126 454226
rect 528182 454170 528278 454226
rect 527658 454102 528278 454170
rect 527658 454046 527754 454102
rect 527810 454046 527878 454102
rect 527934 454046 528002 454102
rect 528058 454046 528126 454102
rect 528182 454046 528278 454102
rect 527658 453978 528278 454046
rect 527658 453922 527754 453978
rect 527810 453922 527878 453978
rect 527934 453922 528002 453978
rect 528058 453922 528126 453978
rect 528182 453922 528278 453978
rect 527658 436350 528278 453922
rect 527658 436294 527754 436350
rect 527810 436294 527878 436350
rect 527934 436294 528002 436350
rect 528058 436294 528126 436350
rect 528182 436294 528278 436350
rect 527658 436226 528278 436294
rect 527658 436170 527754 436226
rect 527810 436170 527878 436226
rect 527934 436170 528002 436226
rect 528058 436170 528126 436226
rect 528182 436170 528278 436226
rect 527658 436102 528278 436170
rect 527658 436046 527754 436102
rect 527810 436046 527878 436102
rect 527934 436046 528002 436102
rect 528058 436046 528126 436102
rect 528182 436046 528278 436102
rect 527658 435978 528278 436046
rect 527658 435922 527754 435978
rect 527810 435922 527878 435978
rect 527934 435922 528002 435978
rect 528058 435922 528126 435978
rect 528182 435922 528278 435978
rect 527658 418350 528278 435922
rect 527658 418294 527754 418350
rect 527810 418294 527878 418350
rect 527934 418294 528002 418350
rect 528058 418294 528126 418350
rect 528182 418294 528278 418350
rect 527658 418226 528278 418294
rect 527658 418170 527754 418226
rect 527810 418170 527878 418226
rect 527934 418170 528002 418226
rect 528058 418170 528126 418226
rect 528182 418170 528278 418226
rect 527658 418102 528278 418170
rect 527658 418046 527754 418102
rect 527810 418046 527878 418102
rect 527934 418046 528002 418102
rect 528058 418046 528126 418102
rect 528182 418046 528278 418102
rect 527658 417978 528278 418046
rect 527658 417922 527754 417978
rect 527810 417922 527878 417978
rect 527934 417922 528002 417978
rect 528058 417922 528126 417978
rect 528182 417922 528278 417978
rect 527658 400350 528278 417922
rect 527658 400294 527754 400350
rect 527810 400294 527878 400350
rect 527934 400294 528002 400350
rect 528058 400294 528126 400350
rect 528182 400294 528278 400350
rect 527658 400226 528278 400294
rect 527658 400170 527754 400226
rect 527810 400170 527878 400226
rect 527934 400170 528002 400226
rect 528058 400170 528126 400226
rect 528182 400170 528278 400226
rect 527658 400102 528278 400170
rect 527658 400046 527754 400102
rect 527810 400046 527878 400102
rect 527934 400046 528002 400102
rect 528058 400046 528126 400102
rect 528182 400046 528278 400102
rect 527658 399978 528278 400046
rect 527658 399922 527754 399978
rect 527810 399922 527878 399978
rect 527934 399922 528002 399978
rect 528058 399922 528126 399978
rect 528182 399922 528278 399978
rect 527658 382350 528278 399922
rect 527658 382294 527754 382350
rect 527810 382294 527878 382350
rect 527934 382294 528002 382350
rect 528058 382294 528126 382350
rect 528182 382294 528278 382350
rect 527658 382226 528278 382294
rect 527658 382170 527754 382226
rect 527810 382170 527878 382226
rect 527934 382170 528002 382226
rect 528058 382170 528126 382226
rect 528182 382170 528278 382226
rect 527658 382102 528278 382170
rect 527658 382046 527754 382102
rect 527810 382046 527878 382102
rect 527934 382046 528002 382102
rect 528058 382046 528126 382102
rect 528182 382046 528278 382102
rect 527658 381978 528278 382046
rect 527658 381922 527754 381978
rect 527810 381922 527878 381978
rect 527934 381922 528002 381978
rect 528058 381922 528126 381978
rect 528182 381922 528278 381978
rect 527658 364350 528278 381922
rect 527658 364294 527754 364350
rect 527810 364294 527878 364350
rect 527934 364294 528002 364350
rect 528058 364294 528126 364350
rect 528182 364294 528278 364350
rect 527658 364226 528278 364294
rect 527658 364170 527754 364226
rect 527810 364170 527878 364226
rect 527934 364170 528002 364226
rect 528058 364170 528126 364226
rect 528182 364170 528278 364226
rect 527658 364102 528278 364170
rect 527658 364046 527754 364102
rect 527810 364046 527878 364102
rect 527934 364046 528002 364102
rect 528058 364046 528126 364102
rect 528182 364046 528278 364102
rect 527658 363978 528278 364046
rect 527658 363922 527754 363978
rect 527810 363922 527878 363978
rect 527934 363922 528002 363978
rect 528058 363922 528126 363978
rect 528182 363922 528278 363978
rect 527658 346350 528278 363922
rect 527658 346294 527754 346350
rect 527810 346294 527878 346350
rect 527934 346294 528002 346350
rect 528058 346294 528126 346350
rect 528182 346294 528278 346350
rect 527658 346226 528278 346294
rect 527658 346170 527754 346226
rect 527810 346170 527878 346226
rect 527934 346170 528002 346226
rect 528058 346170 528126 346226
rect 528182 346170 528278 346226
rect 527658 346102 528278 346170
rect 527658 346046 527754 346102
rect 527810 346046 527878 346102
rect 527934 346046 528002 346102
rect 528058 346046 528126 346102
rect 528182 346046 528278 346102
rect 527658 345978 528278 346046
rect 527658 345922 527754 345978
rect 527810 345922 527878 345978
rect 527934 345922 528002 345978
rect 528058 345922 528126 345978
rect 528182 345922 528278 345978
rect 527658 328350 528278 345922
rect 527658 328294 527754 328350
rect 527810 328294 527878 328350
rect 527934 328294 528002 328350
rect 528058 328294 528126 328350
rect 528182 328294 528278 328350
rect 527658 328226 528278 328294
rect 527658 328170 527754 328226
rect 527810 328170 527878 328226
rect 527934 328170 528002 328226
rect 528058 328170 528126 328226
rect 528182 328170 528278 328226
rect 527658 328102 528278 328170
rect 527658 328046 527754 328102
rect 527810 328046 527878 328102
rect 527934 328046 528002 328102
rect 528058 328046 528126 328102
rect 528182 328046 528278 328102
rect 527658 327978 528278 328046
rect 527658 327922 527754 327978
rect 527810 327922 527878 327978
rect 527934 327922 528002 327978
rect 528058 327922 528126 327978
rect 528182 327922 528278 327978
rect 527658 310350 528278 327922
rect 527658 310294 527754 310350
rect 527810 310294 527878 310350
rect 527934 310294 528002 310350
rect 528058 310294 528126 310350
rect 528182 310294 528278 310350
rect 527658 310226 528278 310294
rect 527658 310170 527754 310226
rect 527810 310170 527878 310226
rect 527934 310170 528002 310226
rect 528058 310170 528126 310226
rect 528182 310170 528278 310226
rect 527658 310102 528278 310170
rect 527658 310046 527754 310102
rect 527810 310046 527878 310102
rect 527934 310046 528002 310102
rect 528058 310046 528126 310102
rect 528182 310046 528278 310102
rect 527658 309978 528278 310046
rect 527658 309922 527754 309978
rect 527810 309922 527878 309978
rect 527934 309922 528002 309978
rect 528058 309922 528126 309978
rect 528182 309922 528278 309978
rect 527658 292350 528278 309922
rect 527658 292294 527754 292350
rect 527810 292294 527878 292350
rect 527934 292294 528002 292350
rect 528058 292294 528126 292350
rect 528182 292294 528278 292350
rect 527658 292226 528278 292294
rect 527658 292170 527754 292226
rect 527810 292170 527878 292226
rect 527934 292170 528002 292226
rect 528058 292170 528126 292226
rect 528182 292170 528278 292226
rect 527658 292102 528278 292170
rect 527658 292046 527754 292102
rect 527810 292046 527878 292102
rect 527934 292046 528002 292102
rect 528058 292046 528126 292102
rect 528182 292046 528278 292102
rect 527658 291978 528278 292046
rect 527658 291922 527754 291978
rect 527810 291922 527878 291978
rect 527934 291922 528002 291978
rect 528058 291922 528126 291978
rect 528182 291922 528278 291978
rect 527658 274350 528278 291922
rect 527658 274294 527754 274350
rect 527810 274294 527878 274350
rect 527934 274294 528002 274350
rect 528058 274294 528126 274350
rect 528182 274294 528278 274350
rect 527658 274226 528278 274294
rect 527658 274170 527754 274226
rect 527810 274170 527878 274226
rect 527934 274170 528002 274226
rect 528058 274170 528126 274226
rect 528182 274170 528278 274226
rect 527658 274102 528278 274170
rect 527658 274046 527754 274102
rect 527810 274046 527878 274102
rect 527934 274046 528002 274102
rect 528058 274046 528126 274102
rect 528182 274046 528278 274102
rect 527658 273978 528278 274046
rect 527658 273922 527754 273978
rect 527810 273922 527878 273978
rect 527934 273922 528002 273978
rect 528058 273922 528126 273978
rect 528182 273922 528278 273978
rect 527658 256350 528278 273922
rect 527658 256294 527754 256350
rect 527810 256294 527878 256350
rect 527934 256294 528002 256350
rect 528058 256294 528126 256350
rect 528182 256294 528278 256350
rect 527658 256226 528278 256294
rect 527658 256170 527754 256226
rect 527810 256170 527878 256226
rect 527934 256170 528002 256226
rect 528058 256170 528126 256226
rect 528182 256170 528278 256226
rect 527658 256102 528278 256170
rect 527658 256046 527754 256102
rect 527810 256046 527878 256102
rect 527934 256046 528002 256102
rect 528058 256046 528126 256102
rect 528182 256046 528278 256102
rect 527658 255978 528278 256046
rect 527658 255922 527754 255978
rect 527810 255922 527878 255978
rect 527934 255922 528002 255978
rect 528058 255922 528126 255978
rect 528182 255922 528278 255978
rect 527658 238350 528278 255922
rect 527658 238294 527754 238350
rect 527810 238294 527878 238350
rect 527934 238294 528002 238350
rect 528058 238294 528126 238350
rect 528182 238294 528278 238350
rect 527658 238226 528278 238294
rect 527658 238170 527754 238226
rect 527810 238170 527878 238226
rect 527934 238170 528002 238226
rect 528058 238170 528126 238226
rect 528182 238170 528278 238226
rect 527658 238102 528278 238170
rect 527658 238046 527754 238102
rect 527810 238046 527878 238102
rect 527934 238046 528002 238102
rect 528058 238046 528126 238102
rect 528182 238046 528278 238102
rect 527658 237978 528278 238046
rect 527658 237922 527754 237978
rect 527810 237922 527878 237978
rect 527934 237922 528002 237978
rect 528058 237922 528126 237978
rect 528182 237922 528278 237978
rect 527658 220350 528278 237922
rect 527658 220294 527754 220350
rect 527810 220294 527878 220350
rect 527934 220294 528002 220350
rect 528058 220294 528126 220350
rect 528182 220294 528278 220350
rect 527658 220226 528278 220294
rect 527658 220170 527754 220226
rect 527810 220170 527878 220226
rect 527934 220170 528002 220226
rect 528058 220170 528126 220226
rect 528182 220170 528278 220226
rect 527658 220102 528278 220170
rect 527658 220046 527754 220102
rect 527810 220046 527878 220102
rect 527934 220046 528002 220102
rect 528058 220046 528126 220102
rect 528182 220046 528278 220102
rect 527658 219978 528278 220046
rect 527658 219922 527754 219978
rect 527810 219922 527878 219978
rect 527934 219922 528002 219978
rect 528058 219922 528126 219978
rect 528182 219922 528278 219978
rect 527658 202350 528278 219922
rect 527658 202294 527754 202350
rect 527810 202294 527878 202350
rect 527934 202294 528002 202350
rect 528058 202294 528126 202350
rect 528182 202294 528278 202350
rect 527658 202226 528278 202294
rect 527658 202170 527754 202226
rect 527810 202170 527878 202226
rect 527934 202170 528002 202226
rect 528058 202170 528126 202226
rect 528182 202170 528278 202226
rect 527658 202102 528278 202170
rect 527658 202046 527754 202102
rect 527810 202046 527878 202102
rect 527934 202046 528002 202102
rect 528058 202046 528126 202102
rect 528182 202046 528278 202102
rect 527658 201978 528278 202046
rect 527658 201922 527754 201978
rect 527810 201922 527878 201978
rect 527934 201922 528002 201978
rect 528058 201922 528126 201978
rect 528182 201922 528278 201978
rect 527658 184350 528278 201922
rect 527658 184294 527754 184350
rect 527810 184294 527878 184350
rect 527934 184294 528002 184350
rect 528058 184294 528126 184350
rect 528182 184294 528278 184350
rect 527658 184226 528278 184294
rect 527658 184170 527754 184226
rect 527810 184170 527878 184226
rect 527934 184170 528002 184226
rect 528058 184170 528126 184226
rect 528182 184170 528278 184226
rect 527658 184102 528278 184170
rect 527658 184046 527754 184102
rect 527810 184046 527878 184102
rect 527934 184046 528002 184102
rect 528058 184046 528126 184102
rect 528182 184046 528278 184102
rect 527658 183978 528278 184046
rect 527658 183922 527754 183978
rect 527810 183922 527878 183978
rect 527934 183922 528002 183978
rect 528058 183922 528126 183978
rect 528182 183922 528278 183978
rect 527658 166350 528278 183922
rect 527658 166294 527754 166350
rect 527810 166294 527878 166350
rect 527934 166294 528002 166350
rect 528058 166294 528126 166350
rect 528182 166294 528278 166350
rect 527658 166226 528278 166294
rect 527658 166170 527754 166226
rect 527810 166170 527878 166226
rect 527934 166170 528002 166226
rect 528058 166170 528126 166226
rect 528182 166170 528278 166226
rect 527658 166102 528278 166170
rect 527658 166046 527754 166102
rect 527810 166046 527878 166102
rect 527934 166046 528002 166102
rect 528058 166046 528126 166102
rect 528182 166046 528278 166102
rect 527658 165978 528278 166046
rect 527658 165922 527754 165978
rect 527810 165922 527878 165978
rect 527934 165922 528002 165978
rect 528058 165922 528126 165978
rect 528182 165922 528278 165978
rect 527658 148350 528278 165922
rect 527658 148294 527754 148350
rect 527810 148294 527878 148350
rect 527934 148294 528002 148350
rect 528058 148294 528126 148350
rect 528182 148294 528278 148350
rect 527658 148226 528278 148294
rect 527658 148170 527754 148226
rect 527810 148170 527878 148226
rect 527934 148170 528002 148226
rect 528058 148170 528126 148226
rect 528182 148170 528278 148226
rect 527658 148102 528278 148170
rect 527658 148046 527754 148102
rect 527810 148046 527878 148102
rect 527934 148046 528002 148102
rect 528058 148046 528126 148102
rect 528182 148046 528278 148102
rect 527658 147978 528278 148046
rect 527658 147922 527754 147978
rect 527810 147922 527878 147978
rect 527934 147922 528002 147978
rect 528058 147922 528126 147978
rect 528182 147922 528278 147978
rect 527658 130350 528278 147922
rect 527658 130294 527754 130350
rect 527810 130294 527878 130350
rect 527934 130294 528002 130350
rect 528058 130294 528126 130350
rect 528182 130294 528278 130350
rect 527658 130226 528278 130294
rect 527658 130170 527754 130226
rect 527810 130170 527878 130226
rect 527934 130170 528002 130226
rect 528058 130170 528126 130226
rect 528182 130170 528278 130226
rect 527658 130102 528278 130170
rect 527658 130046 527754 130102
rect 527810 130046 527878 130102
rect 527934 130046 528002 130102
rect 528058 130046 528126 130102
rect 528182 130046 528278 130102
rect 527658 129978 528278 130046
rect 527658 129922 527754 129978
rect 527810 129922 527878 129978
rect 527934 129922 528002 129978
rect 528058 129922 528126 129978
rect 528182 129922 528278 129978
rect 527658 112350 528278 129922
rect 527658 112294 527754 112350
rect 527810 112294 527878 112350
rect 527934 112294 528002 112350
rect 528058 112294 528126 112350
rect 528182 112294 528278 112350
rect 527658 112226 528278 112294
rect 527658 112170 527754 112226
rect 527810 112170 527878 112226
rect 527934 112170 528002 112226
rect 528058 112170 528126 112226
rect 528182 112170 528278 112226
rect 527658 112102 528278 112170
rect 527658 112046 527754 112102
rect 527810 112046 527878 112102
rect 527934 112046 528002 112102
rect 528058 112046 528126 112102
rect 528182 112046 528278 112102
rect 527658 111978 528278 112046
rect 527658 111922 527754 111978
rect 527810 111922 527878 111978
rect 527934 111922 528002 111978
rect 528058 111922 528126 111978
rect 528182 111922 528278 111978
rect 527658 94350 528278 111922
rect 527658 94294 527754 94350
rect 527810 94294 527878 94350
rect 527934 94294 528002 94350
rect 528058 94294 528126 94350
rect 528182 94294 528278 94350
rect 527658 94226 528278 94294
rect 527658 94170 527754 94226
rect 527810 94170 527878 94226
rect 527934 94170 528002 94226
rect 528058 94170 528126 94226
rect 528182 94170 528278 94226
rect 527658 94102 528278 94170
rect 527658 94046 527754 94102
rect 527810 94046 527878 94102
rect 527934 94046 528002 94102
rect 528058 94046 528126 94102
rect 528182 94046 528278 94102
rect 527658 93978 528278 94046
rect 527658 93922 527754 93978
rect 527810 93922 527878 93978
rect 527934 93922 528002 93978
rect 528058 93922 528126 93978
rect 528182 93922 528278 93978
rect 500658 82294 500754 82350
rect 500810 82294 500878 82350
rect 500934 82294 501002 82350
rect 501058 82294 501126 82350
rect 501182 82294 501278 82350
rect 500658 82226 501278 82294
rect 500658 82170 500754 82226
rect 500810 82170 500878 82226
rect 500934 82170 501002 82226
rect 501058 82170 501126 82226
rect 501182 82170 501278 82226
rect 500658 82102 501278 82170
rect 500658 82046 500754 82102
rect 500810 82046 500878 82102
rect 500934 82046 501002 82102
rect 501058 82046 501126 82102
rect 501182 82046 501278 82102
rect 500658 81978 501278 82046
rect 500658 81922 500754 81978
rect 500810 81922 500878 81978
rect 500934 81922 501002 81978
rect 501058 81922 501126 81978
rect 501182 81922 501278 81978
rect 496938 76294 497034 76350
rect 497090 76294 497158 76350
rect 497214 76294 497282 76350
rect 497338 76294 497406 76350
rect 497462 76294 497558 76350
rect 496938 76226 497558 76294
rect 496938 76170 497034 76226
rect 497090 76170 497158 76226
rect 497214 76170 497282 76226
rect 497338 76170 497406 76226
rect 497462 76170 497558 76226
rect 496938 76102 497558 76170
rect 496938 76046 497034 76102
rect 497090 76046 497158 76102
rect 497214 76046 497282 76102
rect 497338 76046 497406 76102
rect 497462 76046 497558 76102
rect 496938 75978 497558 76046
rect 496938 75922 497034 75978
rect 497090 75922 497158 75978
rect 497214 75922 497282 75978
rect 497338 75922 497406 75978
rect 497462 75922 497558 75978
rect 480508 4162 480564 4172
rect 482188 60778 482244 60788
rect 482188 4228 482244 60722
rect 496938 58350 497558 75922
rect 496938 58294 497034 58350
rect 497090 58294 497158 58350
rect 497214 58294 497282 58350
rect 497338 58294 497406 58350
rect 497462 58294 497558 58350
rect 496938 58226 497558 58294
rect 496938 58170 497034 58226
rect 497090 58170 497158 58226
rect 497214 58170 497282 58226
rect 497338 58170 497406 58226
rect 497462 58170 497558 58226
rect 496938 58102 497558 58170
rect 496938 58046 497034 58102
rect 497090 58046 497158 58102
rect 497214 58046 497282 58102
rect 497338 58046 497406 58102
rect 497462 58046 497558 58102
rect 496938 57978 497558 58046
rect 496938 57922 497034 57978
rect 497090 57922 497158 57978
rect 497214 57922 497282 57978
rect 497338 57922 497406 57978
rect 497462 57922 497558 57978
rect 487228 54298 487284 54308
rect 487228 20188 487284 54242
rect 488908 47278 488964 47288
rect 487228 20132 487396 20188
rect 482188 4162 482244 4172
rect 487340 4228 487396 20132
rect 487340 4162 487396 4172
rect 488908 4228 488964 47222
rect 496938 40350 497558 57922
rect 496938 40294 497034 40350
rect 497090 40294 497158 40350
rect 497214 40294 497282 40350
rect 497338 40294 497406 40350
rect 497462 40294 497558 40350
rect 496938 40226 497558 40294
rect 496938 40170 497034 40226
rect 497090 40170 497158 40226
rect 497214 40170 497282 40226
rect 497338 40170 497406 40226
rect 497462 40170 497558 40226
rect 496938 40102 497558 40170
rect 496938 40046 497034 40102
rect 497090 40046 497158 40102
rect 497214 40046 497282 40102
rect 497338 40046 497406 40102
rect 497462 40046 497558 40102
rect 496938 39978 497558 40046
rect 496938 39922 497034 39978
rect 497090 39922 497158 39978
rect 497214 39922 497282 39978
rect 497338 39922 497406 39978
rect 497462 39922 497558 39978
rect 488908 4162 488964 4172
rect 492268 38818 492324 38828
rect 492268 4228 492324 38762
rect 492268 4162 492324 4172
rect 493948 30358 494004 30368
rect 493948 4228 494004 30302
rect 496938 22350 497558 39922
rect 496938 22294 497034 22350
rect 497090 22294 497158 22350
rect 497214 22294 497282 22350
rect 497338 22294 497406 22350
rect 497462 22294 497558 22350
rect 496938 22226 497558 22294
rect 496938 22170 497034 22226
rect 497090 22170 497158 22226
rect 497214 22170 497282 22226
rect 497338 22170 497406 22226
rect 497462 22170 497558 22226
rect 496938 22102 497558 22170
rect 496938 22046 497034 22102
rect 497090 22046 497158 22102
rect 497214 22046 497282 22102
rect 497338 22046 497406 22102
rect 497462 22046 497558 22102
rect 496938 21978 497558 22046
rect 496938 21922 497034 21978
rect 497090 21922 497158 21978
rect 497214 21922 497282 21978
rect 497338 21922 497406 21978
rect 497462 21922 497558 21978
rect 493948 4162 494004 4172
rect 495628 11818 495684 11828
rect 495628 4228 495684 11762
rect 495628 4162 495684 4172
rect 496938 4350 497558 21922
rect 496938 4294 497034 4350
rect 497090 4294 497158 4350
rect 497214 4294 497282 4350
rect 497338 4294 497406 4350
rect 497462 4294 497558 4350
rect 496938 4226 497558 4294
rect 496938 4170 497034 4226
rect 497090 4170 497158 4226
rect 497214 4170 497282 4226
rect 497338 4170 497406 4226
rect 497462 4170 497558 4226
rect 469938 -1176 470034 -1120
rect 470090 -1176 470158 -1120
rect 470214 -1176 470282 -1120
rect 470338 -1176 470406 -1120
rect 470462 -1176 470558 -1120
rect 469938 -1244 470558 -1176
rect 469938 -1300 470034 -1244
rect 470090 -1300 470158 -1244
rect 470214 -1300 470282 -1244
rect 470338 -1300 470406 -1244
rect 470462 -1300 470558 -1244
rect 469938 -1368 470558 -1300
rect 469938 -1424 470034 -1368
rect 470090 -1424 470158 -1368
rect 470214 -1424 470282 -1368
rect 470338 -1424 470406 -1368
rect 470462 -1424 470558 -1368
rect 469938 -1492 470558 -1424
rect 469938 -1548 470034 -1492
rect 470090 -1548 470158 -1492
rect 470214 -1548 470282 -1492
rect 470338 -1548 470406 -1492
rect 470462 -1548 470558 -1492
rect 469938 -1644 470558 -1548
rect 496938 4102 497558 4170
rect 497644 77338 497700 77348
rect 497644 4228 497700 77282
rect 497644 4162 497700 4172
rect 500658 64350 501278 81922
rect 500658 64294 500754 64350
rect 500810 64294 500878 64350
rect 500934 64294 501002 64350
rect 501058 64294 501126 64350
rect 501182 64294 501278 64350
rect 500658 64226 501278 64294
rect 500658 64170 500754 64226
rect 500810 64170 500878 64226
rect 500934 64170 501002 64226
rect 501058 64170 501126 64226
rect 501182 64170 501278 64226
rect 500658 64102 501278 64170
rect 500658 64046 500754 64102
rect 500810 64046 500878 64102
rect 500934 64046 501002 64102
rect 501058 64046 501126 64102
rect 501182 64046 501278 64102
rect 500658 63978 501278 64046
rect 500658 63922 500754 63978
rect 500810 63922 500878 63978
rect 500934 63922 501002 63978
rect 501058 63922 501126 63978
rect 501182 63922 501278 63978
rect 500658 46350 501278 63922
rect 500658 46294 500754 46350
rect 500810 46294 500878 46350
rect 500934 46294 501002 46350
rect 501058 46294 501126 46350
rect 501182 46294 501278 46350
rect 500658 46226 501278 46294
rect 500658 46170 500754 46226
rect 500810 46170 500878 46226
rect 500934 46170 501002 46226
rect 501058 46170 501126 46226
rect 501182 46170 501278 46226
rect 500658 46102 501278 46170
rect 500658 46046 500754 46102
rect 500810 46046 500878 46102
rect 500934 46046 501002 46102
rect 501058 46046 501126 46102
rect 501182 46046 501278 46102
rect 500658 45978 501278 46046
rect 500658 45922 500754 45978
rect 500810 45922 500878 45978
rect 500934 45922 501002 45978
rect 501058 45922 501126 45978
rect 501182 45922 501278 45978
rect 500658 28350 501278 45922
rect 504812 86436 504868 86446
rect 504812 32788 504868 86380
rect 527658 76350 528278 93922
rect 527658 76294 527754 76350
rect 527810 76294 527878 76350
rect 527934 76294 528002 76350
rect 528058 76294 528126 76350
rect 528182 76294 528278 76350
rect 527658 76226 528278 76294
rect 527658 76170 527754 76226
rect 527810 76170 527878 76226
rect 527934 76170 528002 76226
rect 528058 76170 528126 76226
rect 528182 76170 528278 76226
rect 527658 76102 528278 76170
rect 527658 76046 527754 76102
rect 527810 76046 527878 76102
rect 527934 76046 528002 76102
rect 528058 76046 528126 76102
rect 528182 76046 528278 76102
rect 527658 75978 528278 76046
rect 527658 75922 527754 75978
rect 527810 75922 527878 75978
rect 527934 75922 528002 75978
rect 528058 75922 528126 75978
rect 528182 75922 528278 75978
rect 525868 62218 525924 62228
rect 515788 60598 515844 60608
rect 509068 57358 509124 57368
rect 504812 32722 504868 32732
rect 505708 35398 505764 35408
rect 500658 28294 500754 28350
rect 500810 28294 500878 28350
rect 500934 28294 501002 28350
rect 501058 28294 501126 28350
rect 501182 28294 501278 28350
rect 500658 28226 501278 28294
rect 500658 28170 500754 28226
rect 500810 28170 500878 28226
rect 500934 28170 501002 28226
rect 501058 28170 501126 28226
rect 501182 28170 501278 28226
rect 500658 28102 501278 28170
rect 500658 28046 500754 28102
rect 500810 28046 500878 28102
rect 500934 28046 501002 28102
rect 501058 28046 501126 28102
rect 501182 28046 501278 28102
rect 500658 27978 501278 28046
rect 500658 27922 500754 27978
rect 500810 27922 500878 27978
rect 500934 27922 501002 27978
rect 501058 27922 501126 27978
rect 501182 27922 501278 27978
rect 500658 10350 501278 27922
rect 500658 10294 500754 10350
rect 500810 10294 500878 10350
rect 500934 10294 501002 10350
rect 501058 10294 501126 10350
rect 501182 10294 501278 10350
rect 500658 10226 501278 10294
rect 500658 10170 500754 10226
rect 500810 10170 500878 10226
rect 500934 10170 501002 10226
rect 501058 10170 501126 10226
rect 501182 10170 501278 10226
rect 500658 10102 501278 10170
rect 500658 10046 500754 10102
rect 500810 10046 500878 10102
rect 500934 10046 501002 10102
rect 501058 10046 501126 10102
rect 501182 10046 501278 10102
rect 500658 9978 501278 10046
rect 500658 9922 500754 9978
rect 500810 9922 500878 9978
rect 500934 9922 501002 9978
rect 501058 9922 501126 9978
rect 501182 9922 501278 9978
rect 496938 4046 497034 4102
rect 497090 4046 497158 4102
rect 497214 4046 497282 4102
rect 497338 4046 497406 4102
rect 497462 4046 497558 4102
rect 496938 3978 497558 4046
rect 496938 3922 497034 3978
rect 497090 3922 497158 3978
rect 497214 3922 497282 3978
rect 497338 3922 497406 3978
rect 497462 3922 497558 3978
rect 496938 -160 497558 3922
rect 496938 -216 497034 -160
rect 497090 -216 497158 -160
rect 497214 -216 497282 -160
rect 497338 -216 497406 -160
rect 497462 -216 497558 -160
rect 496938 -284 497558 -216
rect 496938 -340 497034 -284
rect 497090 -340 497158 -284
rect 497214 -340 497282 -284
rect 497338 -340 497406 -284
rect 497462 -340 497558 -284
rect 496938 -408 497558 -340
rect 496938 -464 497034 -408
rect 497090 -464 497158 -408
rect 497214 -464 497282 -408
rect 497338 -464 497406 -408
rect 497462 -464 497558 -408
rect 496938 -532 497558 -464
rect 496938 -588 497034 -532
rect 497090 -588 497158 -532
rect 497214 -588 497282 -532
rect 497338 -588 497406 -532
rect 497462 -588 497558 -532
rect 496938 -1644 497558 -588
rect 500658 -1120 501278 9922
rect 501340 28738 501396 28748
rect 501340 4228 501396 28682
rect 501340 4162 501396 4172
rect 504028 16858 504084 16868
rect 504028 4228 504084 16802
rect 504028 4162 504084 4172
rect 505708 4228 505764 35342
rect 505708 4162 505764 4172
rect 508284 10738 508340 10748
rect 508284 4228 508340 10682
rect 508284 4162 508340 4172
rect 509068 4228 509124 57302
rect 509068 4162 509124 4172
rect 510748 54118 510804 54128
rect 510748 4228 510804 54062
rect 515788 20188 515844 60542
rect 520828 58978 520884 58988
rect 517468 52318 517524 52328
rect 515788 20132 515956 20188
rect 510748 4162 510804 4172
rect 515900 4228 515956 20132
rect 515900 4162 515956 4172
rect 517468 4228 517524 52262
rect 517468 4162 517524 4172
rect 520828 4228 520884 58922
rect 520828 4162 520884 4172
rect 522508 55738 522564 55748
rect 522508 4228 522564 55682
rect 522508 4162 522564 4172
rect 525868 4228 525924 62162
rect 525868 4162 525924 4172
rect 527658 58350 528278 75922
rect 527658 58294 527754 58350
rect 527810 58294 527878 58350
rect 527934 58294 528002 58350
rect 528058 58294 528126 58350
rect 528182 58294 528278 58350
rect 527658 58226 528278 58294
rect 527658 58170 527754 58226
rect 527810 58170 527878 58226
rect 527934 58170 528002 58226
rect 528058 58170 528126 58226
rect 528182 58170 528278 58226
rect 527658 58102 528278 58170
rect 527658 58046 527754 58102
rect 527810 58046 527878 58102
rect 527934 58046 528002 58102
rect 528058 58046 528126 58102
rect 528182 58046 528278 58102
rect 527658 57978 528278 58046
rect 527658 57922 527754 57978
rect 527810 57922 527878 57978
rect 527934 57922 528002 57978
rect 528058 57922 528126 57978
rect 528182 57922 528278 57978
rect 527658 40350 528278 57922
rect 527658 40294 527754 40350
rect 527810 40294 527878 40350
rect 527934 40294 528002 40350
rect 528058 40294 528126 40350
rect 528182 40294 528278 40350
rect 527658 40226 528278 40294
rect 527658 40170 527754 40226
rect 527810 40170 527878 40226
rect 527934 40170 528002 40226
rect 528058 40170 528126 40226
rect 528182 40170 528278 40226
rect 527658 40102 528278 40170
rect 527658 40046 527754 40102
rect 527810 40046 527878 40102
rect 527934 40046 528002 40102
rect 528058 40046 528126 40102
rect 528182 40046 528278 40102
rect 527658 39978 528278 40046
rect 527658 39922 527754 39978
rect 527810 39922 527878 39978
rect 527934 39922 528002 39978
rect 528058 39922 528126 39978
rect 528182 39922 528278 39978
rect 527658 22350 528278 39922
rect 527658 22294 527754 22350
rect 527810 22294 527878 22350
rect 527934 22294 528002 22350
rect 528058 22294 528126 22350
rect 528182 22294 528278 22350
rect 527658 22226 528278 22294
rect 527658 22170 527754 22226
rect 527810 22170 527878 22226
rect 527934 22170 528002 22226
rect 528058 22170 528126 22226
rect 528182 22170 528278 22226
rect 527658 22102 528278 22170
rect 527658 22046 527754 22102
rect 527810 22046 527878 22102
rect 527934 22046 528002 22102
rect 528058 22046 528126 22102
rect 528182 22046 528278 22102
rect 527658 21978 528278 22046
rect 527658 21922 527754 21978
rect 527810 21922 527878 21978
rect 527934 21922 528002 21978
rect 528058 21922 528126 21978
rect 528182 21922 528278 21978
rect 527658 4350 528278 21922
rect 531378 598172 531998 598268
rect 531378 598116 531474 598172
rect 531530 598116 531598 598172
rect 531654 598116 531722 598172
rect 531778 598116 531846 598172
rect 531902 598116 531998 598172
rect 531378 598048 531998 598116
rect 531378 597992 531474 598048
rect 531530 597992 531598 598048
rect 531654 597992 531722 598048
rect 531778 597992 531846 598048
rect 531902 597992 531998 598048
rect 531378 597924 531998 597992
rect 531378 597868 531474 597924
rect 531530 597868 531598 597924
rect 531654 597868 531722 597924
rect 531778 597868 531846 597924
rect 531902 597868 531998 597924
rect 531378 597800 531998 597868
rect 531378 597744 531474 597800
rect 531530 597744 531598 597800
rect 531654 597744 531722 597800
rect 531778 597744 531846 597800
rect 531902 597744 531998 597800
rect 531378 586350 531998 597744
rect 531378 586294 531474 586350
rect 531530 586294 531598 586350
rect 531654 586294 531722 586350
rect 531778 586294 531846 586350
rect 531902 586294 531998 586350
rect 531378 586226 531998 586294
rect 531378 586170 531474 586226
rect 531530 586170 531598 586226
rect 531654 586170 531722 586226
rect 531778 586170 531846 586226
rect 531902 586170 531998 586226
rect 531378 586102 531998 586170
rect 531378 586046 531474 586102
rect 531530 586046 531598 586102
rect 531654 586046 531722 586102
rect 531778 586046 531846 586102
rect 531902 586046 531998 586102
rect 531378 585978 531998 586046
rect 531378 585922 531474 585978
rect 531530 585922 531598 585978
rect 531654 585922 531722 585978
rect 531778 585922 531846 585978
rect 531902 585922 531998 585978
rect 531378 568350 531998 585922
rect 531378 568294 531474 568350
rect 531530 568294 531598 568350
rect 531654 568294 531722 568350
rect 531778 568294 531846 568350
rect 531902 568294 531998 568350
rect 531378 568226 531998 568294
rect 531378 568170 531474 568226
rect 531530 568170 531598 568226
rect 531654 568170 531722 568226
rect 531778 568170 531846 568226
rect 531902 568170 531998 568226
rect 531378 568102 531998 568170
rect 531378 568046 531474 568102
rect 531530 568046 531598 568102
rect 531654 568046 531722 568102
rect 531778 568046 531846 568102
rect 531902 568046 531998 568102
rect 531378 567978 531998 568046
rect 531378 567922 531474 567978
rect 531530 567922 531598 567978
rect 531654 567922 531722 567978
rect 531778 567922 531846 567978
rect 531902 567922 531998 567978
rect 531378 550350 531998 567922
rect 531378 550294 531474 550350
rect 531530 550294 531598 550350
rect 531654 550294 531722 550350
rect 531778 550294 531846 550350
rect 531902 550294 531998 550350
rect 531378 550226 531998 550294
rect 531378 550170 531474 550226
rect 531530 550170 531598 550226
rect 531654 550170 531722 550226
rect 531778 550170 531846 550226
rect 531902 550170 531998 550226
rect 531378 550102 531998 550170
rect 531378 550046 531474 550102
rect 531530 550046 531598 550102
rect 531654 550046 531722 550102
rect 531778 550046 531846 550102
rect 531902 550046 531998 550102
rect 531378 549978 531998 550046
rect 531378 549922 531474 549978
rect 531530 549922 531598 549978
rect 531654 549922 531722 549978
rect 531778 549922 531846 549978
rect 531902 549922 531998 549978
rect 531378 532350 531998 549922
rect 531378 532294 531474 532350
rect 531530 532294 531598 532350
rect 531654 532294 531722 532350
rect 531778 532294 531846 532350
rect 531902 532294 531998 532350
rect 531378 532226 531998 532294
rect 531378 532170 531474 532226
rect 531530 532170 531598 532226
rect 531654 532170 531722 532226
rect 531778 532170 531846 532226
rect 531902 532170 531998 532226
rect 531378 532102 531998 532170
rect 531378 532046 531474 532102
rect 531530 532046 531598 532102
rect 531654 532046 531722 532102
rect 531778 532046 531846 532102
rect 531902 532046 531998 532102
rect 531378 531978 531998 532046
rect 531378 531922 531474 531978
rect 531530 531922 531598 531978
rect 531654 531922 531722 531978
rect 531778 531922 531846 531978
rect 531902 531922 531998 531978
rect 531378 514350 531998 531922
rect 531378 514294 531474 514350
rect 531530 514294 531598 514350
rect 531654 514294 531722 514350
rect 531778 514294 531846 514350
rect 531902 514294 531998 514350
rect 531378 514226 531998 514294
rect 531378 514170 531474 514226
rect 531530 514170 531598 514226
rect 531654 514170 531722 514226
rect 531778 514170 531846 514226
rect 531902 514170 531998 514226
rect 531378 514102 531998 514170
rect 531378 514046 531474 514102
rect 531530 514046 531598 514102
rect 531654 514046 531722 514102
rect 531778 514046 531846 514102
rect 531902 514046 531998 514102
rect 531378 513978 531998 514046
rect 531378 513922 531474 513978
rect 531530 513922 531598 513978
rect 531654 513922 531722 513978
rect 531778 513922 531846 513978
rect 531902 513922 531998 513978
rect 531378 496350 531998 513922
rect 531378 496294 531474 496350
rect 531530 496294 531598 496350
rect 531654 496294 531722 496350
rect 531778 496294 531846 496350
rect 531902 496294 531998 496350
rect 531378 496226 531998 496294
rect 531378 496170 531474 496226
rect 531530 496170 531598 496226
rect 531654 496170 531722 496226
rect 531778 496170 531846 496226
rect 531902 496170 531998 496226
rect 531378 496102 531998 496170
rect 531378 496046 531474 496102
rect 531530 496046 531598 496102
rect 531654 496046 531722 496102
rect 531778 496046 531846 496102
rect 531902 496046 531998 496102
rect 531378 495978 531998 496046
rect 531378 495922 531474 495978
rect 531530 495922 531598 495978
rect 531654 495922 531722 495978
rect 531778 495922 531846 495978
rect 531902 495922 531998 495978
rect 531378 478350 531998 495922
rect 531378 478294 531474 478350
rect 531530 478294 531598 478350
rect 531654 478294 531722 478350
rect 531778 478294 531846 478350
rect 531902 478294 531998 478350
rect 531378 478226 531998 478294
rect 531378 478170 531474 478226
rect 531530 478170 531598 478226
rect 531654 478170 531722 478226
rect 531778 478170 531846 478226
rect 531902 478170 531998 478226
rect 531378 478102 531998 478170
rect 531378 478046 531474 478102
rect 531530 478046 531598 478102
rect 531654 478046 531722 478102
rect 531778 478046 531846 478102
rect 531902 478046 531998 478102
rect 531378 477978 531998 478046
rect 531378 477922 531474 477978
rect 531530 477922 531598 477978
rect 531654 477922 531722 477978
rect 531778 477922 531846 477978
rect 531902 477922 531998 477978
rect 531378 460350 531998 477922
rect 531378 460294 531474 460350
rect 531530 460294 531598 460350
rect 531654 460294 531722 460350
rect 531778 460294 531846 460350
rect 531902 460294 531998 460350
rect 531378 460226 531998 460294
rect 531378 460170 531474 460226
rect 531530 460170 531598 460226
rect 531654 460170 531722 460226
rect 531778 460170 531846 460226
rect 531902 460170 531998 460226
rect 531378 460102 531998 460170
rect 531378 460046 531474 460102
rect 531530 460046 531598 460102
rect 531654 460046 531722 460102
rect 531778 460046 531846 460102
rect 531902 460046 531998 460102
rect 531378 459978 531998 460046
rect 531378 459922 531474 459978
rect 531530 459922 531598 459978
rect 531654 459922 531722 459978
rect 531778 459922 531846 459978
rect 531902 459922 531998 459978
rect 531378 442350 531998 459922
rect 531378 442294 531474 442350
rect 531530 442294 531598 442350
rect 531654 442294 531722 442350
rect 531778 442294 531846 442350
rect 531902 442294 531998 442350
rect 531378 442226 531998 442294
rect 531378 442170 531474 442226
rect 531530 442170 531598 442226
rect 531654 442170 531722 442226
rect 531778 442170 531846 442226
rect 531902 442170 531998 442226
rect 531378 442102 531998 442170
rect 531378 442046 531474 442102
rect 531530 442046 531598 442102
rect 531654 442046 531722 442102
rect 531778 442046 531846 442102
rect 531902 442046 531998 442102
rect 531378 441978 531998 442046
rect 531378 441922 531474 441978
rect 531530 441922 531598 441978
rect 531654 441922 531722 441978
rect 531778 441922 531846 441978
rect 531902 441922 531998 441978
rect 531378 424350 531998 441922
rect 531378 424294 531474 424350
rect 531530 424294 531598 424350
rect 531654 424294 531722 424350
rect 531778 424294 531846 424350
rect 531902 424294 531998 424350
rect 531378 424226 531998 424294
rect 531378 424170 531474 424226
rect 531530 424170 531598 424226
rect 531654 424170 531722 424226
rect 531778 424170 531846 424226
rect 531902 424170 531998 424226
rect 531378 424102 531998 424170
rect 531378 424046 531474 424102
rect 531530 424046 531598 424102
rect 531654 424046 531722 424102
rect 531778 424046 531846 424102
rect 531902 424046 531998 424102
rect 531378 423978 531998 424046
rect 531378 423922 531474 423978
rect 531530 423922 531598 423978
rect 531654 423922 531722 423978
rect 531778 423922 531846 423978
rect 531902 423922 531998 423978
rect 531378 406350 531998 423922
rect 531378 406294 531474 406350
rect 531530 406294 531598 406350
rect 531654 406294 531722 406350
rect 531778 406294 531846 406350
rect 531902 406294 531998 406350
rect 531378 406226 531998 406294
rect 531378 406170 531474 406226
rect 531530 406170 531598 406226
rect 531654 406170 531722 406226
rect 531778 406170 531846 406226
rect 531902 406170 531998 406226
rect 531378 406102 531998 406170
rect 531378 406046 531474 406102
rect 531530 406046 531598 406102
rect 531654 406046 531722 406102
rect 531778 406046 531846 406102
rect 531902 406046 531998 406102
rect 531378 405978 531998 406046
rect 531378 405922 531474 405978
rect 531530 405922 531598 405978
rect 531654 405922 531722 405978
rect 531778 405922 531846 405978
rect 531902 405922 531998 405978
rect 531378 388350 531998 405922
rect 531378 388294 531474 388350
rect 531530 388294 531598 388350
rect 531654 388294 531722 388350
rect 531778 388294 531846 388350
rect 531902 388294 531998 388350
rect 531378 388226 531998 388294
rect 531378 388170 531474 388226
rect 531530 388170 531598 388226
rect 531654 388170 531722 388226
rect 531778 388170 531846 388226
rect 531902 388170 531998 388226
rect 531378 388102 531998 388170
rect 531378 388046 531474 388102
rect 531530 388046 531598 388102
rect 531654 388046 531722 388102
rect 531778 388046 531846 388102
rect 531902 388046 531998 388102
rect 531378 387978 531998 388046
rect 531378 387922 531474 387978
rect 531530 387922 531598 387978
rect 531654 387922 531722 387978
rect 531778 387922 531846 387978
rect 531902 387922 531998 387978
rect 531378 370350 531998 387922
rect 531378 370294 531474 370350
rect 531530 370294 531598 370350
rect 531654 370294 531722 370350
rect 531778 370294 531846 370350
rect 531902 370294 531998 370350
rect 531378 370226 531998 370294
rect 531378 370170 531474 370226
rect 531530 370170 531598 370226
rect 531654 370170 531722 370226
rect 531778 370170 531846 370226
rect 531902 370170 531998 370226
rect 531378 370102 531998 370170
rect 531378 370046 531474 370102
rect 531530 370046 531598 370102
rect 531654 370046 531722 370102
rect 531778 370046 531846 370102
rect 531902 370046 531998 370102
rect 531378 369978 531998 370046
rect 531378 369922 531474 369978
rect 531530 369922 531598 369978
rect 531654 369922 531722 369978
rect 531778 369922 531846 369978
rect 531902 369922 531998 369978
rect 531378 352350 531998 369922
rect 531378 352294 531474 352350
rect 531530 352294 531598 352350
rect 531654 352294 531722 352350
rect 531778 352294 531846 352350
rect 531902 352294 531998 352350
rect 531378 352226 531998 352294
rect 531378 352170 531474 352226
rect 531530 352170 531598 352226
rect 531654 352170 531722 352226
rect 531778 352170 531846 352226
rect 531902 352170 531998 352226
rect 531378 352102 531998 352170
rect 531378 352046 531474 352102
rect 531530 352046 531598 352102
rect 531654 352046 531722 352102
rect 531778 352046 531846 352102
rect 531902 352046 531998 352102
rect 531378 351978 531998 352046
rect 531378 351922 531474 351978
rect 531530 351922 531598 351978
rect 531654 351922 531722 351978
rect 531778 351922 531846 351978
rect 531902 351922 531998 351978
rect 531378 334350 531998 351922
rect 531378 334294 531474 334350
rect 531530 334294 531598 334350
rect 531654 334294 531722 334350
rect 531778 334294 531846 334350
rect 531902 334294 531998 334350
rect 531378 334226 531998 334294
rect 531378 334170 531474 334226
rect 531530 334170 531598 334226
rect 531654 334170 531722 334226
rect 531778 334170 531846 334226
rect 531902 334170 531998 334226
rect 531378 334102 531998 334170
rect 531378 334046 531474 334102
rect 531530 334046 531598 334102
rect 531654 334046 531722 334102
rect 531778 334046 531846 334102
rect 531902 334046 531998 334102
rect 531378 333978 531998 334046
rect 531378 333922 531474 333978
rect 531530 333922 531598 333978
rect 531654 333922 531722 333978
rect 531778 333922 531846 333978
rect 531902 333922 531998 333978
rect 531378 316350 531998 333922
rect 531378 316294 531474 316350
rect 531530 316294 531598 316350
rect 531654 316294 531722 316350
rect 531778 316294 531846 316350
rect 531902 316294 531998 316350
rect 531378 316226 531998 316294
rect 531378 316170 531474 316226
rect 531530 316170 531598 316226
rect 531654 316170 531722 316226
rect 531778 316170 531846 316226
rect 531902 316170 531998 316226
rect 531378 316102 531998 316170
rect 531378 316046 531474 316102
rect 531530 316046 531598 316102
rect 531654 316046 531722 316102
rect 531778 316046 531846 316102
rect 531902 316046 531998 316102
rect 531378 315978 531998 316046
rect 531378 315922 531474 315978
rect 531530 315922 531598 315978
rect 531654 315922 531722 315978
rect 531778 315922 531846 315978
rect 531902 315922 531998 315978
rect 531378 298350 531998 315922
rect 531378 298294 531474 298350
rect 531530 298294 531598 298350
rect 531654 298294 531722 298350
rect 531778 298294 531846 298350
rect 531902 298294 531998 298350
rect 531378 298226 531998 298294
rect 531378 298170 531474 298226
rect 531530 298170 531598 298226
rect 531654 298170 531722 298226
rect 531778 298170 531846 298226
rect 531902 298170 531998 298226
rect 531378 298102 531998 298170
rect 531378 298046 531474 298102
rect 531530 298046 531598 298102
rect 531654 298046 531722 298102
rect 531778 298046 531846 298102
rect 531902 298046 531998 298102
rect 531378 297978 531998 298046
rect 531378 297922 531474 297978
rect 531530 297922 531598 297978
rect 531654 297922 531722 297978
rect 531778 297922 531846 297978
rect 531902 297922 531998 297978
rect 531378 280350 531998 297922
rect 531378 280294 531474 280350
rect 531530 280294 531598 280350
rect 531654 280294 531722 280350
rect 531778 280294 531846 280350
rect 531902 280294 531998 280350
rect 531378 280226 531998 280294
rect 531378 280170 531474 280226
rect 531530 280170 531598 280226
rect 531654 280170 531722 280226
rect 531778 280170 531846 280226
rect 531902 280170 531998 280226
rect 531378 280102 531998 280170
rect 531378 280046 531474 280102
rect 531530 280046 531598 280102
rect 531654 280046 531722 280102
rect 531778 280046 531846 280102
rect 531902 280046 531998 280102
rect 531378 279978 531998 280046
rect 531378 279922 531474 279978
rect 531530 279922 531598 279978
rect 531654 279922 531722 279978
rect 531778 279922 531846 279978
rect 531902 279922 531998 279978
rect 531378 262350 531998 279922
rect 531378 262294 531474 262350
rect 531530 262294 531598 262350
rect 531654 262294 531722 262350
rect 531778 262294 531846 262350
rect 531902 262294 531998 262350
rect 531378 262226 531998 262294
rect 531378 262170 531474 262226
rect 531530 262170 531598 262226
rect 531654 262170 531722 262226
rect 531778 262170 531846 262226
rect 531902 262170 531998 262226
rect 531378 262102 531998 262170
rect 531378 262046 531474 262102
rect 531530 262046 531598 262102
rect 531654 262046 531722 262102
rect 531778 262046 531846 262102
rect 531902 262046 531998 262102
rect 531378 261978 531998 262046
rect 531378 261922 531474 261978
rect 531530 261922 531598 261978
rect 531654 261922 531722 261978
rect 531778 261922 531846 261978
rect 531902 261922 531998 261978
rect 531378 244350 531998 261922
rect 531378 244294 531474 244350
rect 531530 244294 531598 244350
rect 531654 244294 531722 244350
rect 531778 244294 531846 244350
rect 531902 244294 531998 244350
rect 531378 244226 531998 244294
rect 531378 244170 531474 244226
rect 531530 244170 531598 244226
rect 531654 244170 531722 244226
rect 531778 244170 531846 244226
rect 531902 244170 531998 244226
rect 531378 244102 531998 244170
rect 531378 244046 531474 244102
rect 531530 244046 531598 244102
rect 531654 244046 531722 244102
rect 531778 244046 531846 244102
rect 531902 244046 531998 244102
rect 531378 243978 531998 244046
rect 531378 243922 531474 243978
rect 531530 243922 531598 243978
rect 531654 243922 531722 243978
rect 531778 243922 531846 243978
rect 531902 243922 531998 243978
rect 531378 226350 531998 243922
rect 531378 226294 531474 226350
rect 531530 226294 531598 226350
rect 531654 226294 531722 226350
rect 531778 226294 531846 226350
rect 531902 226294 531998 226350
rect 531378 226226 531998 226294
rect 531378 226170 531474 226226
rect 531530 226170 531598 226226
rect 531654 226170 531722 226226
rect 531778 226170 531846 226226
rect 531902 226170 531998 226226
rect 531378 226102 531998 226170
rect 531378 226046 531474 226102
rect 531530 226046 531598 226102
rect 531654 226046 531722 226102
rect 531778 226046 531846 226102
rect 531902 226046 531998 226102
rect 531378 225978 531998 226046
rect 531378 225922 531474 225978
rect 531530 225922 531598 225978
rect 531654 225922 531722 225978
rect 531778 225922 531846 225978
rect 531902 225922 531998 225978
rect 531378 208350 531998 225922
rect 531378 208294 531474 208350
rect 531530 208294 531598 208350
rect 531654 208294 531722 208350
rect 531778 208294 531846 208350
rect 531902 208294 531998 208350
rect 531378 208226 531998 208294
rect 531378 208170 531474 208226
rect 531530 208170 531598 208226
rect 531654 208170 531722 208226
rect 531778 208170 531846 208226
rect 531902 208170 531998 208226
rect 531378 208102 531998 208170
rect 531378 208046 531474 208102
rect 531530 208046 531598 208102
rect 531654 208046 531722 208102
rect 531778 208046 531846 208102
rect 531902 208046 531998 208102
rect 531378 207978 531998 208046
rect 531378 207922 531474 207978
rect 531530 207922 531598 207978
rect 531654 207922 531722 207978
rect 531778 207922 531846 207978
rect 531902 207922 531998 207978
rect 531378 190350 531998 207922
rect 531378 190294 531474 190350
rect 531530 190294 531598 190350
rect 531654 190294 531722 190350
rect 531778 190294 531846 190350
rect 531902 190294 531998 190350
rect 531378 190226 531998 190294
rect 531378 190170 531474 190226
rect 531530 190170 531598 190226
rect 531654 190170 531722 190226
rect 531778 190170 531846 190226
rect 531902 190170 531998 190226
rect 531378 190102 531998 190170
rect 531378 190046 531474 190102
rect 531530 190046 531598 190102
rect 531654 190046 531722 190102
rect 531778 190046 531846 190102
rect 531902 190046 531998 190102
rect 531378 189978 531998 190046
rect 531378 189922 531474 189978
rect 531530 189922 531598 189978
rect 531654 189922 531722 189978
rect 531778 189922 531846 189978
rect 531902 189922 531998 189978
rect 531378 172350 531998 189922
rect 531378 172294 531474 172350
rect 531530 172294 531598 172350
rect 531654 172294 531722 172350
rect 531778 172294 531846 172350
rect 531902 172294 531998 172350
rect 531378 172226 531998 172294
rect 531378 172170 531474 172226
rect 531530 172170 531598 172226
rect 531654 172170 531722 172226
rect 531778 172170 531846 172226
rect 531902 172170 531998 172226
rect 531378 172102 531998 172170
rect 531378 172046 531474 172102
rect 531530 172046 531598 172102
rect 531654 172046 531722 172102
rect 531778 172046 531846 172102
rect 531902 172046 531998 172102
rect 531378 171978 531998 172046
rect 531378 171922 531474 171978
rect 531530 171922 531598 171978
rect 531654 171922 531722 171978
rect 531778 171922 531846 171978
rect 531902 171922 531998 171978
rect 531378 154350 531998 171922
rect 531378 154294 531474 154350
rect 531530 154294 531598 154350
rect 531654 154294 531722 154350
rect 531778 154294 531846 154350
rect 531902 154294 531998 154350
rect 531378 154226 531998 154294
rect 531378 154170 531474 154226
rect 531530 154170 531598 154226
rect 531654 154170 531722 154226
rect 531778 154170 531846 154226
rect 531902 154170 531998 154226
rect 531378 154102 531998 154170
rect 531378 154046 531474 154102
rect 531530 154046 531598 154102
rect 531654 154046 531722 154102
rect 531778 154046 531846 154102
rect 531902 154046 531998 154102
rect 531378 153978 531998 154046
rect 531378 153922 531474 153978
rect 531530 153922 531598 153978
rect 531654 153922 531722 153978
rect 531778 153922 531846 153978
rect 531902 153922 531998 153978
rect 531378 136350 531998 153922
rect 531378 136294 531474 136350
rect 531530 136294 531598 136350
rect 531654 136294 531722 136350
rect 531778 136294 531846 136350
rect 531902 136294 531998 136350
rect 531378 136226 531998 136294
rect 531378 136170 531474 136226
rect 531530 136170 531598 136226
rect 531654 136170 531722 136226
rect 531778 136170 531846 136226
rect 531902 136170 531998 136226
rect 531378 136102 531998 136170
rect 531378 136046 531474 136102
rect 531530 136046 531598 136102
rect 531654 136046 531722 136102
rect 531778 136046 531846 136102
rect 531902 136046 531998 136102
rect 531378 135978 531998 136046
rect 531378 135922 531474 135978
rect 531530 135922 531598 135978
rect 531654 135922 531722 135978
rect 531778 135922 531846 135978
rect 531902 135922 531998 135978
rect 531378 118350 531998 135922
rect 531378 118294 531474 118350
rect 531530 118294 531598 118350
rect 531654 118294 531722 118350
rect 531778 118294 531846 118350
rect 531902 118294 531998 118350
rect 531378 118226 531998 118294
rect 531378 118170 531474 118226
rect 531530 118170 531598 118226
rect 531654 118170 531722 118226
rect 531778 118170 531846 118226
rect 531902 118170 531998 118226
rect 531378 118102 531998 118170
rect 531378 118046 531474 118102
rect 531530 118046 531598 118102
rect 531654 118046 531722 118102
rect 531778 118046 531846 118102
rect 531902 118046 531998 118102
rect 531378 117978 531998 118046
rect 531378 117922 531474 117978
rect 531530 117922 531598 117978
rect 531654 117922 531722 117978
rect 531778 117922 531846 117978
rect 531902 117922 531998 117978
rect 531378 100350 531998 117922
rect 531378 100294 531474 100350
rect 531530 100294 531598 100350
rect 531654 100294 531722 100350
rect 531778 100294 531846 100350
rect 531902 100294 531998 100350
rect 531378 100226 531998 100294
rect 531378 100170 531474 100226
rect 531530 100170 531598 100226
rect 531654 100170 531722 100226
rect 531778 100170 531846 100226
rect 531902 100170 531998 100226
rect 531378 100102 531998 100170
rect 531378 100046 531474 100102
rect 531530 100046 531598 100102
rect 531654 100046 531722 100102
rect 531778 100046 531846 100102
rect 531902 100046 531998 100102
rect 531378 99978 531998 100046
rect 531378 99922 531474 99978
rect 531530 99922 531598 99978
rect 531654 99922 531722 99978
rect 531778 99922 531846 99978
rect 531902 99922 531998 99978
rect 531378 82350 531998 99922
rect 531378 82294 531474 82350
rect 531530 82294 531598 82350
rect 531654 82294 531722 82350
rect 531778 82294 531846 82350
rect 531902 82294 531998 82350
rect 531378 82226 531998 82294
rect 531378 82170 531474 82226
rect 531530 82170 531598 82226
rect 531654 82170 531722 82226
rect 531778 82170 531846 82226
rect 531902 82170 531998 82226
rect 531378 82102 531998 82170
rect 531378 82046 531474 82102
rect 531530 82046 531598 82102
rect 531654 82046 531722 82102
rect 531778 82046 531846 82102
rect 531902 82046 531998 82102
rect 531378 81978 531998 82046
rect 531378 81922 531474 81978
rect 531530 81922 531598 81978
rect 531654 81922 531722 81978
rect 531778 81922 531846 81978
rect 531902 81922 531998 81978
rect 531378 64350 531998 81922
rect 531378 64294 531474 64350
rect 531530 64294 531598 64350
rect 531654 64294 531722 64350
rect 531778 64294 531846 64350
rect 531902 64294 531998 64350
rect 531378 64226 531998 64294
rect 531378 64170 531474 64226
rect 531530 64170 531598 64226
rect 531654 64170 531722 64226
rect 531778 64170 531846 64226
rect 531902 64170 531998 64226
rect 531378 64102 531998 64170
rect 531378 64046 531474 64102
rect 531530 64046 531598 64102
rect 531654 64046 531722 64102
rect 531778 64046 531846 64102
rect 531902 64046 531998 64102
rect 531378 63978 531998 64046
rect 531378 63922 531474 63978
rect 531530 63922 531598 63978
rect 531654 63922 531722 63978
rect 531778 63922 531846 63978
rect 531902 63922 531998 63978
rect 531378 46350 531998 63922
rect 558378 597212 558998 598268
rect 558378 597156 558474 597212
rect 558530 597156 558598 597212
rect 558654 597156 558722 597212
rect 558778 597156 558846 597212
rect 558902 597156 558998 597212
rect 558378 597088 558998 597156
rect 558378 597032 558474 597088
rect 558530 597032 558598 597088
rect 558654 597032 558722 597088
rect 558778 597032 558846 597088
rect 558902 597032 558998 597088
rect 558378 596964 558998 597032
rect 558378 596908 558474 596964
rect 558530 596908 558598 596964
rect 558654 596908 558722 596964
rect 558778 596908 558846 596964
rect 558902 596908 558998 596964
rect 558378 596840 558998 596908
rect 558378 596784 558474 596840
rect 558530 596784 558598 596840
rect 558654 596784 558722 596840
rect 558778 596784 558846 596840
rect 558902 596784 558998 596840
rect 558378 580350 558998 596784
rect 558378 580294 558474 580350
rect 558530 580294 558598 580350
rect 558654 580294 558722 580350
rect 558778 580294 558846 580350
rect 558902 580294 558998 580350
rect 558378 580226 558998 580294
rect 558378 580170 558474 580226
rect 558530 580170 558598 580226
rect 558654 580170 558722 580226
rect 558778 580170 558846 580226
rect 558902 580170 558998 580226
rect 558378 580102 558998 580170
rect 558378 580046 558474 580102
rect 558530 580046 558598 580102
rect 558654 580046 558722 580102
rect 558778 580046 558846 580102
rect 558902 580046 558998 580102
rect 558378 579978 558998 580046
rect 558378 579922 558474 579978
rect 558530 579922 558598 579978
rect 558654 579922 558722 579978
rect 558778 579922 558846 579978
rect 558902 579922 558998 579978
rect 558378 562350 558998 579922
rect 558378 562294 558474 562350
rect 558530 562294 558598 562350
rect 558654 562294 558722 562350
rect 558778 562294 558846 562350
rect 558902 562294 558998 562350
rect 558378 562226 558998 562294
rect 558378 562170 558474 562226
rect 558530 562170 558598 562226
rect 558654 562170 558722 562226
rect 558778 562170 558846 562226
rect 558902 562170 558998 562226
rect 558378 562102 558998 562170
rect 558378 562046 558474 562102
rect 558530 562046 558598 562102
rect 558654 562046 558722 562102
rect 558778 562046 558846 562102
rect 558902 562046 558998 562102
rect 558378 561978 558998 562046
rect 558378 561922 558474 561978
rect 558530 561922 558598 561978
rect 558654 561922 558722 561978
rect 558778 561922 558846 561978
rect 558902 561922 558998 561978
rect 558378 544350 558998 561922
rect 558378 544294 558474 544350
rect 558530 544294 558598 544350
rect 558654 544294 558722 544350
rect 558778 544294 558846 544350
rect 558902 544294 558998 544350
rect 558378 544226 558998 544294
rect 558378 544170 558474 544226
rect 558530 544170 558598 544226
rect 558654 544170 558722 544226
rect 558778 544170 558846 544226
rect 558902 544170 558998 544226
rect 558378 544102 558998 544170
rect 558378 544046 558474 544102
rect 558530 544046 558598 544102
rect 558654 544046 558722 544102
rect 558778 544046 558846 544102
rect 558902 544046 558998 544102
rect 558378 543978 558998 544046
rect 558378 543922 558474 543978
rect 558530 543922 558598 543978
rect 558654 543922 558722 543978
rect 558778 543922 558846 543978
rect 558902 543922 558998 543978
rect 558378 526350 558998 543922
rect 558378 526294 558474 526350
rect 558530 526294 558598 526350
rect 558654 526294 558722 526350
rect 558778 526294 558846 526350
rect 558902 526294 558998 526350
rect 558378 526226 558998 526294
rect 558378 526170 558474 526226
rect 558530 526170 558598 526226
rect 558654 526170 558722 526226
rect 558778 526170 558846 526226
rect 558902 526170 558998 526226
rect 558378 526102 558998 526170
rect 558378 526046 558474 526102
rect 558530 526046 558598 526102
rect 558654 526046 558722 526102
rect 558778 526046 558846 526102
rect 558902 526046 558998 526102
rect 558378 525978 558998 526046
rect 558378 525922 558474 525978
rect 558530 525922 558598 525978
rect 558654 525922 558722 525978
rect 558778 525922 558846 525978
rect 558902 525922 558998 525978
rect 558378 508350 558998 525922
rect 558378 508294 558474 508350
rect 558530 508294 558598 508350
rect 558654 508294 558722 508350
rect 558778 508294 558846 508350
rect 558902 508294 558998 508350
rect 558378 508226 558998 508294
rect 558378 508170 558474 508226
rect 558530 508170 558598 508226
rect 558654 508170 558722 508226
rect 558778 508170 558846 508226
rect 558902 508170 558998 508226
rect 558378 508102 558998 508170
rect 558378 508046 558474 508102
rect 558530 508046 558598 508102
rect 558654 508046 558722 508102
rect 558778 508046 558846 508102
rect 558902 508046 558998 508102
rect 558378 507978 558998 508046
rect 558378 507922 558474 507978
rect 558530 507922 558598 507978
rect 558654 507922 558722 507978
rect 558778 507922 558846 507978
rect 558902 507922 558998 507978
rect 558378 490350 558998 507922
rect 558378 490294 558474 490350
rect 558530 490294 558598 490350
rect 558654 490294 558722 490350
rect 558778 490294 558846 490350
rect 558902 490294 558998 490350
rect 558378 490226 558998 490294
rect 558378 490170 558474 490226
rect 558530 490170 558598 490226
rect 558654 490170 558722 490226
rect 558778 490170 558846 490226
rect 558902 490170 558998 490226
rect 558378 490102 558998 490170
rect 558378 490046 558474 490102
rect 558530 490046 558598 490102
rect 558654 490046 558722 490102
rect 558778 490046 558846 490102
rect 558902 490046 558998 490102
rect 558378 489978 558998 490046
rect 558378 489922 558474 489978
rect 558530 489922 558598 489978
rect 558654 489922 558722 489978
rect 558778 489922 558846 489978
rect 558902 489922 558998 489978
rect 558378 472350 558998 489922
rect 558378 472294 558474 472350
rect 558530 472294 558598 472350
rect 558654 472294 558722 472350
rect 558778 472294 558846 472350
rect 558902 472294 558998 472350
rect 558378 472226 558998 472294
rect 558378 472170 558474 472226
rect 558530 472170 558598 472226
rect 558654 472170 558722 472226
rect 558778 472170 558846 472226
rect 558902 472170 558998 472226
rect 558378 472102 558998 472170
rect 558378 472046 558474 472102
rect 558530 472046 558598 472102
rect 558654 472046 558722 472102
rect 558778 472046 558846 472102
rect 558902 472046 558998 472102
rect 558378 471978 558998 472046
rect 558378 471922 558474 471978
rect 558530 471922 558598 471978
rect 558654 471922 558722 471978
rect 558778 471922 558846 471978
rect 558902 471922 558998 471978
rect 558378 454350 558998 471922
rect 558378 454294 558474 454350
rect 558530 454294 558598 454350
rect 558654 454294 558722 454350
rect 558778 454294 558846 454350
rect 558902 454294 558998 454350
rect 558378 454226 558998 454294
rect 558378 454170 558474 454226
rect 558530 454170 558598 454226
rect 558654 454170 558722 454226
rect 558778 454170 558846 454226
rect 558902 454170 558998 454226
rect 558378 454102 558998 454170
rect 558378 454046 558474 454102
rect 558530 454046 558598 454102
rect 558654 454046 558722 454102
rect 558778 454046 558846 454102
rect 558902 454046 558998 454102
rect 558378 453978 558998 454046
rect 558378 453922 558474 453978
rect 558530 453922 558598 453978
rect 558654 453922 558722 453978
rect 558778 453922 558846 453978
rect 558902 453922 558998 453978
rect 558378 436350 558998 453922
rect 558378 436294 558474 436350
rect 558530 436294 558598 436350
rect 558654 436294 558722 436350
rect 558778 436294 558846 436350
rect 558902 436294 558998 436350
rect 558378 436226 558998 436294
rect 558378 436170 558474 436226
rect 558530 436170 558598 436226
rect 558654 436170 558722 436226
rect 558778 436170 558846 436226
rect 558902 436170 558998 436226
rect 558378 436102 558998 436170
rect 558378 436046 558474 436102
rect 558530 436046 558598 436102
rect 558654 436046 558722 436102
rect 558778 436046 558846 436102
rect 558902 436046 558998 436102
rect 558378 435978 558998 436046
rect 558378 435922 558474 435978
rect 558530 435922 558598 435978
rect 558654 435922 558722 435978
rect 558778 435922 558846 435978
rect 558902 435922 558998 435978
rect 558378 418350 558998 435922
rect 558378 418294 558474 418350
rect 558530 418294 558598 418350
rect 558654 418294 558722 418350
rect 558778 418294 558846 418350
rect 558902 418294 558998 418350
rect 558378 418226 558998 418294
rect 558378 418170 558474 418226
rect 558530 418170 558598 418226
rect 558654 418170 558722 418226
rect 558778 418170 558846 418226
rect 558902 418170 558998 418226
rect 558378 418102 558998 418170
rect 558378 418046 558474 418102
rect 558530 418046 558598 418102
rect 558654 418046 558722 418102
rect 558778 418046 558846 418102
rect 558902 418046 558998 418102
rect 558378 417978 558998 418046
rect 558378 417922 558474 417978
rect 558530 417922 558598 417978
rect 558654 417922 558722 417978
rect 558778 417922 558846 417978
rect 558902 417922 558998 417978
rect 558378 400350 558998 417922
rect 558378 400294 558474 400350
rect 558530 400294 558598 400350
rect 558654 400294 558722 400350
rect 558778 400294 558846 400350
rect 558902 400294 558998 400350
rect 558378 400226 558998 400294
rect 558378 400170 558474 400226
rect 558530 400170 558598 400226
rect 558654 400170 558722 400226
rect 558778 400170 558846 400226
rect 558902 400170 558998 400226
rect 558378 400102 558998 400170
rect 558378 400046 558474 400102
rect 558530 400046 558598 400102
rect 558654 400046 558722 400102
rect 558778 400046 558846 400102
rect 558902 400046 558998 400102
rect 558378 399978 558998 400046
rect 558378 399922 558474 399978
rect 558530 399922 558598 399978
rect 558654 399922 558722 399978
rect 558778 399922 558846 399978
rect 558902 399922 558998 399978
rect 558378 382350 558998 399922
rect 558378 382294 558474 382350
rect 558530 382294 558598 382350
rect 558654 382294 558722 382350
rect 558778 382294 558846 382350
rect 558902 382294 558998 382350
rect 558378 382226 558998 382294
rect 558378 382170 558474 382226
rect 558530 382170 558598 382226
rect 558654 382170 558722 382226
rect 558778 382170 558846 382226
rect 558902 382170 558998 382226
rect 558378 382102 558998 382170
rect 558378 382046 558474 382102
rect 558530 382046 558598 382102
rect 558654 382046 558722 382102
rect 558778 382046 558846 382102
rect 558902 382046 558998 382102
rect 558378 381978 558998 382046
rect 558378 381922 558474 381978
rect 558530 381922 558598 381978
rect 558654 381922 558722 381978
rect 558778 381922 558846 381978
rect 558902 381922 558998 381978
rect 558378 364350 558998 381922
rect 558378 364294 558474 364350
rect 558530 364294 558598 364350
rect 558654 364294 558722 364350
rect 558778 364294 558846 364350
rect 558902 364294 558998 364350
rect 558378 364226 558998 364294
rect 558378 364170 558474 364226
rect 558530 364170 558598 364226
rect 558654 364170 558722 364226
rect 558778 364170 558846 364226
rect 558902 364170 558998 364226
rect 558378 364102 558998 364170
rect 558378 364046 558474 364102
rect 558530 364046 558598 364102
rect 558654 364046 558722 364102
rect 558778 364046 558846 364102
rect 558902 364046 558998 364102
rect 558378 363978 558998 364046
rect 558378 363922 558474 363978
rect 558530 363922 558598 363978
rect 558654 363922 558722 363978
rect 558778 363922 558846 363978
rect 558902 363922 558998 363978
rect 558378 346350 558998 363922
rect 558378 346294 558474 346350
rect 558530 346294 558598 346350
rect 558654 346294 558722 346350
rect 558778 346294 558846 346350
rect 558902 346294 558998 346350
rect 558378 346226 558998 346294
rect 558378 346170 558474 346226
rect 558530 346170 558598 346226
rect 558654 346170 558722 346226
rect 558778 346170 558846 346226
rect 558902 346170 558998 346226
rect 558378 346102 558998 346170
rect 558378 346046 558474 346102
rect 558530 346046 558598 346102
rect 558654 346046 558722 346102
rect 558778 346046 558846 346102
rect 558902 346046 558998 346102
rect 558378 345978 558998 346046
rect 558378 345922 558474 345978
rect 558530 345922 558598 345978
rect 558654 345922 558722 345978
rect 558778 345922 558846 345978
rect 558902 345922 558998 345978
rect 558378 328350 558998 345922
rect 558378 328294 558474 328350
rect 558530 328294 558598 328350
rect 558654 328294 558722 328350
rect 558778 328294 558846 328350
rect 558902 328294 558998 328350
rect 558378 328226 558998 328294
rect 558378 328170 558474 328226
rect 558530 328170 558598 328226
rect 558654 328170 558722 328226
rect 558778 328170 558846 328226
rect 558902 328170 558998 328226
rect 558378 328102 558998 328170
rect 558378 328046 558474 328102
rect 558530 328046 558598 328102
rect 558654 328046 558722 328102
rect 558778 328046 558846 328102
rect 558902 328046 558998 328102
rect 558378 327978 558998 328046
rect 558378 327922 558474 327978
rect 558530 327922 558598 327978
rect 558654 327922 558722 327978
rect 558778 327922 558846 327978
rect 558902 327922 558998 327978
rect 558378 310350 558998 327922
rect 558378 310294 558474 310350
rect 558530 310294 558598 310350
rect 558654 310294 558722 310350
rect 558778 310294 558846 310350
rect 558902 310294 558998 310350
rect 558378 310226 558998 310294
rect 558378 310170 558474 310226
rect 558530 310170 558598 310226
rect 558654 310170 558722 310226
rect 558778 310170 558846 310226
rect 558902 310170 558998 310226
rect 558378 310102 558998 310170
rect 558378 310046 558474 310102
rect 558530 310046 558598 310102
rect 558654 310046 558722 310102
rect 558778 310046 558846 310102
rect 558902 310046 558998 310102
rect 558378 309978 558998 310046
rect 558378 309922 558474 309978
rect 558530 309922 558598 309978
rect 558654 309922 558722 309978
rect 558778 309922 558846 309978
rect 558902 309922 558998 309978
rect 558378 292350 558998 309922
rect 558378 292294 558474 292350
rect 558530 292294 558598 292350
rect 558654 292294 558722 292350
rect 558778 292294 558846 292350
rect 558902 292294 558998 292350
rect 558378 292226 558998 292294
rect 558378 292170 558474 292226
rect 558530 292170 558598 292226
rect 558654 292170 558722 292226
rect 558778 292170 558846 292226
rect 558902 292170 558998 292226
rect 558378 292102 558998 292170
rect 558378 292046 558474 292102
rect 558530 292046 558598 292102
rect 558654 292046 558722 292102
rect 558778 292046 558846 292102
rect 558902 292046 558998 292102
rect 558378 291978 558998 292046
rect 558378 291922 558474 291978
rect 558530 291922 558598 291978
rect 558654 291922 558722 291978
rect 558778 291922 558846 291978
rect 558902 291922 558998 291978
rect 558378 274350 558998 291922
rect 558378 274294 558474 274350
rect 558530 274294 558598 274350
rect 558654 274294 558722 274350
rect 558778 274294 558846 274350
rect 558902 274294 558998 274350
rect 558378 274226 558998 274294
rect 558378 274170 558474 274226
rect 558530 274170 558598 274226
rect 558654 274170 558722 274226
rect 558778 274170 558846 274226
rect 558902 274170 558998 274226
rect 558378 274102 558998 274170
rect 558378 274046 558474 274102
rect 558530 274046 558598 274102
rect 558654 274046 558722 274102
rect 558778 274046 558846 274102
rect 558902 274046 558998 274102
rect 558378 273978 558998 274046
rect 558378 273922 558474 273978
rect 558530 273922 558598 273978
rect 558654 273922 558722 273978
rect 558778 273922 558846 273978
rect 558902 273922 558998 273978
rect 558378 256350 558998 273922
rect 558378 256294 558474 256350
rect 558530 256294 558598 256350
rect 558654 256294 558722 256350
rect 558778 256294 558846 256350
rect 558902 256294 558998 256350
rect 558378 256226 558998 256294
rect 558378 256170 558474 256226
rect 558530 256170 558598 256226
rect 558654 256170 558722 256226
rect 558778 256170 558846 256226
rect 558902 256170 558998 256226
rect 558378 256102 558998 256170
rect 558378 256046 558474 256102
rect 558530 256046 558598 256102
rect 558654 256046 558722 256102
rect 558778 256046 558846 256102
rect 558902 256046 558998 256102
rect 558378 255978 558998 256046
rect 558378 255922 558474 255978
rect 558530 255922 558598 255978
rect 558654 255922 558722 255978
rect 558778 255922 558846 255978
rect 558902 255922 558998 255978
rect 558378 238350 558998 255922
rect 558378 238294 558474 238350
rect 558530 238294 558598 238350
rect 558654 238294 558722 238350
rect 558778 238294 558846 238350
rect 558902 238294 558998 238350
rect 558378 238226 558998 238294
rect 558378 238170 558474 238226
rect 558530 238170 558598 238226
rect 558654 238170 558722 238226
rect 558778 238170 558846 238226
rect 558902 238170 558998 238226
rect 558378 238102 558998 238170
rect 558378 238046 558474 238102
rect 558530 238046 558598 238102
rect 558654 238046 558722 238102
rect 558778 238046 558846 238102
rect 558902 238046 558998 238102
rect 558378 237978 558998 238046
rect 558378 237922 558474 237978
rect 558530 237922 558598 237978
rect 558654 237922 558722 237978
rect 558778 237922 558846 237978
rect 558902 237922 558998 237978
rect 558378 220350 558998 237922
rect 558378 220294 558474 220350
rect 558530 220294 558598 220350
rect 558654 220294 558722 220350
rect 558778 220294 558846 220350
rect 558902 220294 558998 220350
rect 558378 220226 558998 220294
rect 558378 220170 558474 220226
rect 558530 220170 558598 220226
rect 558654 220170 558722 220226
rect 558778 220170 558846 220226
rect 558902 220170 558998 220226
rect 558378 220102 558998 220170
rect 558378 220046 558474 220102
rect 558530 220046 558598 220102
rect 558654 220046 558722 220102
rect 558778 220046 558846 220102
rect 558902 220046 558998 220102
rect 558378 219978 558998 220046
rect 558378 219922 558474 219978
rect 558530 219922 558598 219978
rect 558654 219922 558722 219978
rect 558778 219922 558846 219978
rect 558902 219922 558998 219978
rect 558378 202350 558998 219922
rect 558378 202294 558474 202350
rect 558530 202294 558598 202350
rect 558654 202294 558722 202350
rect 558778 202294 558846 202350
rect 558902 202294 558998 202350
rect 558378 202226 558998 202294
rect 558378 202170 558474 202226
rect 558530 202170 558598 202226
rect 558654 202170 558722 202226
rect 558778 202170 558846 202226
rect 558902 202170 558998 202226
rect 558378 202102 558998 202170
rect 558378 202046 558474 202102
rect 558530 202046 558598 202102
rect 558654 202046 558722 202102
rect 558778 202046 558846 202102
rect 558902 202046 558998 202102
rect 558378 201978 558998 202046
rect 558378 201922 558474 201978
rect 558530 201922 558598 201978
rect 558654 201922 558722 201978
rect 558778 201922 558846 201978
rect 558902 201922 558998 201978
rect 558378 184350 558998 201922
rect 558378 184294 558474 184350
rect 558530 184294 558598 184350
rect 558654 184294 558722 184350
rect 558778 184294 558846 184350
rect 558902 184294 558998 184350
rect 558378 184226 558998 184294
rect 558378 184170 558474 184226
rect 558530 184170 558598 184226
rect 558654 184170 558722 184226
rect 558778 184170 558846 184226
rect 558902 184170 558998 184226
rect 558378 184102 558998 184170
rect 558378 184046 558474 184102
rect 558530 184046 558598 184102
rect 558654 184046 558722 184102
rect 558778 184046 558846 184102
rect 558902 184046 558998 184102
rect 558378 183978 558998 184046
rect 558378 183922 558474 183978
rect 558530 183922 558598 183978
rect 558654 183922 558722 183978
rect 558778 183922 558846 183978
rect 558902 183922 558998 183978
rect 558378 166350 558998 183922
rect 558378 166294 558474 166350
rect 558530 166294 558598 166350
rect 558654 166294 558722 166350
rect 558778 166294 558846 166350
rect 558902 166294 558998 166350
rect 558378 166226 558998 166294
rect 558378 166170 558474 166226
rect 558530 166170 558598 166226
rect 558654 166170 558722 166226
rect 558778 166170 558846 166226
rect 558902 166170 558998 166226
rect 558378 166102 558998 166170
rect 558378 166046 558474 166102
rect 558530 166046 558598 166102
rect 558654 166046 558722 166102
rect 558778 166046 558846 166102
rect 558902 166046 558998 166102
rect 558378 165978 558998 166046
rect 558378 165922 558474 165978
rect 558530 165922 558598 165978
rect 558654 165922 558722 165978
rect 558778 165922 558846 165978
rect 558902 165922 558998 165978
rect 558378 148350 558998 165922
rect 558378 148294 558474 148350
rect 558530 148294 558598 148350
rect 558654 148294 558722 148350
rect 558778 148294 558846 148350
rect 558902 148294 558998 148350
rect 558378 148226 558998 148294
rect 558378 148170 558474 148226
rect 558530 148170 558598 148226
rect 558654 148170 558722 148226
rect 558778 148170 558846 148226
rect 558902 148170 558998 148226
rect 558378 148102 558998 148170
rect 558378 148046 558474 148102
rect 558530 148046 558598 148102
rect 558654 148046 558722 148102
rect 558778 148046 558846 148102
rect 558902 148046 558998 148102
rect 558378 147978 558998 148046
rect 558378 147922 558474 147978
rect 558530 147922 558598 147978
rect 558654 147922 558722 147978
rect 558778 147922 558846 147978
rect 558902 147922 558998 147978
rect 558378 130350 558998 147922
rect 558378 130294 558474 130350
rect 558530 130294 558598 130350
rect 558654 130294 558722 130350
rect 558778 130294 558846 130350
rect 558902 130294 558998 130350
rect 558378 130226 558998 130294
rect 558378 130170 558474 130226
rect 558530 130170 558598 130226
rect 558654 130170 558722 130226
rect 558778 130170 558846 130226
rect 558902 130170 558998 130226
rect 558378 130102 558998 130170
rect 558378 130046 558474 130102
rect 558530 130046 558598 130102
rect 558654 130046 558722 130102
rect 558778 130046 558846 130102
rect 558902 130046 558998 130102
rect 558378 129978 558998 130046
rect 558378 129922 558474 129978
rect 558530 129922 558598 129978
rect 558654 129922 558722 129978
rect 558778 129922 558846 129978
rect 558902 129922 558998 129978
rect 558378 112350 558998 129922
rect 558378 112294 558474 112350
rect 558530 112294 558598 112350
rect 558654 112294 558722 112350
rect 558778 112294 558846 112350
rect 558902 112294 558998 112350
rect 558378 112226 558998 112294
rect 558378 112170 558474 112226
rect 558530 112170 558598 112226
rect 558654 112170 558722 112226
rect 558778 112170 558846 112226
rect 558902 112170 558998 112226
rect 558378 112102 558998 112170
rect 558378 112046 558474 112102
rect 558530 112046 558598 112102
rect 558654 112046 558722 112102
rect 558778 112046 558846 112102
rect 558902 112046 558998 112102
rect 558378 111978 558998 112046
rect 558378 111922 558474 111978
rect 558530 111922 558598 111978
rect 558654 111922 558722 111978
rect 558778 111922 558846 111978
rect 558902 111922 558998 111978
rect 558378 94350 558998 111922
rect 558378 94294 558474 94350
rect 558530 94294 558598 94350
rect 558654 94294 558722 94350
rect 558778 94294 558846 94350
rect 558902 94294 558998 94350
rect 558378 94226 558998 94294
rect 558378 94170 558474 94226
rect 558530 94170 558598 94226
rect 558654 94170 558722 94226
rect 558778 94170 558846 94226
rect 558902 94170 558998 94226
rect 558378 94102 558998 94170
rect 558378 94046 558474 94102
rect 558530 94046 558598 94102
rect 558654 94046 558722 94102
rect 558778 94046 558846 94102
rect 558902 94046 558998 94102
rect 558378 93978 558998 94046
rect 558378 93922 558474 93978
rect 558530 93922 558598 93978
rect 558654 93922 558722 93978
rect 558778 93922 558846 93978
rect 558902 93922 558998 93978
rect 558378 76350 558998 93922
rect 558378 76294 558474 76350
rect 558530 76294 558598 76350
rect 558654 76294 558722 76350
rect 558778 76294 558846 76350
rect 558902 76294 558998 76350
rect 558378 76226 558998 76294
rect 558378 76170 558474 76226
rect 558530 76170 558598 76226
rect 558654 76170 558722 76226
rect 558778 76170 558846 76226
rect 558902 76170 558998 76226
rect 558378 76102 558998 76170
rect 558378 76046 558474 76102
rect 558530 76046 558598 76102
rect 558654 76046 558722 76102
rect 558778 76046 558846 76102
rect 558902 76046 558998 76102
rect 558378 75978 558998 76046
rect 558378 75922 558474 75978
rect 558530 75922 558598 75978
rect 558654 75922 558722 75978
rect 558778 75922 558846 75978
rect 558902 75922 558998 75978
rect 558378 58350 558998 75922
rect 558378 58294 558474 58350
rect 558530 58294 558598 58350
rect 558654 58294 558722 58350
rect 558778 58294 558846 58350
rect 558902 58294 558998 58350
rect 558378 58226 558998 58294
rect 558378 58170 558474 58226
rect 558530 58170 558598 58226
rect 558654 58170 558722 58226
rect 558778 58170 558846 58226
rect 558902 58170 558998 58226
rect 558378 58102 558998 58170
rect 558378 58046 558474 58102
rect 558530 58046 558598 58102
rect 558654 58046 558722 58102
rect 558778 58046 558846 58102
rect 558902 58046 558998 58102
rect 558378 57978 558998 58046
rect 558378 57922 558474 57978
rect 558530 57922 558598 57978
rect 558654 57922 558722 57978
rect 558778 57922 558846 57978
rect 558902 57922 558998 57978
rect 539308 57178 539364 57188
rect 534268 50698 534324 50708
rect 531378 46294 531474 46350
rect 531530 46294 531598 46350
rect 531654 46294 531722 46350
rect 531778 46294 531846 46350
rect 531902 46294 531998 46350
rect 531378 46226 531998 46294
rect 531378 46170 531474 46226
rect 531530 46170 531598 46226
rect 531654 46170 531722 46226
rect 531778 46170 531846 46226
rect 531902 46170 531998 46226
rect 531378 46102 531998 46170
rect 531378 46046 531474 46102
rect 531530 46046 531598 46102
rect 531654 46046 531722 46102
rect 531778 46046 531846 46102
rect 531902 46046 531998 46102
rect 531378 45978 531998 46046
rect 531378 45922 531474 45978
rect 531530 45922 531598 45978
rect 531654 45922 531722 45978
rect 531778 45922 531846 45978
rect 531902 45922 531998 45978
rect 531378 28350 531998 45922
rect 531378 28294 531474 28350
rect 531530 28294 531598 28350
rect 531654 28294 531722 28350
rect 531778 28294 531846 28350
rect 531902 28294 531998 28350
rect 531378 28226 531998 28294
rect 531378 28170 531474 28226
rect 531530 28170 531598 28226
rect 531654 28170 531722 28226
rect 531778 28170 531846 28226
rect 531902 28170 531998 28226
rect 531378 28102 531998 28170
rect 531378 28046 531474 28102
rect 531530 28046 531598 28102
rect 531654 28046 531722 28102
rect 531778 28046 531846 28102
rect 531902 28046 531998 28102
rect 531378 27978 531998 28046
rect 531378 27922 531474 27978
rect 531530 27922 531598 27978
rect 531654 27922 531722 27978
rect 531778 27922 531846 27978
rect 531902 27922 531998 27978
rect 527658 4294 527754 4350
rect 527810 4294 527878 4350
rect 527934 4294 528002 4350
rect 528058 4294 528126 4350
rect 528182 4294 528278 4350
rect 527658 4226 528278 4294
rect 527658 4170 527754 4226
rect 527810 4170 527878 4226
rect 527934 4170 528002 4226
rect 528058 4170 528126 4226
rect 528182 4170 528278 4226
rect 500658 -1176 500754 -1120
rect 500810 -1176 500878 -1120
rect 500934 -1176 501002 -1120
rect 501058 -1176 501126 -1120
rect 501182 -1176 501278 -1120
rect 500658 -1244 501278 -1176
rect 500658 -1300 500754 -1244
rect 500810 -1300 500878 -1244
rect 500934 -1300 501002 -1244
rect 501058 -1300 501126 -1244
rect 501182 -1300 501278 -1244
rect 500658 -1368 501278 -1300
rect 500658 -1424 500754 -1368
rect 500810 -1424 500878 -1368
rect 500934 -1424 501002 -1368
rect 501058 -1424 501126 -1368
rect 501182 -1424 501278 -1368
rect 500658 -1492 501278 -1424
rect 500658 -1548 500754 -1492
rect 500810 -1548 500878 -1492
rect 500934 -1548 501002 -1492
rect 501058 -1548 501126 -1492
rect 501182 -1548 501278 -1492
rect 500658 -1644 501278 -1548
rect 527658 4102 528278 4170
rect 531132 15238 531188 15248
rect 531132 4228 531188 15182
rect 531132 4162 531188 4172
rect 531378 10350 531998 27922
rect 531378 10294 531474 10350
rect 531530 10294 531598 10350
rect 531654 10294 531722 10350
rect 531778 10294 531846 10350
rect 531902 10294 531998 10350
rect 531378 10226 531998 10294
rect 531378 10170 531474 10226
rect 531530 10170 531598 10226
rect 531654 10170 531722 10226
rect 531778 10170 531846 10226
rect 531902 10170 531998 10226
rect 531378 10102 531998 10170
rect 531378 10046 531474 10102
rect 531530 10046 531598 10102
rect 531654 10046 531722 10102
rect 531778 10046 531846 10102
rect 531902 10046 531998 10102
rect 531378 9978 531998 10046
rect 531378 9922 531474 9978
rect 531530 9922 531598 9978
rect 531654 9922 531722 9978
rect 531778 9922 531846 9978
rect 531902 9922 531998 9978
rect 527658 4046 527754 4102
rect 527810 4046 527878 4102
rect 527934 4046 528002 4102
rect 528058 4046 528126 4102
rect 528182 4046 528278 4102
rect 527658 3978 528278 4046
rect 527658 3922 527754 3978
rect 527810 3922 527878 3978
rect 527934 3922 528002 3978
rect 528058 3922 528126 3978
rect 528182 3922 528278 3978
rect 527658 -160 528278 3922
rect 527658 -216 527754 -160
rect 527810 -216 527878 -160
rect 527934 -216 528002 -160
rect 528058 -216 528126 -160
rect 528182 -216 528278 -160
rect 527658 -284 528278 -216
rect 527658 -340 527754 -284
rect 527810 -340 527878 -284
rect 527934 -340 528002 -284
rect 528058 -340 528126 -284
rect 528182 -340 528278 -284
rect 527658 -408 528278 -340
rect 527658 -464 527754 -408
rect 527810 -464 527878 -408
rect 527934 -464 528002 -408
rect 528058 -464 528126 -408
rect 528182 -464 528278 -408
rect 527658 -532 528278 -464
rect 527658 -588 527754 -532
rect 527810 -588 527878 -532
rect 527934 -588 528002 -532
rect 528058 -588 528126 -532
rect 528182 -588 528278 -532
rect 527658 -1644 528278 -588
rect 531378 -1120 531998 9922
rect 532588 47098 532644 47108
rect 532588 4228 532644 47042
rect 532588 4162 532644 4172
rect 534268 4228 534324 50642
rect 534268 4162 534324 4172
rect 537628 50518 537684 50528
rect 537628 4228 537684 50462
rect 537628 4162 537684 4172
rect 539308 4228 539364 57122
rect 554428 52138 554484 52148
rect 549388 48898 549444 48908
rect 544348 40618 544404 40628
rect 544348 20188 544404 40562
rect 544348 20132 544516 20188
rect 539308 4162 539364 4172
rect 544460 4228 544516 20132
rect 544460 4162 544516 4172
rect 549388 4228 549444 48842
rect 549388 4162 549444 4172
rect 554428 4228 554484 52082
rect 554428 4162 554484 4172
rect 558378 40350 558998 57922
rect 562098 598172 562718 598268
rect 562098 598116 562194 598172
rect 562250 598116 562318 598172
rect 562374 598116 562442 598172
rect 562498 598116 562566 598172
rect 562622 598116 562718 598172
rect 562098 598048 562718 598116
rect 562098 597992 562194 598048
rect 562250 597992 562318 598048
rect 562374 597992 562442 598048
rect 562498 597992 562566 598048
rect 562622 597992 562718 598048
rect 562098 597924 562718 597992
rect 562098 597868 562194 597924
rect 562250 597868 562318 597924
rect 562374 597868 562442 597924
rect 562498 597868 562566 597924
rect 562622 597868 562718 597924
rect 562098 597800 562718 597868
rect 562098 597744 562194 597800
rect 562250 597744 562318 597800
rect 562374 597744 562442 597800
rect 562498 597744 562566 597800
rect 562622 597744 562718 597800
rect 562098 586350 562718 597744
rect 562098 586294 562194 586350
rect 562250 586294 562318 586350
rect 562374 586294 562442 586350
rect 562498 586294 562566 586350
rect 562622 586294 562718 586350
rect 562098 586226 562718 586294
rect 562098 586170 562194 586226
rect 562250 586170 562318 586226
rect 562374 586170 562442 586226
rect 562498 586170 562566 586226
rect 562622 586170 562718 586226
rect 562098 586102 562718 586170
rect 562098 586046 562194 586102
rect 562250 586046 562318 586102
rect 562374 586046 562442 586102
rect 562498 586046 562566 586102
rect 562622 586046 562718 586102
rect 562098 585978 562718 586046
rect 562098 585922 562194 585978
rect 562250 585922 562318 585978
rect 562374 585922 562442 585978
rect 562498 585922 562566 585978
rect 562622 585922 562718 585978
rect 562098 568350 562718 585922
rect 562098 568294 562194 568350
rect 562250 568294 562318 568350
rect 562374 568294 562442 568350
rect 562498 568294 562566 568350
rect 562622 568294 562718 568350
rect 562098 568226 562718 568294
rect 562098 568170 562194 568226
rect 562250 568170 562318 568226
rect 562374 568170 562442 568226
rect 562498 568170 562566 568226
rect 562622 568170 562718 568226
rect 562098 568102 562718 568170
rect 562098 568046 562194 568102
rect 562250 568046 562318 568102
rect 562374 568046 562442 568102
rect 562498 568046 562566 568102
rect 562622 568046 562718 568102
rect 562098 567978 562718 568046
rect 562098 567922 562194 567978
rect 562250 567922 562318 567978
rect 562374 567922 562442 567978
rect 562498 567922 562566 567978
rect 562622 567922 562718 567978
rect 562098 550350 562718 567922
rect 562098 550294 562194 550350
rect 562250 550294 562318 550350
rect 562374 550294 562442 550350
rect 562498 550294 562566 550350
rect 562622 550294 562718 550350
rect 562098 550226 562718 550294
rect 562098 550170 562194 550226
rect 562250 550170 562318 550226
rect 562374 550170 562442 550226
rect 562498 550170 562566 550226
rect 562622 550170 562718 550226
rect 562098 550102 562718 550170
rect 562098 550046 562194 550102
rect 562250 550046 562318 550102
rect 562374 550046 562442 550102
rect 562498 550046 562566 550102
rect 562622 550046 562718 550102
rect 562098 549978 562718 550046
rect 562098 549922 562194 549978
rect 562250 549922 562318 549978
rect 562374 549922 562442 549978
rect 562498 549922 562566 549978
rect 562622 549922 562718 549978
rect 562098 532350 562718 549922
rect 562098 532294 562194 532350
rect 562250 532294 562318 532350
rect 562374 532294 562442 532350
rect 562498 532294 562566 532350
rect 562622 532294 562718 532350
rect 562098 532226 562718 532294
rect 562098 532170 562194 532226
rect 562250 532170 562318 532226
rect 562374 532170 562442 532226
rect 562498 532170 562566 532226
rect 562622 532170 562718 532226
rect 562098 532102 562718 532170
rect 562098 532046 562194 532102
rect 562250 532046 562318 532102
rect 562374 532046 562442 532102
rect 562498 532046 562566 532102
rect 562622 532046 562718 532102
rect 562098 531978 562718 532046
rect 562098 531922 562194 531978
rect 562250 531922 562318 531978
rect 562374 531922 562442 531978
rect 562498 531922 562566 531978
rect 562622 531922 562718 531978
rect 562098 514350 562718 531922
rect 562098 514294 562194 514350
rect 562250 514294 562318 514350
rect 562374 514294 562442 514350
rect 562498 514294 562566 514350
rect 562622 514294 562718 514350
rect 562098 514226 562718 514294
rect 562098 514170 562194 514226
rect 562250 514170 562318 514226
rect 562374 514170 562442 514226
rect 562498 514170 562566 514226
rect 562622 514170 562718 514226
rect 562098 514102 562718 514170
rect 562098 514046 562194 514102
rect 562250 514046 562318 514102
rect 562374 514046 562442 514102
rect 562498 514046 562566 514102
rect 562622 514046 562718 514102
rect 562098 513978 562718 514046
rect 562098 513922 562194 513978
rect 562250 513922 562318 513978
rect 562374 513922 562442 513978
rect 562498 513922 562566 513978
rect 562622 513922 562718 513978
rect 562098 496350 562718 513922
rect 562098 496294 562194 496350
rect 562250 496294 562318 496350
rect 562374 496294 562442 496350
rect 562498 496294 562566 496350
rect 562622 496294 562718 496350
rect 562098 496226 562718 496294
rect 562098 496170 562194 496226
rect 562250 496170 562318 496226
rect 562374 496170 562442 496226
rect 562498 496170 562566 496226
rect 562622 496170 562718 496226
rect 562098 496102 562718 496170
rect 562098 496046 562194 496102
rect 562250 496046 562318 496102
rect 562374 496046 562442 496102
rect 562498 496046 562566 496102
rect 562622 496046 562718 496102
rect 562098 495978 562718 496046
rect 562098 495922 562194 495978
rect 562250 495922 562318 495978
rect 562374 495922 562442 495978
rect 562498 495922 562566 495978
rect 562622 495922 562718 495978
rect 562098 478350 562718 495922
rect 562098 478294 562194 478350
rect 562250 478294 562318 478350
rect 562374 478294 562442 478350
rect 562498 478294 562566 478350
rect 562622 478294 562718 478350
rect 562098 478226 562718 478294
rect 562098 478170 562194 478226
rect 562250 478170 562318 478226
rect 562374 478170 562442 478226
rect 562498 478170 562566 478226
rect 562622 478170 562718 478226
rect 562098 478102 562718 478170
rect 562098 478046 562194 478102
rect 562250 478046 562318 478102
rect 562374 478046 562442 478102
rect 562498 478046 562566 478102
rect 562622 478046 562718 478102
rect 562098 477978 562718 478046
rect 562098 477922 562194 477978
rect 562250 477922 562318 477978
rect 562374 477922 562442 477978
rect 562498 477922 562566 477978
rect 562622 477922 562718 477978
rect 562098 460350 562718 477922
rect 562098 460294 562194 460350
rect 562250 460294 562318 460350
rect 562374 460294 562442 460350
rect 562498 460294 562566 460350
rect 562622 460294 562718 460350
rect 562098 460226 562718 460294
rect 562098 460170 562194 460226
rect 562250 460170 562318 460226
rect 562374 460170 562442 460226
rect 562498 460170 562566 460226
rect 562622 460170 562718 460226
rect 562098 460102 562718 460170
rect 562098 460046 562194 460102
rect 562250 460046 562318 460102
rect 562374 460046 562442 460102
rect 562498 460046 562566 460102
rect 562622 460046 562718 460102
rect 562098 459978 562718 460046
rect 562098 459922 562194 459978
rect 562250 459922 562318 459978
rect 562374 459922 562442 459978
rect 562498 459922 562566 459978
rect 562622 459922 562718 459978
rect 562098 442350 562718 459922
rect 562098 442294 562194 442350
rect 562250 442294 562318 442350
rect 562374 442294 562442 442350
rect 562498 442294 562566 442350
rect 562622 442294 562718 442350
rect 562098 442226 562718 442294
rect 562098 442170 562194 442226
rect 562250 442170 562318 442226
rect 562374 442170 562442 442226
rect 562498 442170 562566 442226
rect 562622 442170 562718 442226
rect 562098 442102 562718 442170
rect 562098 442046 562194 442102
rect 562250 442046 562318 442102
rect 562374 442046 562442 442102
rect 562498 442046 562566 442102
rect 562622 442046 562718 442102
rect 562098 441978 562718 442046
rect 562098 441922 562194 441978
rect 562250 441922 562318 441978
rect 562374 441922 562442 441978
rect 562498 441922 562566 441978
rect 562622 441922 562718 441978
rect 562098 424350 562718 441922
rect 562098 424294 562194 424350
rect 562250 424294 562318 424350
rect 562374 424294 562442 424350
rect 562498 424294 562566 424350
rect 562622 424294 562718 424350
rect 562098 424226 562718 424294
rect 562098 424170 562194 424226
rect 562250 424170 562318 424226
rect 562374 424170 562442 424226
rect 562498 424170 562566 424226
rect 562622 424170 562718 424226
rect 562098 424102 562718 424170
rect 562098 424046 562194 424102
rect 562250 424046 562318 424102
rect 562374 424046 562442 424102
rect 562498 424046 562566 424102
rect 562622 424046 562718 424102
rect 562098 423978 562718 424046
rect 562098 423922 562194 423978
rect 562250 423922 562318 423978
rect 562374 423922 562442 423978
rect 562498 423922 562566 423978
rect 562622 423922 562718 423978
rect 562098 406350 562718 423922
rect 562098 406294 562194 406350
rect 562250 406294 562318 406350
rect 562374 406294 562442 406350
rect 562498 406294 562566 406350
rect 562622 406294 562718 406350
rect 562098 406226 562718 406294
rect 562098 406170 562194 406226
rect 562250 406170 562318 406226
rect 562374 406170 562442 406226
rect 562498 406170 562566 406226
rect 562622 406170 562718 406226
rect 562098 406102 562718 406170
rect 562098 406046 562194 406102
rect 562250 406046 562318 406102
rect 562374 406046 562442 406102
rect 562498 406046 562566 406102
rect 562622 406046 562718 406102
rect 562098 405978 562718 406046
rect 562098 405922 562194 405978
rect 562250 405922 562318 405978
rect 562374 405922 562442 405978
rect 562498 405922 562566 405978
rect 562622 405922 562718 405978
rect 562098 388350 562718 405922
rect 562098 388294 562194 388350
rect 562250 388294 562318 388350
rect 562374 388294 562442 388350
rect 562498 388294 562566 388350
rect 562622 388294 562718 388350
rect 562098 388226 562718 388294
rect 562098 388170 562194 388226
rect 562250 388170 562318 388226
rect 562374 388170 562442 388226
rect 562498 388170 562566 388226
rect 562622 388170 562718 388226
rect 562098 388102 562718 388170
rect 562098 388046 562194 388102
rect 562250 388046 562318 388102
rect 562374 388046 562442 388102
rect 562498 388046 562566 388102
rect 562622 388046 562718 388102
rect 562098 387978 562718 388046
rect 562098 387922 562194 387978
rect 562250 387922 562318 387978
rect 562374 387922 562442 387978
rect 562498 387922 562566 387978
rect 562622 387922 562718 387978
rect 562098 370350 562718 387922
rect 562098 370294 562194 370350
rect 562250 370294 562318 370350
rect 562374 370294 562442 370350
rect 562498 370294 562566 370350
rect 562622 370294 562718 370350
rect 562098 370226 562718 370294
rect 562098 370170 562194 370226
rect 562250 370170 562318 370226
rect 562374 370170 562442 370226
rect 562498 370170 562566 370226
rect 562622 370170 562718 370226
rect 562098 370102 562718 370170
rect 562098 370046 562194 370102
rect 562250 370046 562318 370102
rect 562374 370046 562442 370102
rect 562498 370046 562566 370102
rect 562622 370046 562718 370102
rect 562098 369978 562718 370046
rect 562098 369922 562194 369978
rect 562250 369922 562318 369978
rect 562374 369922 562442 369978
rect 562498 369922 562566 369978
rect 562622 369922 562718 369978
rect 562098 352350 562718 369922
rect 589098 597212 589718 598268
rect 589098 597156 589194 597212
rect 589250 597156 589318 597212
rect 589374 597156 589442 597212
rect 589498 597156 589566 597212
rect 589622 597156 589718 597212
rect 589098 597088 589718 597156
rect 589098 597032 589194 597088
rect 589250 597032 589318 597088
rect 589374 597032 589442 597088
rect 589498 597032 589566 597088
rect 589622 597032 589718 597088
rect 589098 596964 589718 597032
rect 589098 596908 589194 596964
rect 589250 596908 589318 596964
rect 589374 596908 589442 596964
rect 589498 596908 589566 596964
rect 589622 596908 589718 596964
rect 589098 596840 589718 596908
rect 589098 596784 589194 596840
rect 589250 596784 589318 596840
rect 589374 596784 589442 596840
rect 589498 596784 589566 596840
rect 589622 596784 589718 596840
rect 589098 580350 589718 596784
rect 589098 580294 589194 580350
rect 589250 580294 589318 580350
rect 589374 580294 589442 580350
rect 589498 580294 589566 580350
rect 589622 580294 589718 580350
rect 589098 580226 589718 580294
rect 589098 580170 589194 580226
rect 589250 580170 589318 580226
rect 589374 580170 589442 580226
rect 589498 580170 589566 580226
rect 589622 580170 589718 580226
rect 589098 580102 589718 580170
rect 589098 580046 589194 580102
rect 589250 580046 589318 580102
rect 589374 580046 589442 580102
rect 589498 580046 589566 580102
rect 589622 580046 589718 580102
rect 589098 579978 589718 580046
rect 589098 579922 589194 579978
rect 589250 579922 589318 579978
rect 589374 579922 589442 579978
rect 589498 579922 589566 579978
rect 589622 579922 589718 579978
rect 589098 562350 589718 579922
rect 589098 562294 589194 562350
rect 589250 562294 589318 562350
rect 589374 562294 589442 562350
rect 589498 562294 589566 562350
rect 589622 562294 589718 562350
rect 589098 562226 589718 562294
rect 589098 562170 589194 562226
rect 589250 562170 589318 562226
rect 589374 562170 589442 562226
rect 589498 562170 589566 562226
rect 589622 562170 589718 562226
rect 592818 598172 593438 598268
rect 592818 598116 592914 598172
rect 592970 598116 593038 598172
rect 593094 598116 593162 598172
rect 593218 598116 593286 598172
rect 593342 598116 593438 598172
rect 592818 598048 593438 598116
rect 592818 597992 592914 598048
rect 592970 597992 593038 598048
rect 593094 597992 593162 598048
rect 593218 597992 593286 598048
rect 593342 597992 593438 598048
rect 592818 597924 593438 597992
rect 592818 597868 592914 597924
rect 592970 597868 593038 597924
rect 593094 597868 593162 597924
rect 593218 597868 593286 597924
rect 593342 597868 593438 597924
rect 592818 597800 593438 597868
rect 592818 597744 592914 597800
rect 592970 597744 593038 597800
rect 593094 597744 593162 597800
rect 593218 597744 593286 597800
rect 593342 597744 593438 597800
rect 592818 586350 593438 597744
rect 597360 598172 597980 598268
rect 597360 598116 597456 598172
rect 597512 598116 597580 598172
rect 597636 598116 597704 598172
rect 597760 598116 597828 598172
rect 597884 598116 597980 598172
rect 597360 598048 597980 598116
rect 597360 597992 597456 598048
rect 597512 597992 597580 598048
rect 597636 597992 597704 598048
rect 597760 597992 597828 598048
rect 597884 597992 597980 598048
rect 597360 597924 597980 597992
rect 597360 597868 597456 597924
rect 597512 597868 597580 597924
rect 597636 597868 597704 597924
rect 597760 597868 597828 597924
rect 597884 597868 597980 597924
rect 597360 597800 597980 597868
rect 597360 597744 597456 597800
rect 597512 597744 597580 597800
rect 597636 597744 597704 597800
rect 597760 597744 597828 597800
rect 597884 597744 597980 597800
rect 592818 586294 592914 586350
rect 592970 586294 593038 586350
rect 593094 586294 593162 586350
rect 593218 586294 593286 586350
rect 593342 586294 593438 586350
rect 592818 586226 593438 586294
rect 592818 586170 592914 586226
rect 592970 586170 593038 586226
rect 593094 586170 593162 586226
rect 593218 586170 593286 586226
rect 593342 586170 593438 586226
rect 592818 586102 593438 586170
rect 592818 586046 592914 586102
rect 592970 586046 593038 586102
rect 593094 586046 593162 586102
rect 593218 586046 593286 586102
rect 593342 586046 593438 586102
rect 592818 585978 593438 586046
rect 592818 585922 592914 585978
rect 592970 585922 593038 585978
rect 593094 585922 593162 585978
rect 593218 585922 593286 585978
rect 593342 585922 593438 585978
rect 592818 568350 593438 585922
rect 592818 568294 592914 568350
rect 592970 568294 593038 568350
rect 593094 568294 593162 568350
rect 593218 568294 593286 568350
rect 593342 568294 593438 568350
rect 592818 568226 593438 568294
rect 592818 568170 592914 568226
rect 592970 568170 593038 568226
rect 593094 568170 593162 568226
rect 593218 568170 593286 568226
rect 593342 568170 593438 568226
rect 592818 568102 593438 568170
rect 592818 568046 592914 568102
rect 592970 568046 593038 568102
rect 593094 568046 593162 568102
rect 593218 568046 593286 568102
rect 593342 568046 593438 568102
rect 592818 567978 593438 568046
rect 592818 567922 592914 567978
rect 592970 567922 593038 567978
rect 593094 567922 593162 567978
rect 593218 567922 593286 567978
rect 593342 567922 593438 567978
rect 589098 562102 589718 562170
rect 589098 562046 589194 562102
rect 589250 562046 589318 562102
rect 589374 562046 589442 562102
rect 589498 562046 589566 562102
rect 589622 562046 589718 562102
rect 589098 561978 589718 562046
rect 589098 561922 589194 561978
rect 589250 561922 589318 561978
rect 589374 561922 589442 561978
rect 589498 561922 589566 561978
rect 589622 561922 589718 561978
rect 589098 544350 589718 561922
rect 589098 544294 589194 544350
rect 589250 544294 589318 544350
rect 589374 544294 589442 544350
rect 589498 544294 589566 544350
rect 589622 544294 589718 544350
rect 589098 544226 589718 544294
rect 589098 544170 589194 544226
rect 589250 544170 589318 544226
rect 589374 544170 589442 544226
rect 589498 544170 589566 544226
rect 589622 544170 589718 544226
rect 589098 544102 589718 544170
rect 589098 544046 589194 544102
rect 589250 544046 589318 544102
rect 589374 544046 589442 544102
rect 589498 544046 589566 544102
rect 589622 544046 589718 544102
rect 589098 543978 589718 544046
rect 589098 543922 589194 543978
rect 589250 543922 589318 543978
rect 589374 543922 589442 543978
rect 589498 543922 589566 543978
rect 589622 543922 589718 543978
rect 589098 526350 589718 543922
rect 589098 526294 589194 526350
rect 589250 526294 589318 526350
rect 589374 526294 589442 526350
rect 589498 526294 589566 526350
rect 589622 526294 589718 526350
rect 589098 526226 589718 526294
rect 589098 526170 589194 526226
rect 589250 526170 589318 526226
rect 589374 526170 589442 526226
rect 589498 526170 589566 526226
rect 589622 526170 589718 526226
rect 589098 526102 589718 526170
rect 589098 526046 589194 526102
rect 589250 526046 589318 526102
rect 589374 526046 589442 526102
rect 589498 526046 589566 526102
rect 589622 526046 589718 526102
rect 589098 525978 589718 526046
rect 589098 525922 589194 525978
rect 589250 525922 589318 525978
rect 589374 525922 589442 525978
rect 589498 525922 589566 525978
rect 589622 525922 589718 525978
rect 589098 508350 589718 525922
rect 590716 562212 590772 562222
rect 590716 523348 590772 562156
rect 590716 523282 590772 523292
rect 592818 550350 593438 567922
rect 592818 550294 592914 550350
rect 592970 550294 593038 550350
rect 593094 550294 593162 550350
rect 593218 550294 593286 550350
rect 593342 550294 593438 550350
rect 592818 550226 593438 550294
rect 592818 550170 592914 550226
rect 592970 550170 593038 550226
rect 593094 550170 593162 550226
rect 593218 550170 593286 550226
rect 593342 550170 593438 550226
rect 592818 550102 593438 550170
rect 592818 550046 592914 550102
rect 592970 550046 593038 550102
rect 593094 550046 593162 550102
rect 593218 550046 593286 550102
rect 593342 550046 593438 550102
rect 592818 549978 593438 550046
rect 592818 549922 592914 549978
rect 592970 549922 593038 549978
rect 593094 549922 593162 549978
rect 593218 549922 593286 549978
rect 593342 549922 593438 549978
rect 592818 532350 593438 549922
rect 592818 532294 592914 532350
rect 592970 532294 593038 532350
rect 593094 532294 593162 532350
rect 593218 532294 593286 532350
rect 593342 532294 593438 532350
rect 592818 532226 593438 532294
rect 592818 532170 592914 532226
rect 592970 532170 593038 532226
rect 593094 532170 593162 532226
rect 593218 532170 593286 532226
rect 593342 532170 593438 532226
rect 592818 532102 593438 532170
rect 592818 532046 592914 532102
rect 592970 532046 593038 532102
rect 593094 532046 593162 532102
rect 593218 532046 593286 532102
rect 593342 532046 593438 532102
rect 592818 531978 593438 532046
rect 592818 531922 592914 531978
rect 592970 531922 593038 531978
rect 593094 531922 593162 531978
rect 593218 531922 593286 531978
rect 593342 531922 593438 531978
rect 589098 508294 589194 508350
rect 589250 508294 589318 508350
rect 589374 508294 589442 508350
rect 589498 508294 589566 508350
rect 589622 508294 589718 508350
rect 589098 508226 589718 508294
rect 589098 508170 589194 508226
rect 589250 508170 589318 508226
rect 589374 508170 589442 508226
rect 589498 508170 589566 508226
rect 589622 508170 589718 508226
rect 589098 508102 589718 508170
rect 589098 508046 589194 508102
rect 589250 508046 589318 508102
rect 589374 508046 589442 508102
rect 589498 508046 589566 508102
rect 589622 508046 589718 508102
rect 589098 507978 589718 508046
rect 589098 507922 589194 507978
rect 589250 507922 589318 507978
rect 589374 507922 589442 507978
rect 589498 507922 589566 507978
rect 589622 507922 589718 507978
rect 589098 490350 589718 507922
rect 590492 522564 590548 522574
rect 590156 496132 590212 496142
rect 590156 494788 590212 496076
rect 590156 494722 590212 494732
rect 589098 490294 589194 490350
rect 589250 490294 589318 490350
rect 589374 490294 589442 490350
rect 589498 490294 589566 490350
rect 589622 490294 589718 490350
rect 589098 490226 589718 490294
rect 589098 490170 589194 490226
rect 589250 490170 589318 490226
rect 589374 490170 589442 490226
rect 589498 490170 589566 490226
rect 589622 490170 589718 490226
rect 589098 490102 589718 490170
rect 589098 490046 589194 490102
rect 589250 490046 589318 490102
rect 589374 490046 589442 490102
rect 589498 490046 589566 490102
rect 589622 490046 589718 490102
rect 589098 489978 589718 490046
rect 589098 489922 589194 489978
rect 589250 489922 589318 489978
rect 589374 489922 589442 489978
rect 589498 489922 589566 489978
rect 589622 489922 589718 489978
rect 589098 472350 589718 489922
rect 589098 472294 589194 472350
rect 589250 472294 589318 472350
rect 589374 472294 589442 472350
rect 589498 472294 589566 472350
rect 589622 472294 589718 472350
rect 589098 472226 589718 472294
rect 589098 472170 589194 472226
rect 589250 472170 589318 472226
rect 589374 472170 589442 472226
rect 589498 472170 589566 472226
rect 589622 472170 589718 472226
rect 589098 472102 589718 472170
rect 589098 472046 589194 472102
rect 589250 472046 589318 472102
rect 589374 472046 589442 472102
rect 589498 472046 589566 472102
rect 589622 472046 589718 472102
rect 589098 471978 589718 472046
rect 589098 471922 589194 471978
rect 589250 471922 589318 471978
rect 589374 471922 589442 471978
rect 589498 471922 589566 471978
rect 589622 471922 589718 471978
rect 589098 454350 589718 471922
rect 589098 454294 589194 454350
rect 589250 454294 589318 454350
rect 589374 454294 589442 454350
rect 589498 454294 589566 454350
rect 589622 454294 589718 454350
rect 589098 454226 589718 454294
rect 589098 454170 589194 454226
rect 589250 454170 589318 454226
rect 589374 454170 589442 454226
rect 589498 454170 589566 454226
rect 589622 454170 589718 454226
rect 589098 454102 589718 454170
rect 589098 454046 589194 454102
rect 589250 454046 589318 454102
rect 589374 454046 589442 454102
rect 589498 454046 589566 454102
rect 589622 454046 589718 454102
rect 589098 453978 589718 454046
rect 589098 453922 589194 453978
rect 589250 453922 589318 453978
rect 589374 453922 589442 453978
rect 589498 453922 589566 453978
rect 589622 453922 589718 453978
rect 589098 436350 589718 453922
rect 589098 436294 589194 436350
rect 589250 436294 589318 436350
rect 589374 436294 589442 436350
rect 589498 436294 589566 436350
rect 589622 436294 589718 436350
rect 589098 436226 589718 436294
rect 589098 436170 589194 436226
rect 589250 436170 589318 436226
rect 589374 436170 589442 436226
rect 589498 436170 589566 436226
rect 589622 436170 589718 436226
rect 589098 436102 589718 436170
rect 589098 436046 589194 436102
rect 589250 436046 589318 436102
rect 589374 436046 589442 436102
rect 589498 436046 589566 436102
rect 589622 436046 589718 436102
rect 589098 435978 589718 436046
rect 589098 435922 589194 435978
rect 589250 435922 589318 435978
rect 589374 435922 589442 435978
rect 589498 435922 589566 435978
rect 589622 435922 589718 435978
rect 589098 418350 589718 435922
rect 589098 418294 589194 418350
rect 589250 418294 589318 418350
rect 589374 418294 589442 418350
rect 589498 418294 589566 418350
rect 589622 418294 589718 418350
rect 589098 418226 589718 418294
rect 589098 418170 589194 418226
rect 589250 418170 589318 418226
rect 589374 418170 589442 418226
rect 589498 418170 589566 418226
rect 589622 418170 589718 418226
rect 589098 418102 589718 418170
rect 589098 418046 589194 418102
rect 589250 418046 589318 418102
rect 589374 418046 589442 418102
rect 589498 418046 589566 418102
rect 589622 418046 589718 418102
rect 589098 417978 589718 418046
rect 589098 417922 589194 417978
rect 589250 417922 589318 417978
rect 589374 417922 589442 417978
rect 589498 417922 589566 417978
rect 589622 417922 589718 417978
rect 589098 400350 589718 417922
rect 589098 400294 589194 400350
rect 589250 400294 589318 400350
rect 589374 400294 589442 400350
rect 589498 400294 589566 400350
rect 589622 400294 589718 400350
rect 589098 400226 589718 400294
rect 589098 400170 589194 400226
rect 589250 400170 589318 400226
rect 589374 400170 589442 400226
rect 589498 400170 589566 400226
rect 589622 400170 589718 400226
rect 589098 400102 589718 400170
rect 589098 400046 589194 400102
rect 589250 400046 589318 400102
rect 589374 400046 589442 400102
rect 589498 400046 589566 400102
rect 589622 400046 589718 400102
rect 589098 399978 589718 400046
rect 589098 399922 589194 399978
rect 589250 399922 589318 399978
rect 589374 399922 589442 399978
rect 589498 399922 589566 399978
rect 589622 399922 589718 399978
rect 589098 382350 589718 399922
rect 589098 382294 589194 382350
rect 589250 382294 589318 382350
rect 589374 382294 589442 382350
rect 589498 382294 589566 382350
rect 589622 382294 589718 382350
rect 589098 382226 589718 382294
rect 589098 382170 589194 382226
rect 589250 382170 589318 382226
rect 589374 382170 589442 382226
rect 589498 382170 589566 382226
rect 589622 382170 589718 382226
rect 589098 382102 589718 382170
rect 589098 382046 589194 382102
rect 589250 382046 589318 382102
rect 589374 382046 589442 382102
rect 589498 382046 589566 382102
rect 589622 382046 589718 382102
rect 589098 381978 589718 382046
rect 589098 381922 589194 381978
rect 589250 381922 589318 381978
rect 589374 381922 589442 381978
rect 589498 381922 589566 381978
rect 589622 381922 589718 381978
rect 589098 364350 589718 381922
rect 589098 364294 589194 364350
rect 589250 364294 589318 364350
rect 589374 364294 589442 364350
rect 589498 364294 589566 364350
rect 589622 364294 589718 364350
rect 589098 364226 589718 364294
rect 589098 364170 589194 364226
rect 589250 364170 589318 364226
rect 589374 364170 589442 364226
rect 589498 364170 589566 364226
rect 589622 364170 589718 364226
rect 589098 364102 589718 364170
rect 589098 364046 589194 364102
rect 589250 364046 589318 364102
rect 589374 364046 589442 364102
rect 589498 364046 589566 364102
rect 589622 364046 589718 364102
rect 562098 352294 562194 352350
rect 562250 352294 562318 352350
rect 562374 352294 562442 352350
rect 562498 352294 562566 352350
rect 562622 352294 562718 352350
rect 562098 352226 562718 352294
rect 562098 352170 562194 352226
rect 562250 352170 562318 352226
rect 562374 352170 562442 352226
rect 562498 352170 562566 352226
rect 562622 352170 562718 352226
rect 562098 352102 562718 352170
rect 562098 352046 562194 352102
rect 562250 352046 562318 352102
rect 562374 352046 562442 352102
rect 562498 352046 562566 352102
rect 562622 352046 562718 352102
rect 562098 351978 562718 352046
rect 562098 351922 562194 351978
rect 562250 351922 562318 351978
rect 562374 351922 562442 351978
rect 562498 351922 562566 351978
rect 562622 351922 562718 351978
rect 562098 334350 562718 351922
rect 562098 334294 562194 334350
rect 562250 334294 562318 334350
rect 562374 334294 562442 334350
rect 562498 334294 562566 334350
rect 562622 334294 562718 334350
rect 562098 334226 562718 334294
rect 562098 334170 562194 334226
rect 562250 334170 562318 334226
rect 562374 334170 562442 334226
rect 562498 334170 562566 334226
rect 562622 334170 562718 334226
rect 562098 334102 562718 334170
rect 562098 334046 562194 334102
rect 562250 334046 562318 334102
rect 562374 334046 562442 334102
rect 562498 334046 562566 334102
rect 562622 334046 562718 334102
rect 562098 333978 562718 334046
rect 562098 333922 562194 333978
rect 562250 333922 562318 333978
rect 562374 333922 562442 333978
rect 562498 333922 562566 333978
rect 562622 333922 562718 333978
rect 562098 316350 562718 333922
rect 562098 316294 562194 316350
rect 562250 316294 562318 316350
rect 562374 316294 562442 316350
rect 562498 316294 562566 316350
rect 562622 316294 562718 316350
rect 562098 316226 562718 316294
rect 562098 316170 562194 316226
rect 562250 316170 562318 316226
rect 562374 316170 562442 316226
rect 562498 316170 562566 316226
rect 562622 316170 562718 316226
rect 562098 316102 562718 316170
rect 562098 316046 562194 316102
rect 562250 316046 562318 316102
rect 562374 316046 562442 316102
rect 562498 316046 562566 316102
rect 562622 316046 562718 316102
rect 562098 315978 562718 316046
rect 562098 315922 562194 315978
rect 562250 315922 562318 315978
rect 562374 315922 562442 315978
rect 562498 315922 562566 315978
rect 562622 315922 562718 315978
rect 562098 298350 562718 315922
rect 562098 298294 562194 298350
rect 562250 298294 562318 298350
rect 562374 298294 562442 298350
rect 562498 298294 562566 298350
rect 562622 298294 562718 298350
rect 562098 298226 562718 298294
rect 562098 298170 562194 298226
rect 562250 298170 562318 298226
rect 562374 298170 562442 298226
rect 562498 298170 562566 298226
rect 562622 298170 562718 298226
rect 562098 298102 562718 298170
rect 562098 298046 562194 298102
rect 562250 298046 562318 298102
rect 562374 298046 562442 298102
rect 562498 298046 562566 298102
rect 562622 298046 562718 298102
rect 562098 297978 562718 298046
rect 562098 297922 562194 297978
rect 562250 297922 562318 297978
rect 562374 297922 562442 297978
rect 562498 297922 562566 297978
rect 562622 297922 562718 297978
rect 562098 280350 562718 297922
rect 562098 280294 562194 280350
rect 562250 280294 562318 280350
rect 562374 280294 562442 280350
rect 562498 280294 562566 280350
rect 562622 280294 562718 280350
rect 562098 280226 562718 280294
rect 562098 280170 562194 280226
rect 562250 280170 562318 280226
rect 562374 280170 562442 280226
rect 562498 280170 562566 280226
rect 562622 280170 562718 280226
rect 562098 280102 562718 280170
rect 562098 280046 562194 280102
rect 562250 280046 562318 280102
rect 562374 280046 562442 280102
rect 562498 280046 562566 280102
rect 562622 280046 562718 280102
rect 562098 279978 562718 280046
rect 562098 279922 562194 279978
rect 562250 279922 562318 279978
rect 562374 279922 562442 279978
rect 562498 279922 562566 279978
rect 562622 279922 562718 279978
rect 562098 262350 562718 279922
rect 562098 262294 562194 262350
rect 562250 262294 562318 262350
rect 562374 262294 562442 262350
rect 562498 262294 562566 262350
rect 562622 262294 562718 262350
rect 562098 262226 562718 262294
rect 562098 262170 562194 262226
rect 562250 262170 562318 262226
rect 562374 262170 562442 262226
rect 562498 262170 562566 262226
rect 562622 262170 562718 262226
rect 562098 262102 562718 262170
rect 562098 262046 562194 262102
rect 562250 262046 562318 262102
rect 562374 262046 562442 262102
rect 562498 262046 562566 262102
rect 562622 262046 562718 262102
rect 562098 261978 562718 262046
rect 562098 261922 562194 261978
rect 562250 261922 562318 261978
rect 562374 261922 562442 261978
rect 562498 261922 562566 261978
rect 562622 261922 562718 261978
rect 562098 244350 562718 261922
rect 562098 244294 562194 244350
rect 562250 244294 562318 244350
rect 562374 244294 562442 244350
rect 562498 244294 562566 244350
rect 562622 244294 562718 244350
rect 562098 244226 562718 244294
rect 562098 244170 562194 244226
rect 562250 244170 562318 244226
rect 562374 244170 562442 244226
rect 562498 244170 562566 244226
rect 562622 244170 562718 244226
rect 562098 244102 562718 244170
rect 562098 244046 562194 244102
rect 562250 244046 562318 244102
rect 562374 244046 562442 244102
rect 562498 244046 562566 244102
rect 562622 244046 562718 244102
rect 562098 243978 562718 244046
rect 562098 243922 562194 243978
rect 562250 243922 562318 243978
rect 562374 243922 562442 243978
rect 562498 243922 562566 243978
rect 562622 243922 562718 243978
rect 562098 226350 562718 243922
rect 562098 226294 562194 226350
rect 562250 226294 562318 226350
rect 562374 226294 562442 226350
rect 562498 226294 562566 226350
rect 562622 226294 562718 226350
rect 562098 226226 562718 226294
rect 562098 226170 562194 226226
rect 562250 226170 562318 226226
rect 562374 226170 562442 226226
rect 562498 226170 562566 226226
rect 562622 226170 562718 226226
rect 562098 226102 562718 226170
rect 562098 226046 562194 226102
rect 562250 226046 562318 226102
rect 562374 226046 562442 226102
rect 562498 226046 562566 226102
rect 562622 226046 562718 226102
rect 562098 225978 562718 226046
rect 562098 225922 562194 225978
rect 562250 225922 562318 225978
rect 562374 225922 562442 225978
rect 562498 225922 562566 225978
rect 562622 225922 562718 225978
rect 562098 208350 562718 225922
rect 562098 208294 562194 208350
rect 562250 208294 562318 208350
rect 562374 208294 562442 208350
rect 562498 208294 562566 208350
rect 562622 208294 562718 208350
rect 562098 208226 562718 208294
rect 562098 208170 562194 208226
rect 562250 208170 562318 208226
rect 562374 208170 562442 208226
rect 562498 208170 562566 208226
rect 562622 208170 562718 208226
rect 562098 208102 562718 208170
rect 562098 208046 562194 208102
rect 562250 208046 562318 208102
rect 562374 208046 562442 208102
rect 562498 208046 562566 208102
rect 562622 208046 562718 208102
rect 562098 207978 562718 208046
rect 562098 207922 562194 207978
rect 562250 207922 562318 207978
rect 562374 207922 562442 207978
rect 562498 207922 562566 207978
rect 562622 207922 562718 207978
rect 562098 190350 562718 207922
rect 562098 190294 562194 190350
rect 562250 190294 562318 190350
rect 562374 190294 562442 190350
rect 562498 190294 562566 190350
rect 562622 190294 562718 190350
rect 562098 190226 562718 190294
rect 562098 190170 562194 190226
rect 562250 190170 562318 190226
rect 562374 190170 562442 190226
rect 562498 190170 562566 190226
rect 562622 190170 562718 190226
rect 562098 190102 562718 190170
rect 562098 190046 562194 190102
rect 562250 190046 562318 190102
rect 562374 190046 562442 190102
rect 562498 190046 562566 190102
rect 562622 190046 562718 190102
rect 562098 189978 562718 190046
rect 562098 189922 562194 189978
rect 562250 189922 562318 189978
rect 562374 189922 562442 189978
rect 562498 189922 562566 189978
rect 562622 189922 562718 189978
rect 562098 172350 562718 189922
rect 562098 172294 562194 172350
rect 562250 172294 562318 172350
rect 562374 172294 562442 172350
rect 562498 172294 562566 172350
rect 562622 172294 562718 172350
rect 562098 172226 562718 172294
rect 562098 172170 562194 172226
rect 562250 172170 562318 172226
rect 562374 172170 562442 172226
rect 562498 172170 562566 172226
rect 562622 172170 562718 172226
rect 562098 172102 562718 172170
rect 562098 172046 562194 172102
rect 562250 172046 562318 172102
rect 562374 172046 562442 172102
rect 562498 172046 562566 172102
rect 562622 172046 562718 172102
rect 562098 171978 562718 172046
rect 562098 171922 562194 171978
rect 562250 171922 562318 171978
rect 562374 171922 562442 171978
rect 562498 171922 562566 171978
rect 562622 171922 562718 171978
rect 562098 154350 562718 171922
rect 562098 154294 562194 154350
rect 562250 154294 562318 154350
rect 562374 154294 562442 154350
rect 562498 154294 562566 154350
rect 562622 154294 562718 154350
rect 562098 154226 562718 154294
rect 562098 154170 562194 154226
rect 562250 154170 562318 154226
rect 562374 154170 562442 154226
rect 562498 154170 562566 154226
rect 562622 154170 562718 154226
rect 562098 154102 562718 154170
rect 562098 154046 562194 154102
rect 562250 154046 562318 154102
rect 562374 154046 562442 154102
rect 562498 154046 562566 154102
rect 562622 154046 562718 154102
rect 562098 153978 562718 154046
rect 562098 153922 562194 153978
rect 562250 153922 562318 153978
rect 562374 153922 562442 153978
rect 562498 153922 562566 153978
rect 562622 153922 562718 153978
rect 562098 136350 562718 153922
rect 562098 136294 562194 136350
rect 562250 136294 562318 136350
rect 562374 136294 562442 136350
rect 562498 136294 562566 136350
rect 562622 136294 562718 136350
rect 562098 136226 562718 136294
rect 562098 136170 562194 136226
rect 562250 136170 562318 136226
rect 562374 136170 562442 136226
rect 562498 136170 562566 136226
rect 562622 136170 562718 136226
rect 562098 136102 562718 136170
rect 562098 136046 562194 136102
rect 562250 136046 562318 136102
rect 562374 136046 562442 136102
rect 562498 136046 562566 136102
rect 562622 136046 562718 136102
rect 562098 135978 562718 136046
rect 562098 135922 562194 135978
rect 562250 135922 562318 135978
rect 562374 135922 562442 135978
rect 562498 135922 562566 135978
rect 562622 135922 562718 135978
rect 562098 118350 562718 135922
rect 562098 118294 562194 118350
rect 562250 118294 562318 118350
rect 562374 118294 562442 118350
rect 562498 118294 562566 118350
rect 562622 118294 562718 118350
rect 562098 118226 562718 118294
rect 562098 118170 562194 118226
rect 562250 118170 562318 118226
rect 562374 118170 562442 118226
rect 562498 118170 562566 118226
rect 562622 118170 562718 118226
rect 562098 118102 562718 118170
rect 562098 118046 562194 118102
rect 562250 118046 562318 118102
rect 562374 118046 562442 118102
rect 562498 118046 562566 118102
rect 562622 118046 562718 118102
rect 562098 117978 562718 118046
rect 562098 117922 562194 117978
rect 562250 117922 562318 117978
rect 562374 117922 562442 117978
rect 562498 117922 562566 117978
rect 562622 117922 562718 117978
rect 562098 100350 562718 117922
rect 587132 363972 587188 363982
rect 587132 105028 587188 363916
rect 587132 104962 587188 104972
rect 589098 363978 589718 364046
rect 589098 363922 589194 363978
rect 589250 363922 589318 363978
rect 589374 363922 589442 363978
rect 589498 363922 589566 363978
rect 589622 363922 589718 363978
rect 589098 346350 589718 363922
rect 589098 346294 589194 346350
rect 589250 346294 589318 346350
rect 589374 346294 589442 346350
rect 589498 346294 589566 346350
rect 589622 346294 589718 346350
rect 589098 346226 589718 346294
rect 589098 346170 589194 346226
rect 589250 346170 589318 346226
rect 589374 346170 589442 346226
rect 589498 346170 589566 346226
rect 589622 346170 589718 346226
rect 589098 346102 589718 346170
rect 589098 346046 589194 346102
rect 589250 346046 589318 346102
rect 589374 346046 589442 346102
rect 589498 346046 589566 346102
rect 589622 346046 589718 346102
rect 589098 345978 589718 346046
rect 589098 345922 589194 345978
rect 589250 345922 589318 345978
rect 589374 345922 589442 345978
rect 589498 345922 589566 345978
rect 589622 345922 589718 345978
rect 589098 328350 589718 345922
rect 589098 328294 589194 328350
rect 589250 328294 589318 328350
rect 589374 328294 589442 328350
rect 589498 328294 589566 328350
rect 589622 328294 589718 328350
rect 589098 328226 589718 328294
rect 589098 328170 589194 328226
rect 589250 328170 589318 328226
rect 589374 328170 589442 328226
rect 589498 328170 589566 328226
rect 589622 328170 589718 328226
rect 589098 328102 589718 328170
rect 589098 328046 589194 328102
rect 589250 328046 589318 328102
rect 589374 328046 589442 328102
rect 589498 328046 589566 328102
rect 589622 328046 589718 328102
rect 589098 327978 589718 328046
rect 589098 327922 589194 327978
rect 589250 327922 589318 327978
rect 589374 327922 589442 327978
rect 589498 327922 589566 327978
rect 589622 327922 589718 327978
rect 589098 310350 589718 327922
rect 589098 310294 589194 310350
rect 589250 310294 589318 310350
rect 589374 310294 589442 310350
rect 589498 310294 589566 310350
rect 589622 310294 589718 310350
rect 589098 310226 589718 310294
rect 589098 310170 589194 310226
rect 589250 310170 589318 310226
rect 589374 310170 589442 310226
rect 589498 310170 589566 310226
rect 589622 310170 589718 310226
rect 589098 310102 589718 310170
rect 589098 310046 589194 310102
rect 589250 310046 589318 310102
rect 589374 310046 589442 310102
rect 589498 310046 589566 310102
rect 589622 310046 589718 310102
rect 589098 309978 589718 310046
rect 589098 309922 589194 309978
rect 589250 309922 589318 309978
rect 589374 309922 589442 309978
rect 589498 309922 589566 309978
rect 589622 309922 589718 309978
rect 589098 292350 589718 309922
rect 590156 297892 590212 297902
rect 590156 296548 590212 297836
rect 590156 296482 590212 296492
rect 589098 292294 589194 292350
rect 589250 292294 589318 292350
rect 589374 292294 589442 292350
rect 589498 292294 589566 292350
rect 589622 292294 589718 292350
rect 589098 292226 589718 292294
rect 589098 292170 589194 292226
rect 589250 292170 589318 292226
rect 589374 292170 589442 292226
rect 589498 292170 589566 292226
rect 589622 292170 589718 292226
rect 589098 292102 589718 292170
rect 589098 292046 589194 292102
rect 589250 292046 589318 292102
rect 589374 292046 589442 292102
rect 589498 292046 589566 292102
rect 589622 292046 589718 292102
rect 589098 291978 589718 292046
rect 589098 291922 589194 291978
rect 589250 291922 589318 291978
rect 589374 291922 589442 291978
rect 589498 291922 589566 291978
rect 589622 291922 589718 291978
rect 589098 274350 589718 291922
rect 589098 274294 589194 274350
rect 589250 274294 589318 274350
rect 589374 274294 589442 274350
rect 589498 274294 589566 274350
rect 589622 274294 589718 274350
rect 589098 274226 589718 274294
rect 589098 274170 589194 274226
rect 589250 274170 589318 274226
rect 589374 274170 589442 274226
rect 589498 274170 589566 274226
rect 589622 274170 589718 274226
rect 589098 274102 589718 274170
rect 589098 274046 589194 274102
rect 589250 274046 589318 274102
rect 589374 274046 589442 274102
rect 589498 274046 589566 274102
rect 589622 274046 589718 274102
rect 589098 273978 589718 274046
rect 589098 273922 589194 273978
rect 589250 273922 589318 273978
rect 589374 273922 589442 273978
rect 589498 273922 589566 273978
rect 589622 273922 589718 273978
rect 589098 256350 589718 273922
rect 589098 256294 589194 256350
rect 589250 256294 589318 256350
rect 589374 256294 589442 256350
rect 589498 256294 589566 256350
rect 589622 256294 589718 256350
rect 589098 256226 589718 256294
rect 589098 256170 589194 256226
rect 589250 256170 589318 256226
rect 589374 256170 589442 256226
rect 589498 256170 589566 256226
rect 589622 256170 589718 256226
rect 589098 256102 589718 256170
rect 589098 256046 589194 256102
rect 589250 256046 589318 256102
rect 589374 256046 589442 256102
rect 589498 256046 589566 256102
rect 589622 256046 589718 256102
rect 589098 255978 589718 256046
rect 589098 255922 589194 255978
rect 589250 255922 589318 255978
rect 589374 255922 589442 255978
rect 589498 255922 589566 255978
rect 589622 255922 589718 255978
rect 589098 238350 589718 255922
rect 589098 238294 589194 238350
rect 589250 238294 589318 238350
rect 589374 238294 589442 238350
rect 589498 238294 589566 238350
rect 589622 238294 589718 238350
rect 589098 238226 589718 238294
rect 589098 238170 589194 238226
rect 589250 238170 589318 238226
rect 589374 238170 589442 238226
rect 589498 238170 589566 238226
rect 589622 238170 589718 238226
rect 589098 238102 589718 238170
rect 589098 238046 589194 238102
rect 589250 238046 589318 238102
rect 589374 238046 589442 238102
rect 589498 238046 589566 238102
rect 589622 238046 589718 238102
rect 589098 237978 589718 238046
rect 589098 237922 589194 237978
rect 589250 237922 589318 237978
rect 589374 237922 589442 237978
rect 589498 237922 589566 237978
rect 589622 237922 589718 237978
rect 589098 220350 589718 237922
rect 589098 220294 589194 220350
rect 589250 220294 589318 220350
rect 589374 220294 589442 220350
rect 589498 220294 589566 220350
rect 589622 220294 589718 220350
rect 589098 220226 589718 220294
rect 589098 220170 589194 220226
rect 589250 220170 589318 220226
rect 589374 220170 589442 220226
rect 589498 220170 589566 220226
rect 589622 220170 589718 220226
rect 589098 220102 589718 220170
rect 589098 220046 589194 220102
rect 589250 220046 589318 220102
rect 589374 220046 589442 220102
rect 589498 220046 589566 220102
rect 589622 220046 589718 220102
rect 589098 219978 589718 220046
rect 589098 219922 589194 219978
rect 589250 219922 589318 219978
rect 589374 219922 589442 219978
rect 589498 219922 589566 219978
rect 589622 219922 589718 219978
rect 589098 202350 589718 219922
rect 589098 202294 589194 202350
rect 589250 202294 589318 202350
rect 589374 202294 589442 202350
rect 589498 202294 589566 202350
rect 589622 202294 589718 202350
rect 589098 202226 589718 202294
rect 589098 202170 589194 202226
rect 589250 202170 589318 202226
rect 589374 202170 589442 202226
rect 589498 202170 589566 202226
rect 589622 202170 589718 202226
rect 589098 202102 589718 202170
rect 589098 202046 589194 202102
rect 589250 202046 589318 202102
rect 589374 202046 589442 202102
rect 589498 202046 589566 202102
rect 589622 202046 589718 202102
rect 589098 201978 589718 202046
rect 589098 201922 589194 201978
rect 589250 201922 589318 201978
rect 589374 201922 589442 201978
rect 589498 201922 589566 201978
rect 589622 201922 589718 201978
rect 589098 184350 589718 201922
rect 589098 184294 589194 184350
rect 589250 184294 589318 184350
rect 589374 184294 589442 184350
rect 589498 184294 589566 184350
rect 589622 184294 589718 184350
rect 589098 184226 589718 184294
rect 589098 184170 589194 184226
rect 589250 184170 589318 184226
rect 589374 184170 589442 184226
rect 589498 184170 589566 184226
rect 589622 184170 589718 184226
rect 589098 184102 589718 184170
rect 589098 184046 589194 184102
rect 589250 184046 589318 184102
rect 589374 184046 589442 184102
rect 589498 184046 589566 184102
rect 589622 184046 589718 184102
rect 589098 183978 589718 184046
rect 589098 183922 589194 183978
rect 589250 183922 589318 183978
rect 589374 183922 589442 183978
rect 589498 183922 589566 183978
rect 589622 183922 589718 183978
rect 589098 166350 589718 183922
rect 589098 166294 589194 166350
rect 589250 166294 589318 166350
rect 589374 166294 589442 166350
rect 589498 166294 589566 166350
rect 589622 166294 589718 166350
rect 589098 166226 589718 166294
rect 589098 166170 589194 166226
rect 589250 166170 589318 166226
rect 589374 166170 589442 166226
rect 589498 166170 589566 166226
rect 589622 166170 589718 166226
rect 589098 166102 589718 166170
rect 589098 166046 589194 166102
rect 589250 166046 589318 166102
rect 589374 166046 589442 166102
rect 589498 166046 589566 166102
rect 589622 166046 589718 166102
rect 589098 165978 589718 166046
rect 589098 165922 589194 165978
rect 589250 165922 589318 165978
rect 589374 165922 589442 165978
rect 589498 165922 589566 165978
rect 589622 165922 589718 165978
rect 589098 148350 589718 165922
rect 590156 165732 590212 165742
rect 590156 163828 590212 165676
rect 590156 163762 590212 163772
rect 589098 148294 589194 148350
rect 589250 148294 589318 148350
rect 589374 148294 589442 148350
rect 589498 148294 589566 148350
rect 589622 148294 589718 148350
rect 589098 148226 589718 148294
rect 589098 148170 589194 148226
rect 589250 148170 589318 148226
rect 589374 148170 589442 148226
rect 589498 148170 589566 148226
rect 589622 148170 589718 148226
rect 589098 148102 589718 148170
rect 589098 148046 589194 148102
rect 589250 148046 589318 148102
rect 589374 148046 589442 148102
rect 589498 148046 589566 148102
rect 589622 148046 589718 148102
rect 589098 147978 589718 148046
rect 589098 147922 589194 147978
rect 589250 147922 589318 147978
rect 589374 147922 589442 147978
rect 589498 147922 589566 147978
rect 589622 147922 589718 147978
rect 589098 130350 589718 147922
rect 589098 130294 589194 130350
rect 589250 130294 589318 130350
rect 589374 130294 589442 130350
rect 589498 130294 589566 130350
rect 589622 130294 589718 130350
rect 589098 130226 589718 130294
rect 589098 130170 589194 130226
rect 589250 130170 589318 130226
rect 589374 130170 589442 130226
rect 589498 130170 589566 130226
rect 589622 130170 589718 130226
rect 589098 130102 589718 130170
rect 589098 130046 589194 130102
rect 589250 130046 589318 130102
rect 589374 130046 589442 130102
rect 589498 130046 589566 130102
rect 589622 130046 589718 130102
rect 589098 129978 589718 130046
rect 589098 129922 589194 129978
rect 589250 129922 589318 129978
rect 589374 129922 589442 129978
rect 589498 129922 589566 129978
rect 589622 129922 589718 129978
rect 589098 112350 589718 129922
rect 589098 112294 589194 112350
rect 589250 112294 589318 112350
rect 589374 112294 589442 112350
rect 589498 112294 589566 112350
rect 589622 112294 589718 112350
rect 589098 112226 589718 112294
rect 589098 112170 589194 112226
rect 589250 112170 589318 112226
rect 589374 112170 589442 112226
rect 589498 112170 589566 112226
rect 589622 112170 589718 112226
rect 589098 112102 589718 112170
rect 589098 112046 589194 112102
rect 589250 112046 589318 112102
rect 589374 112046 589442 112102
rect 589498 112046 589566 112102
rect 589622 112046 589718 112102
rect 589098 111978 589718 112046
rect 589098 111922 589194 111978
rect 589250 111922 589318 111978
rect 589374 111922 589442 111978
rect 589498 111922 589566 111978
rect 589622 111922 589718 111978
rect 562098 100294 562194 100350
rect 562250 100294 562318 100350
rect 562374 100294 562442 100350
rect 562498 100294 562566 100350
rect 562622 100294 562718 100350
rect 562098 100226 562718 100294
rect 562098 100170 562194 100226
rect 562250 100170 562318 100226
rect 562374 100170 562442 100226
rect 562498 100170 562566 100226
rect 562622 100170 562718 100226
rect 562098 100102 562718 100170
rect 562098 100046 562194 100102
rect 562250 100046 562318 100102
rect 562374 100046 562442 100102
rect 562498 100046 562566 100102
rect 562622 100046 562718 100102
rect 562098 99978 562718 100046
rect 562098 99922 562194 99978
rect 562250 99922 562318 99978
rect 562374 99922 562442 99978
rect 562498 99922 562566 99978
rect 562622 99922 562718 99978
rect 562098 82350 562718 99922
rect 562098 82294 562194 82350
rect 562250 82294 562318 82350
rect 562374 82294 562442 82350
rect 562498 82294 562566 82350
rect 562622 82294 562718 82350
rect 562098 82226 562718 82294
rect 562098 82170 562194 82226
rect 562250 82170 562318 82226
rect 562374 82170 562442 82226
rect 562498 82170 562566 82226
rect 562622 82170 562718 82226
rect 562098 82102 562718 82170
rect 562098 82046 562194 82102
rect 562250 82046 562318 82102
rect 562374 82046 562442 82102
rect 562498 82046 562566 82102
rect 562622 82046 562718 82102
rect 562098 81978 562718 82046
rect 562098 81922 562194 81978
rect 562250 81922 562318 81978
rect 562374 81922 562442 81978
rect 562498 81922 562566 81978
rect 562622 81922 562718 81978
rect 562098 64350 562718 81922
rect 589098 94350 589718 111922
rect 590156 99652 590212 99662
rect 590156 98308 590212 99596
rect 590156 98242 590212 98252
rect 589098 94294 589194 94350
rect 589250 94294 589318 94350
rect 589374 94294 589442 94350
rect 589498 94294 589566 94350
rect 589622 94294 589718 94350
rect 589098 94226 589718 94294
rect 589098 94170 589194 94226
rect 589250 94170 589318 94226
rect 589374 94170 589442 94226
rect 589498 94170 589566 94226
rect 589622 94170 589718 94226
rect 589098 94102 589718 94170
rect 589098 94046 589194 94102
rect 589250 94046 589318 94102
rect 589374 94046 589442 94102
rect 589498 94046 589566 94102
rect 589622 94046 589718 94102
rect 589098 93978 589718 94046
rect 589098 93922 589194 93978
rect 589250 93922 589318 93978
rect 589374 93922 589442 93978
rect 589498 93922 589566 93978
rect 589622 93922 589718 93978
rect 589098 76350 589718 93922
rect 590492 78058 590548 522508
rect 592818 514350 593438 531922
rect 592818 514294 592914 514350
rect 592970 514294 593038 514350
rect 593094 514294 593162 514350
rect 593218 514294 593286 514350
rect 593342 514294 593438 514350
rect 592818 514226 593438 514294
rect 592818 514170 592914 514226
rect 592970 514170 593038 514226
rect 593094 514170 593162 514226
rect 593218 514170 593286 514226
rect 593342 514170 593438 514226
rect 592818 514102 593438 514170
rect 592818 514046 592914 514102
rect 592970 514046 593038 514102
rect 593094 514046 593162 514102
rect 593218 514046 593286 514102
rect 593342 514046 593438 514102
rect 592818 513978 593438 514046
rect 592818 513922 592914 513978
rect 592970 513922 593038 513978
rect 593094 513922 593162 513978
rect 593218 513922 593286 513978
rect 593342 513922 593438 513978
rect 592818 496350 593438 513922
rect 592818 496294 592914 496350
rect 592970 496294 593038 496350
rect 593094 496294 593162 496350
rect 593218 496294 593286 496350
rect 593342 496294 593438 496350
rect 592818 496226 593438 496294
rect 592818 496170 592914 496226
rect 592970 496170 593038 496226
rect 593094 496170 593162 496226
rect 593218 496170 593286 496226
rect 593342 496170 593438 496226
rect 592818 496102 593438 496170
rect 592818 496046 592914 496102
rect 592970 496046 593038 496102
rect 593094 496046 593162 496102
rect 593218 496046 593286 496102
rect 593342 496046 593438 496102
rect 592818 495978 593438 496046
rect 592818 495922 592914 495978
rect 592970 495922 593038 495978
rect 593094 495922 593162 495978
rect 593218 495922 593286 495978
rect 593342 495922 593438 495978
rect 592818 478350 593438 495922
rect 592818 478294 592914 478350
rect 592970 478294 593038 478350
rect 593094 478294 593162 478350
rect 593218 478294 593286 478350
rect 593342 478294 593438 478350
rect 592818 478226 593438 478294
rect 592818 478170 592914 478226
rect 592970 478170 593038 478226
rect 593094 478170 593162 478226
rect 593218 478170 593286 478226
rect 593342 478170 593438 478226
rect 592818 478102 593438 478170
rect 592818 478046 592914 478102
rect 592970 478046 593038 478102
rect 593094 478046 593162 478102
rect 593218 478046 593286 478102
rect 593342 478046 593438 478102
rect 592818 477978 593438 478046
rect 592818 477922 592914 477978
rect 592970 477922 593038 477978
rect 593094 477922 593162 477978
rect 593218 477922 593286 477978
rect 593342 477922 593438 477978
rect 592818 460350 593438 477922
rect 592818 460294 592914 460350
rect 592970 460294 593038 460350
rect 593094 460294 593162 460350
rect 593218 460294 593286 460350
rect 593342 460294 593438 460350
rect 592818 460226 593438 460294
rect 592818 460170 592914 460226
rect 592970 460170 593038 460226
rect 593094 460170 593162 460226
rect 593218 460170 593286 460226
rect 593342 460170 593438 460226
rect 592818 460102 593438 460170
rect 592818 460046 592914 460102
rect 592970 460046 593038 460102
rect 593094 460046 593162 460102
rect 593218 460046 593286 460102
rect 593342 460046 593438 460102
rect 592818 459978 593438 460046
rect 592818 459922 592914 459978
rect 592970 459922 593038 459978
rect 593094 459922 593162 459978
rect 593218 459922 593286 459978
rect 593342 459922 593438 459978
rect 592818 442350 593438 459922
rect 592818 442294 592914 442350
rect 592970 442294 593038 442350
rect 593094 442294 593162 442350
rect 593218 442294 593286 442350
rect 593342 442294 593438 442350
rect 592818 442226 593438 442294
rect 592818 442170 592914 442226
rect 592970 442170 593038 442226
rect 593094 442170 593162 442226
rect 593218 442170 593286 442226
rect 593342 442170 593438 442226
rect 592818 442102 593438 442170
rect 592818 442046 592914 442102
rect 592970 442046 593038 442102
rect 593094 442046 593162 442102
rect 593218 442046 593286 442102
rect 593342 442046 593438 442102
rect 592818 441978 593438 442046
rect 592818 441922 592914 441978
rect 592970 441922 593038 441978
rect 593094 441922 593162 441978
rect 593218 441922 593286 441978
rect 593342 441922 593438 441978
rect 592818 424350 593438 441922
rect 592818 424294 592914 424350
rect 592970 424294 593038 424350
rect 593094 424294 593162 424350
rect 593218 424294 593286 424350
rect 593342 424294 593438 424350
rect 592818 424226 593438 424294
rect 592818 424170 592914 424226
rect 592970 424170 593038 424226
rect 593094 424170 593162 424226
rect 593218 424170 593286 424226
rect 593342 424170 593438 424226
rect 592818 424102 593438 424170
rect 592818 424046 592914 424102
rect 592970 424046 593038 424102
rect 593094 424046 593162 424102
rect 593218 424046 593286 424102
rect 593342 424046 593438 424102
rect 592818 423978 593438 424046
rect 592818 423922 592914 423978
rect 592970 423922 593038 423978
rect 593094 423922 593162 423978
rect 593218 423922 593286 423978
rect 593342 423922 593438 423978
rect 592818 406350 593438 423922
rect 592818 406294 592914 406350
rect 592970 406294 593038 406350
rect 593094 406294 593162 406350
rect 593218 406294 593286 406350
rect 593342 406294 593438 406350
rect 592818 406226 593438 406294
rect 592818 406170 592914 406226
rect 592970 406170 593038 406226
rect 593094 406170 593162 406226
rect 593218 406170 593286 406226
rect 593342 406170 593438 406226
rect 592818 406102 593438 406170
rect 592818 406046 592914 406102
rect 592970 406046 593038 406102
rect 593094 406046 593162 406102
rect 593218 406046 593286 406102
rect 593342 406046 593438 406102
rect 592818 405978 593438 406046
rect 592818 405922 592914 405978
rect 592970 405922 593038 405978
rect 593094 405922 593162 405978
rect 593218 405922 593286 405978
rect 593342 405922 593438 405978
rect 592818 388350 593438 405922
rect 592818 388294 592914 388350
rect 592970 388294 593038 388350
rect 593094 388294 593162 388350
rect 593218 388294 593286 388350
rect 593342 388294 593438 388350
rect 592818 388226 593438 388294
rect 592818 388170 592914 388226
rect 592970 388170 593038 388226
rect 593094 388170 593162 388226
rect 593218 388170 593286 388226
rect 593342 388170 593438 388226
rect 592818 388102 593438 388170
rect 592818 388046 592914 388102
rect 592970 388046 593038 388102
rect 593094 388046 593162 388102
rect 593218 388046 593286 388102
rect 593342 388046 593438 388102
rect 592818 387978 593438 388046
rect 592818 387922 592914 387978
rect 592970 387922 593038 387978
rect 593094 387922 593162 387978
rect 593218 387922 593286 387978
rect 593342 387922 593438 387978
rect 592818 370350 593438 387922
rect 592818 370294 592914 370350
rect 592970 370294 593038 370350
rect 593094 370294 593162 370350
rect 593218 370294 593286 370350
rect 593342 370294 593438 370350
rect 592818 370226 593438 370294
rect 592818 370170 592914 370226
rect 592970 370170 593038 370226
rect 593094 370170 593162 370226
rect 593218 370170 593286 370226
rect 593342 370170 593438 370226
rect 592818 370102 593438 370170
rect 592818 370046 592914 370102
rect 592970 370046 593038 370102
rect 593094 370046 593162 370102
rect 593218 370046 593286 370102
rect 593342 370046 593438 370102
rect 592818 369978 593438 370046
rect 592818 369922 592914 369978
rect 592970 369922 593038 369978
rect 593094 369922 593162 369978
rect 593218 369922 593286 369978
rect 593342 369922 593438 369978
rect 592818 352350 593438 369922
rect 592818 352294 592914 352350
rect 592970 352294 593038 352350
rect 593094 352294 593162 352350
rect 593218 352294 593286 352350
rect 593342 352294 593438 352350
rect 592818 352226 593438 352294
rect 592818 352170 592914 352226
rect 592970 352170 593038 352226
rect 593094 352170 593162 352226
rect 593218 352170 593286 352226
rect 593342 352170 593438 352226
rect 592818 352102 593438 352170
rect 592818 352046 592914 352102
rect 592970 352046 593038 352102
rect 593094 352046 593162 352102
rect 593218 352046 593286 352102
rect 593342 352046 593438 352102
rect 592818 351978 593438 352046
rect 592818 351922 592914 351978
rect 592970 351922 593038 351978
rect 593094 351922 593162 351978
rect 593218 351922 593286 351978
rect 593342 351922 593438 351978
rect 592818 334350 593438 351922
rect 592818 334294 592914 334350
rect 592970 334294 593038 334350
rect 593094 334294 593162 334350
rect 593218 334294 593286 334350
rect 593342 334294 593438 334350
rect 592818 334226 593438 334294
rect 592818 334170 592914 334226
rect 592970 334170 593038 334226
rect 593094 334170 593162 334226
rect 593218 334170 593286 334226
rect 593342 334170 593438 334226
rect 592818 334102 593438 334170
rect 592818 334046 592914 334102
rect 592970 334046 593038 334102
rect 593094 334046 593162 334102
rect 593218 334046 593286 334102
rect 593342 334046 593438 334102
rect 592818 333978 593438 334046
rect 592818 333922 592914 333978
rect 592970 333922 593038 333978
rect 593094 333922 593162 333978
rect 593218 333922 593286 333978
rect 593342 333922 593438 333978
rect 592818 316350 593438 333922
rect 592818 316294 592914 316350
rect 592970 316294 593038 316350
rect 593094 316294 593162 316350
rect 593218 316294 593286 316350
rect 593342 316294 593438 316350
rect 592818 316226 593438 316294
rect 592818 316170 592914 316226
rect 592970 316170 593038 316226
rect 593094 316170 593162 316226
rect 593218 316170 593286 316226
rect 593342 316170 593438 316226
rect 592818 316102 593438 316170
rect 592818 316046 592914 316102
rect 592970 316046 593038 316102
rect 593094 316046 593162 316102
rect 593218 316046 593286 316102
rect 593342 316046 593438 316102
rect 592818 315978 593438 316046
rect 592818 315922 592914 315978
rect 592970 315922 593038 315978
rect 593094 315922 593162 315978
rect 593218 315922 593286 315978
rect 593342 315922 593438 315978
rect 592818 298350 593438 315922
rect 592818 298294 592914 298350
rect 592970 298294 593038 298350
rect 593094 298294 593162 298350
rect 593218 298294 593286 298350
rect 593342 298294 593438 298350
rect 592818 298226 593438 298294
rect 592818 298170 592914 298226
rect 592970 298170 593038 298226
rect 593094 298170 593162 298226
rect 593218 298170 593286 298226
rect 593342 298170 593438 298226
rect 592818 298102 593438 298170
rect 592818 298046 592914 298102
rect 592970 298046 593038 298102
rect 593094 298046 593162 298102
rect 593218 298046 593286 298102
rect 593342 298046 593438 298102
rect 592818 297978 593438 298046
rect 592818 297922 592914 297978
rect 592970 297922 593038 297978
rect 593094 297922 593162 297978
rect 593218 297922 593286 297978
rect 593342 297922 593438 297978
rect 592818 280350 593438 297922
rect 592818 280294 592914 280350
rect 592970 280294 593038 280350
rect 593094 280294 593162 280350
rect 593218 280294 593286 280350
rect 593342 280294 593438 280350
rect 592818 280226 593438 280294
rect 592818 280170 592914 280226
rect 592970 280170 593038 280226
rect 593094 280170 593162 280226
rect 593218 280170 593286 280226
rect 593342 280170 593438 280226
rect 592818 280102 593438 280170
rect 592818 280046 592914 280102
rect 592970 280046 593038 280102
rect 593094 280046 593162 280102
rect 593218 280046 593286 280102
rect 593342 280046 593438 280102
rect 592818 279978 593438 280046
rect 592818 279922 592914 279978
rect 592970 279922 593038 279978
rect 593094 279922 593162 279978
rect 593218 279922 593286 279978
rect 593342 279922 593438 279978
rect 592818 262350 593438 279922
rect 592818 262294 592914 262350
rect 592970 262294 593038 262350
rect 593094 262294 593162 262350
rect 593218 262294 593286 262350
rect 593342 262294 593438 262350
rect 592818 262226 593438 262294
rect 592818 262170 592914 262226
rect 592970 262170 593038 262226
rect 593094 262170 593162 262226
rect 593218 262170 593286 262226
rect 593342 262170 593438 262226
rect 592818 262102 593438 262170
rect 592818 262046 592914 262102
rect 592970 262046 593038 262102
rect 593094 262046 593162 262102
rect 593218 262046 593286 262102
rect 593342 262046 593438 262102
rect 592818 261978 593438 262046
rect 592818 261922 592914 261978
rect 592970 261922 593038 261978
rect 593094 261922 593162 261978
rect 593218 261922 593286 261978
rect 593342 261922 593438 261978
rect 591276 245028 591332 245038
rect 591276 242788 591332 244972
rect 591276 242722 591332 242732
rect 592818 244350 593438 261922
rect 592818 244294 592914 244350
rect 592970 244294 593038 244350
rect 593094 244294 593162 244350
rect 593218 244294 593286 244350
rect 593342 244294 593438 244350
rect 592818 244226 593438 244294
rect 592818 244170 592914 244226
rect 592970 244170 593038 244226
rect 593094 244170 593162 244226
rect 593218 244170 593286 244226
rect 593342 244170 593438 244226
rect 592818 244102 593438 244170
rect 592818 244046 592914 244102
rect 592970 244046 593038 244102
rect 593094 244046 593162 244102
rect 593218 244046 593286 244102
rect 593342 244046 593438 244102
rect 592818 243978 593438 244046
rect 592818 243922 592914 243978
rect 592970 243922 593038 243978
rect 593094 243922 593162 243978
rect 593218 243922 593286 243978
rect 593342 243922 593438 243978
rect 590492 77992 590548 78002
rect 592818 226350 593438 243922
rect 592818 226294 592914 226350
rect 592970 226294 593038 226350
rect 593094 226294 593162 226350
rect 593218 226294 593286 226350
rect 593342 226294 593438 226350
rect 592818 226226 593438 226294
rect 592818 226170 592914 226226
rect 592970 226170 593038 226226
rect 593094 226170 593162 226226
rect 593218 226170 593286 226226
rect 593342 226170 593438 226226
rect 592818 226102 593438 226170
rect 592818 226046 592914 226102
rect 592970 226046 593038 226102
rect 593094 226046 593162 226102
rect 593218 226046 593286 226102
rect 593342 226046 593438 226102
rect 592818 225978 593438 226046
rect 592818 225922 592914 225978
rect 592970 225922 593038 225978
rect 593094 225922 593162 225978
rect 593218 225922 593286 225978
rect 593342 225922 593438 225978
rect 592818 208350 593438 225922
rect 592818 208294 592914 208350
rect 592970 208294 593038 208350
rect 593094 208294 593162 208350
rect 593218 208294 593286 208350
rect 593342 208294 593438 208350
rect 592818 208226 593438 208294
rect 592818 208170 592914 208226
rect 592970 208170 593038 208226
rect 593094 208170 593162 208226
rect 593218 208170 593286 208226
rect 593342 208170 593438 208226
rect 592818 208102 593438 208170
rect 592818 208046 592914 208102
rect 592970 208046 593038 208102
rect 593094 208046 593162 208102
rect 593218 208046 593286 208102
rect 593342 208046 593438 208102
rect 592818 207978 593438 208046
rect 592818 207922 592914 207978
rect 592970 207922 593038 207978
rect 593094 207922 593162 207978
rect 593218 207922 593286 207978
rect 593342 207922 593438 207978
rect 592818 190350 593438 207922
rect 592818 190294 592914 190350
rect 592970 190294 593038 190350
rect 593094 190294 593162 190350
rect 593218 190294 593286 190350
rect 593342 190294 593438 190350
rect 592818 190226 593438 190294
rect 592818 190170 592914 190226
rect 592970 190170 593038 190226
rect 593094 190170 593162 190226
rect 593218 190170 593286 190226
rect 593342 190170 593438 190226
rect 592818 190102 593438 190170
rect 592818 190046 592914 190102
rect 592970 190046 593038 190102
rect 593094 190046 593162 190102
rect 593218 190046 593286 190102
rect 593342 190046 593438 190102
rect 592818 189978 593438 190046
rect 592818 189922 592914 189978
rect 592970 189922 593038 189978
rect 593094 189922 593162 189978
rect 593218 189922 593286 189978
rect 593342 189922 593438 189978
rect 592818 172350 593438 189922
rect 592818 172294 592914 172350
rect 592970 172294 593038 172350
rect 593094 172294 593162 172350
rect 593218 172294 593286 172350
rect 593342 172294 593438 172350
rect 592818 172226 593438 172294
rect 592818 172170 592914 172226
rect 592970 172170 593038 172226
rect 593094 172170 593162 172226
rect 593218 172170 593286 172226
rect 593342 172170 593438 172226
rect 592818 172102 593438 172170
rect 592818 172046 592914 172102
rect 592970 172046 593038 172102
rect 593094 172046 593162 172102
rect 593218 172046 593286 172102
rect 593342 172046 593438 172102
rect 592818 171978 593438 172046
rect 592818 171922 592914 171978
rect 592970 171922 593038 171978
rect 593094 171922 593162 171978
rect 593218 171922 593286 171978
rect 593342 171922 593438 171978
rect 592818 154350 593438 171922
rect 592818 154294 592914 154350
rect 592970 154294 593038 154350
rect 593094 154294 593162 154350
rect 593218 154294 593286 154350
rect 593342 154294 593438 154350
rect 592818 154226 593438 154294
rect 592818 154170 592914 154226
rect 592970 154170 593038 154226
rect 593094 154170 593162 154226
rect 593218 154170 593286 154226
rect 593342 154170 593438 154226
rect 592818 154102 593438 154170
rect 592818 154046 592914 154102
rect 592970 154046 593038 154102
rect 593094 154046 593162 154102
rect 593218 154046 593286 154102
rect 593342 154046 593438 154102
rect 592818 153978 593438 154046
rect 592818 153922 592914 153978
rect 592970 153922 593038 153978
rect 593094 153922 593162 153978
rect 593218 153922 593286 153978
rect 593342 153922 593438 153978
rect 592818 136350 593438 153922
rect 592818 136294 592914 136350
rect 592970 136294 593038 136350
rect 593094 136294 593162 136350
rect 593218 136294 593286 136350
rect 593342 136294 593438 136350
rect 592818 136226 593438 136294
rect 592818 136170 592914 136226
rect 592970 136170 593038 136226
rect 593094 136170 593162 136226
rect 593218 136170 593286 136226
rect 593342 136170 593438 136226
rect 592818 136102 593438 136170
rect 592818 136046 592914 136102
rect 592970 136046 593038 136102
rect 593094 136046 593162 136102
rect 593218 136046 593286 136102
rect 593342 136046 593438 136102
rect 592818 135978 593438 136046
rect 592818 135922 592914 135978
rect 592970 135922 593038 135978
rect 593094 135922 593162 135978
rect 593218 135922 593286 135978
rect 593342 135922 593438 135978
rect 592818 118350 593438 135922
rect 592818 118294 592914 118350
rect 592970 118294 593038 118350
rect 593094 118294 593162 118350
rect 593218 118294 593286 118350
rect 593342 118294 593438 118350
rect 592818 118226 593438 118294
rect 592818 118170 592914 118226
rect 592970 118170 593038 118226
rect 593094 118170 593162 118226
rect 593218 118170 593286 118226
rect 593342 118170 593438 118226
rect 592818 118102 593438 118170
rect 592818 118046 592914 118102
rect 592970 118046 593038 118102
rect 593094 118046 593162 118102
rect 593218 118046 593286 118102
rect 593342 118046 593438 118102
rect 592818 117978 593438 118046
rect 592818 117922 592914 117978
rect 592970 117922 593038 117978
rect 593094 117922 593162 117978
rect 593218 117922 593286 117978
rect 593342 117922 593438 117978
rect 592818 100350 593438 117922
rect 592818 100294 592914 100350
rect 592970 100294 593038 100350
rect 593094 100294 593162 100350
rect 593218 100294 593286 100350
rect 593342 100294 593438 100350
rect 592818 100226 593438 100294
rect 592818 100170 592914 100226
rect 592970 100170 593038 100226
rect 593094 100170 593162 100226
rect 593218 100170 593286 100226
rect 593342 100170 593438 100226
rect 592818 100102 593438 100170
rect 592818 100046 592914 100102
rect 592970 100046 593038 100102
rect 593094 100046 593162 100102
rect 593218 100046 593286 100102
rect 593342 100046 593438 100102
rect 592818 99978 593438 100046
rect 592818 99922 592914 99978
rect 592970 99922 593038 99978
rect 593094 99922 593162 99978
rect 593218 99922 593286 99978
rect 593342 99922 593438 99978
rect 592818 82350 593438 99922
rect 592818 82294 592914 82350
rect 592970 82294 593038 82350
rect 593094 82294 593162 82350
rect 593218 82294 593286 82350
rect 593342 82294 593438 82350
rect 592818 82226 593438 82294
rect 592818 82170 592914 82226
rect 592970 82170 593038 82226
rect 593094 82170 593162 82226
rect 593218 82170 593286 82226
rect 593342 82170 593438 82226
rect 592818 82102 593438 82170
rect 592818 82046 592914 82102
rect 592970 82046 593038 82102
rect 593094 82046 593162 82102
rect 593218 82046 593286 82102
rect 593342 82046 593438 82102
rect 592818 81978 593438 82046
rect 592818 81922 592914 81978
rect 592970 81922 593038 81978
rect 593094 81922 593162 81978
rect 593218 81922 593286 81978
rect 593342 81922 593438 81978
rect 589098 76294 589194 76350
rect 589250 76294 589318 76350
rect 589374 76294 589442 76350
rect 589498 76294 589566 76350
rect 589622 76294 589718 76350
rect 589098 76226 589718 76294
rect 589098 76170 589194 76226
rect 589250 76170 589318 76226
rect 589374 76170 589442 76226
rect 589498 76170 589566 76226
rect 589622 76170 589718 76226
rect 589098 76102 589718 76170
rect 589098 76046 589194 76102
rect 589250 76046 589318 76102
rect 589374 76046 589442 76102
rect 589498 76046 589566 76102
rect 589622 76046 589718 76102
rect 589098 75978 589718 76046
rect 589098 75922 589194 75978
rect 589250 75922 589318 75978
rect 589374 75922 589442 75978
rect 589498 75922 589566 75978
rect 589622 75922 589718 75978
rect 562098 64294 562194 64350
rect 562250 64294 562318 64350
rect 562374 64294 562442 64350
rect 562498 64294 562566 64350
rect 562622 64294 562718 64350
rect 562098 64226 562718 64294
rect 562098 64170 562194 64226
rect 562250 64170 562318 64226
rect 562374 64170 562442 64226
rect 562498 64170 562566 64226
rect 562622 64170 562718 64226
rect 562098 64102 562718 64170
rect 562098 64046 562194 64102
rect 562250 64046 562318 64102
rect 562374 64046 562442 64102
rect 562498 64046 562566 64102
rect 562622 64046 562718 64102
rect 562098 63978 562718 64046
rect 562098 63922 562194 63978
rect 562250 63922 562318 63978
rect 562374 63922 562442 63978
rect 562498 63922 562566 63978
rect 562622 63922 562718 63978
rect 558378 40294 558474 40350
rect 558530 40294 558598 40350
rect 558654 40294 558722 40350
rect 558778 40294 558846 40350
rect 558902 40294 558998 40350
rect 558378 40226 558998 40294
rect 558378 40170 558474 40226
rect 558530 40170 558598 40226
rect 558654 40170 558722 40226
rect 558778 40170 558846 40226
rect 558902 40170 558998 40226
rect 558378 40102 558998 40170
rect 558378 40046 558474 40102
rect 558530 40046 558598 40102
rect 558654 40046 558722 40102
rect 558778 40046 558846 40102
rect 558902 40046 558998 40102
rect 558378 39978 558998 40046
rect 558378 39922 558474 39978
rect 558530 39922 558598 39978
rect 558654 39922 558722 39978
rect 558778 39922 558846 39978
rect 558902 39922 558998 39978
rect 558378 22350 558998 39922
rect 558378 22294 558474 22350
rect 558530 22294 558598 22350
rect 558654 22294 558722 22350
rect 558778 22294 558846 22350
rect 558902 22294 558998 22350
rect 558378 22226 558998 22294
rect 558378 22170 558474 22226
rect 558530 22170 558598 22226
rect 558654 22170 558722 22226
rect 558778 22170 558846 22226
rect 558902 22170 558998 22226
rect 558378 22102 558998 22170
rect 558378 22046 558474 22102
rect 558530 22046 558598 22102
rect 558654 22046 558722 22102
rect 558778 22046 558846 22102
rect 558902 22046 558998 22102
rect 558378 21978 558998 22046
rect 558378 21922 558474 21978
rect 558530 21922 558598 21978
rect 558654 21922 558722 21978
rect 558778 21922 558846 21978
rect 558902 21922 558998 21978
rect 558378 4350 558998 21922
rect 558378 4294 558474 4350
rect 558530 4294 558598 4350
rect 558654 4294 558722 4350
rect 558778 4294 558846 4350
rect 558902 4294 558998 4350
rect 558378 4226 558998 4294
rect 558378 4170 558474 4226
rect 558530 4170 558598 4226
rect 558654 4170 558722 4226
rect 558778 4170 558846 4226
rect 558902 4170 558998 4226
rect 558378 4102 558998 4170
rect 561148 55558 561204 55568
rect 561148 4228 561204 55502
rect 561148 4162 561204 4172
rect 562098 46350 562718 63922
rect 572908 67258 572964 67268
rect 562098 46294 562194 46350
rect 562250 46294 562318 46350
rect 562374 46294 562442 46350
rect 562498 46294 562566 46350
rect 562622 46294 562718 46350
rect 562098 46226 562718 46294
rect 562098 46170 562194 46226
rect 562250 46170 562318 46226
rect 562374 46170 562442 46226
rect 562498 46170 562566 46226
rect 562622 46170 562718 46226
rect 562098 46102 562718 46170
rect 562098 46046 562194 46102
rect 562250 46046 562318 46102
rect 562374 46046 562442 46102
rect 562498 46046 562566 46102
rect 562622 46046 562718 46102
rect 562098 45978 562718 46046
rect 562098 45922 562194 45978
rect 562250 45922 562318 45978
rect 562374 45922 562442 45978
rect 562498 45922 562566 45978
rect 562622 45922 562718 45978
rect 562098 28350 562718 45922
rect 566188 53938 566244 53948
rect 562098 28294 562194 28350
rect 562250 28294 562318 28350
rect 562374 28294 562442 28350
rect 562498 28294 562566 28350
rect 562622 28294 562718 28350
rect 562098 28226 562718 28294
rect 562098 28170 562194 28226
rect 562250 28170 562318 28226
rect 562374 28170 562442 28226
rect 562498 28170 562566 28226
rect 562622 28170 562718 28226
rect 562098 28102 562718 28170
rect 562098 28046 562194 28102
rect 562250 28046 562318 28102
rect 562374 28046 562442 28102
rect 562498 28046 562566 28102
rect 562622 28046 562718 28102
rect 562098 27978 562718 28046
rect 562098 27922 562194 27978
rect 562250 27922 562318 27978
rect 562374 27922 562442 27978
rect 562498 27922 562566 27978
rect 562622 27922 562718 27978
rect 562098 10350 562718 27922
rect 562098 10294 562194 10350
rect 562250 10294 562318 10350
rect 562374 10294 562442 10350
rect 562498 10294 562566 10350
rect 562622 10294 562718 10350
rect 562098 10226 562718 10294
rect 562098 10170 562194 10226
rect 562250 10170 562318 10226
rect 562374 10170 562442 10226
rect 562498 10170 562566 10226
rect 562622 10170 562718 10226
rect 562098 10102 562718 10170
rect 562098 10046 562194 10102
rect 562250 10046 562318 10102
rect 562374 10046 562442 10102
rect 562498 10046 562566 10102
rect 562622 10046 562718 10102
rect 562098 9978 562718 10046
rect 562098 9922 562194 9978
rect 562250 9922 562318 9978
rect 562374 9922 562442 9978
rect 562498 9922 562566 9978
rect 562622 9922 562718 9978
rect 558378 4046 558474 4102
rect 558530 4046 558598 4102
rect 558654 4046 558722 4102
rect 558778 4046 558846 4102
rect 558902 4046 558998 4102
rect 558378 3978 558998 4046
rect 558378 3922 558474 3978
rect 558530 3922 558598 3978
rect 558654 3922 558722 3978
rect 558778 3922 558846 3978
rect 558902 3922 558998 3978
rect 557788 3178 557844 3188
rect 542556 1876 542612 1886
rect 542556 1378 542612 1820
rect 557788 1764 557844 3122
rect 557788 1698 557844 1708
rect 542556 1312 542612 1322
rect 531378 -1176 531474 -1120
rect 531530 -1176 531598 -1120
rect 531654 -1176 531722 -1120
rect 531778 -1176 531846 -1120
rect 531902 -1176 531998 -1120
rect 531378 -1244 531998 -1176
rect 531378 -1300 531474 -1244
rect 531530 -1300 531598 -1244
rect 531654 -1300 531722 -1244
rect 531778 -1300 531846 -1244
rect 531902 -1300 531998 -1244
rect 531378 -1368 531998 -1300
rect 531378 -1424 531474 -1368
rect 531530 -1424 531598 -1368
rect 531654 -1424 531722 -1368
rect 531778 -1424 531846 -1368
rect 531902 -1424 531998 -1368
rect 531378 -1492 531998 -1424
rect 531378 -1548 531474 -1492
rect 531530 -1548 531598 -1492
rect 531654 -1548 531722 -1492
rect 531778 -1548 531846 -1492
rect 531902 -1548 531998 -1492
rect 531378 -1644 531998 -1548
rect 558378 -160 558998 3922
rect 558378 -216 558474 -160
rect 558530 -216 558598 -160
rect 558654 -216 558722 -160
rect 558778 -216 558846 -160
rect 558902 -216 558998 -160
rect 558378 -284 558998 -216
rect 558378 -340 558474 -284
rect 558530 -340 558598 -284
rect 558654 -340 558722 -284
rect 558778 -340 558846 -284
rect 558902 -340 558998 -284
rect 558378 -408 558998 -340
rect 558378 -464 558474 -408
rect 558530 -464 558598 -408
rect 558654 -464 558722 -408
rect 558778 -464 558846 -408
rect 558902 -464 558998 -408
rect 558378 -532 558998 -464
rect 558378 -588 558474 -532
rect 558530 -588 558598 -532
rect 558654 -588 558722 -532
rect 558778 -588 558846 -532
rect 558902 -588 558998 -532
rect 558378 -1644 558998 -588
rect 562098 -1120 562718 9922
rect 564508 31978 564564 31988
rect 563500 6778 563556 6788
rect 563500 3444 563556 6722
rect 564508 4228 564564 31922
rect 564508 4162 564564 4172
rect 566188 4228 566244 53882
rect 572908 20188 572964 67202
rect 576268 65638 576324 65648
rect 575372 30324 575428 30334
rect 574588 25318 574644 25328
rect 572908 20132 573076 20188
rect 566188 4162 566244 4172
rect 573020 4228 573076 20132
rect 573020 4162 573076 4172
rect 574588 4228 574644 25262
rect 575372 7140 575428 30268
rect 575372 7074 575428 7084
rect 574588 4162 574644 4172
rect 576268 4228 576324 65582
rect 589098 58350 589718 75922
rect 589098 58294 589194 58350
rect 589250 58294 589318 58350
rect 589374 58294 589442 58350
rect 589498 58294 589566 58350
rect 589622 58294 589718 58350
rect 589098 58226 589718 58294
rect 589098 58170 589194 58226
rect 589250 58170 589318 58226
rect 589374 58170 589442 58226
rect 589498 58170 589566 58226
rect 589622 58170 589718 58226
rect 589098 58102 589718 58170
rect 589098 58046 589194 58102
rect 589250 58046 589318 58102
rect 589374 58046 589442 58102
rect 589498 58046 589566 58102
rect 589622 58046 589718 58102
rect 589098 57978 589718 58046
rect 589098 57922 589194 57978
rect 589250 57922 589318 57978
rect 589374 57922 589442 57978
rect 589498 57922 589566 57978
rect 589622 57922 589718 57978
rect 589098 40350 589718 57922
rect 592818 64350 593438 81922
rect 592818 64294 592914 64350
rect 592970 64294 593038 64350
rect 593094 64294 593162 64350
rect 593218 64294 593286 64350
rect 593342 64294 593438 64350
rect 592818 64226 593438 64294
rect 592818 64170 592914 64226
rect 592970 64170 593038 64226
rect 593094 64170 593162 64226
rect 593218 64170 593286 64226
rect 593342 64170 593438 64226
rect 592818 64102 593438 64170
rect 592818 64046 592914 64102
rect 592970 64046 593038 64102
rect 593094 64046 593162 64102
rect 593218 64046 593286 64102
rect 593342 64046 593438 64102
rect 592818 63978 593438 64046
rect 592818 63922 592914 63978
rect 592970 63922 593038 63978
rect 593094 63922 593162 63978
rect 593218 63922 593286 63978
rect 593342 63922 593438 63978
rect 589098 40294 589194 40350
rect 589250 40294 589318 40350
rect 589374 40294 589442 40350
rect 589498 40294 589566 40350
rect 589622 40294 589718 40350
rect 589098 40226 589718 40294
rect 589098 40170 589194 40226
rect 589250 40170 589318 40226
rect 589374 40170 589442 40226
rect 589498 40170 589566 40226
rect 589622 40170 589718 40226
rect 589098 40102 589718 40170
rect 589098 40046 589194 40102
rect 589250 40046 589318 40102
rect 589374 40046 589442 40102
rect 589498 40046 589566 40102
rect 589622 40046 589718 40102
rect 589098 39978 589718 40046
rect 589098 39922 589194 39978
rect 589250 39922 589318 39978
rect 589374 39922 589442 39978
rect 589498 39922 589566 39978
rect 589622 39922 589718 39978
rect 587132 32004 587188 32014
rect 587132 20580 587188 31948
rect 587132 20514 587188 20524
rect 589098 22350 589718 39922
rect 590492 46788 590548 46798
rect 590492 31108 590548 46732
rect 590492 31042 590548 31052
rect 592818 46350 593438 63922
rect 592818 46294 592914 46350
rect 592970 46294 593038 46350
rect 593094 46294 593162 46350
rect 593218 46294 593286 46350
rect 593342 46294 593438 46350
rect 592818 46226 593438 46294
rect 592818 46170 592914 46226
rect 592970 46170 593038 46226
rect 593094 46170 593162 46226
rect 593218 46170 593286 46226
rect 593342 46170 593438 46226
rect 592818 46102 593438 46170
rect 592818 46046 592914 46102
rect 592970 46046 593038 46102
rect 593094 46046 593162 46102
rect 593218 46046 593286 46102
rect 593342 46046 593438 46102
rect 592818 45978 593438 46046
rect 592818 45922 592914 45978
rect 592970 45922 593038 45978
rect 593094 45922 593162 45978
rect 593218 45922 593286 45978
rect 593342 45922 593438 45978
rect 589098 22294 589194 22350
rect 589250 22294 589318 22350
rect 589374 22294 589442 22350
rect 589498 22294 589566 22350
rect 589622 22294 589718 22350
rect 589098 22226 589718 22294
rect 589098 22170 589194 22226
rect 589250 22170 589318 22226
rect 589374 22170 589442 22226
rect 589498 22170 589566 22226
rect 589622 22170 589718 22226
rect 589098 22102 589718 22170
rect 589098 22046 589194 22102
rect 589250 22046 589318 22102
rect 589374 22046 589442 22102
rect 589498 22046 589566 22102
rect 589622 22046 589718 22102
rect 589098 21978 589718 22046
rect 589098 21922 589194 21978
rect 589250 21922 589318 21978
rect 589374 21922 589442 21978
rect 589498 21922 589566 21978
rect 589622 21922 589718 21978
rect 576268 4162 576324 4172
rect 589098 4350 589718 21922
rect 589098 4294 589194 4350
rect 589250 4294 589318 4350
rect 589374 4294 589442 4350
rect 589498 4294 589566 4350
rect 589622 4294 589718 4350
rect 589098 4226 589718 4294
rect 589098 4170 589194 4226
rect 589250 4170 589318 4226
rect 589374 4170 589442 4226
rect 589498 4170 589566 4226
rect 589622 4170 589718 4226
rect 563500 3378 563556 3388
rect 589098 4102 589718 4170
rect 589098 4046 589194 4102
rect 589250 4046 589318 4102
rect 589374 4046 589442 4102
rect 589498 4046 589566 4102
rect 589622 4046 589718 4102
rect 589098 3978 589718 4046
rect 589098 3922 589194 3978
rect 589250 3922 589318 3978
rect 589374 3922 589442 3978
rect 589498 3922 589566 3978
rect 589622 3922 589718 3978
rect 569548 1764 569604 1774
rect 569548 1558 569604 1708
rect 569548 1492 569604 1502
rect 562098 -1176 562194 -1120
rect 562250 -1176 562318 -1120
rect 562374 -1176 562442 -1120
rect 562498 -1176 562566 -1120
rect 562622 -1176 562718 -1120
rect 562098 -1244 562718 -1176
rect 562098 -1300 562194 -1244
rect 562250 -1300 562318 -1244
rect 562374 -1300 562442 -1244
rect 562498 -1300 562566 -1244
rect 562622 -1300 562718 -1244
rect 562098 -1368 562718 -1300
rect 562098 -1424 562194 -1368
rect 562250 -1424 562318 -1368
rect 562374 -1424 562442 -1368
rect 562498 -1424 562566 -1368
rect 562622 -1424 562718 -1368
rect 562098 -1492 562718 -1424
rect 562098 -1548 562194 -1492
rect 562250 -1548 562318 -1492
rect 562374 -1548 562442 -1492
rect 562498 -1548 562566 -1492
rect 562622 -1548 562718 -1492
rect 562098 -1644 562718 -1548
rect 589098 -160 589718 3922
rect 589098 -216 589194 -160
rect 589250 -216 589318 -160
rect 589374 -216 589442 -160
rect 589498 -216 589566 -160
rect 589622 -216 589718 -160
rect 589098 -284 589718 -216
rect 589098 -340 589194 -284
rect 589250 -340 589318 -284
rect 589374 -340 589442 -284
rect 589498 -340 589566 -284
rect 589622 -340 589718 -284
rect 589098 -408 589718 -340
rect 589098 -464 589194 -408
rect 589250 -464 589318 -408
rect 589374 -464 589442 -408
rect 589498 -464 589566 -408
rect 589622 -464 589718 -408
rect 589098 -532 589718 -464
rect 589098 -588 589194 -532
rect 589250 -588 589318 -532
rect 589374 -588 589442 -532
rect 589498 -588 589566 -532
rect 589622 -588 589718 -532
rect 589098 -1644 589718 -588
rect 592818 28350 593438 45922
rect 592818 28294 592914 28350
rect 592970 28294 593038 28350
rect 593094 28294 593162 28350
rect 593218 28294 593286 28350
rect 593342 28294 593438 28350
rect 592818 28226 593438 28294
rect 592818 28170 592914 28226
rect 592970 28170 593038 28226
rect 593094 28170 593162 28226
rect 593218 28170 593286 28226
rect 593342 28170 593438 28226
rect 592818 28102 593438 28170
rect 592818 28046 592914 28102
rect 592970 28046 593038 28102
rect 593094 28046 593162 28102
rect 593218 28046 593286 28102
rect 593342 28046 593438 28102
rect 592818 27978 593438 28046
rect 592818 27922 592914 27978
rect 592970 27922 593038 27978
rect 593094 27922 593162 27978
rect 593218 27922 593286 27978
rect 593342 27922 593438 27978
rect 592818 10350 593438 27922
rect 592818 10294 592914 10350
rect 592970 10294 593038 10350
rect 593094 10294 593162 10350
rect 593218 10294 593286 10350
rect 593342 10294 593438 10350
rect 592818 10226 593438 10294
rect 592818 10170 592914 10226
rect 592970 10170 593038 10226
rect 593094 10170 593162 10226
rect 593218 10170 593286 10226
rect 593342 10170 593438 10226
rect 592818 10102 593438 10170
rect 592818 10046 592914 10102
rect 592970 10046 593038 10102
rect 593094 10046 593162 10102
rect 593218 10046 593286 10102
rect 593342 10046 593438 10102
rect 592818 9978 593438 10046
rect 592818 9922 592914 9978
rect 592970 9922 593038 9978
rect 593094 9922 593162 9978
rect 593218 9922 593286 9978
rect 593342 9922 593438 9978
rect 592818 -1120 593438 9922
rect 596400 597212 597020 597308
rect 596400 597156 596496 597212
rect 596552 597156 596620 597212
rect 596676 597156 596744 597212
rect 596800 597156 596868 597212
rect 596924 597156 597020 597212
rect 596400 597088 597020 597156
rect 596400 597032 596496 597088
rect 596552 597032 596620 597088
rect 596676 597032 596744 597088
rect 596800 597032 596868 597088
rect 596924 597032 597020 597088
rect 596400 596964 597020 597032
rect 596400 596908 596496 596964
rect 596552 596908 596620 596964
rect 596676 596908 596744 596964
rect 596800 596908 596868 596964
rect 596924 596908 597020 596964
rect 596400 596840 597020 596908
rect 596400 596784 596496 596840
rect 596552 596784 596620 596840
rect 596676 596784 596744 596840
rect 596800 596784 596868 596840
rect 596924 596784 597020 596840
rect 596400 580350 597020 596784
rect 596400 580294 596496 580350
rect 596552 580294 596620 580350
rect 596676 580294 596744 580350
rect 596800 580294 596868 580350
rect 596924 580294 597020 580350
rect 596400 580226 597020 580294
rect 596400 580170 596496 580226
rect 596552 580170 596620 580226
rect 596676 580170 596744 580226
rect 596800 580170 596868 580226
rect 596924 580170 597020 580226
rect 596400 580102 597020 580170
rect 596400 580046 596496 580102
rect 596552 580046 596620 580102
rect 596676 580046 596744 580102
rect 596800 580046 596868 580102
rect 596924 580046 597020 580102
rect 596400 579978 597020 580046
rect 596400 579922 596496 579978
rect 596552 579922 596620 579978
rect 596676 579922 596744 579978
rect 596800 579922 596868 579978
rect 596924 579922 597020 579978
rect 596400 562350 597020 579922
rect 596400 562294 596496 562350
rect 596552 562294 596620 562350
rect 596676 562294 596744 562350
rect 596800 562294 596868 562350
rect 596924 562294 597020 562350
rect 596400 562226 597020 562294
rect 596400 562170 596496 562226
rect 596552 562170 596620 562226
rect 596676 562170 596744 562226
rect 596800 562170 596868 562226
rect 596924 562170 597020 562226
rect 596400 562102 597020 562170
rect 596400 562046 596496 562102
rect 596552 562046 596620 562102
rect 596676 562046 596744 562102
rect 596800 562046 596868 562102
rect 596924 562046 597020 562102
rect 596400 561978 597020 562046
rect 596400 561922 596496 561978
rect 596552 561922 596620 561978
rect 596676 561922 596744 561978
rect 596800 561922 596868 561978
rect 596924 561922 597020 561978
rect 596400 544350 597020 561922
rect 596400 544294 596496 544350
rect 596552 544294 596620 544350
rect 596676 544294 596744 544350
rect 596800 544294 596868 544350
rect 596924 544294 597020 544350
rect 596400 544226 597020 544294
rect 596400 544170 596496 544226
rect 596552 544170 596620 544226
rect 596676 544170 596744 544226
rect 596800 544170 596868 544226
rect 596924 544170 597020 544226
rect 596400 544102 597020 544170
rect 596400 544046 596496 544102
rect 596552 544046 596620 544102
rect 596676 544046 596744 544102
rect 596800 544046 596868 544102
rect 596924 544046 597020 544102
rect 596400 543978 597020 544046
rect 596400 543922 596496 543978
rect 596552 543922 596620 543978
rect 596676 543922 596744 543978
rect 596800 543922 596868 543978
rect 596924 543922 597020 543978
rect 596400 526350 597020 543922
rect 596400 526294 596496 526350
rect 596552 526294 596620 526350
rect 596676 526294 596744 526350
rect 596800 526294 596868 526350
rect 596924 526294 597020 526350
rect 596400 526226 597020 526294
rect 596400 526170 596496 526226
rect 596552 526170 596620 526226
rect 596676 526170 596744 526226
rect 596800 526170 596868 526226
rect 596924 526170 597020 526226
rect 596400 526102 597020 526170
rect 596400 526046 596496 526102
rect 596552 526046 596620 526102
rect 596676 526046 596744 526102
rect 596800 526046 596868 526102
rect 596924 526046 597020 526102
rect 596400 525978 597020 526046
rect 596400 525922 596496 525978
rect 596552 525922 596620 525978
rect 596676 525922 596744 525978
rect 596800 525922 596868 525978
rect 596924 525922 597020 525978
rect 596400 508350 597020 525922
rect 596400 508294 596496 508350
rect 596552 508294 596620 508350
rect 596676 508294 596744 508350
rect 596800 508294 596868 508350
rect 596924 508294 597020 508350
rect 596400 508226 597020 508294
rect 596400 508170 596496 508226
rect 596552 508170 596620 508226
rect 596676 508170 596744 508226
rect 596800 508170 596868 508226
rect 596924 508170 597020 508226
rect 596400 508102 597020 508170
rect 596400 508046 596496 508102
rect 596552 508046 596620 508102
rect 596676 508046 596744 508102
rect 596800 508046 596868 508102
rect 596924 508046 597020 508102
rect 596400 507978 597020 508046
rect 596400 507922 596496 507978
rect 596552 507922 596620 507978
rect 596676 507922 596744 507978
rect 596800 507922 596868 507978
rect 596924 507922 597020 507978
rect 596400 490350 597020 507922
rect 596400 490294 596496 490350
rect 596552 490294 596620 490350
rect 596676 490294 596744 490350
rect 596800 490294 596868 490350
rect 596924 490294 597020 490350
rect 596400 490226 597020 490294
rect 596400 490170 596496 490226
rect 596552 490170 596620 490226
rect 596676 490170 596744 490226
rect 596800 490170 596868 490226
rect 596924 490170 597020 490226
rect 596400 490102 597020 490170
rect 596400 490046 596496 490102
rect 596552 490046 596620 490102
rect 596676 490046 596744 490102
rect 596800 490046 596868 490102
rect 596924 490046 597020 490102
rect 596400 489978 597020 490046
rect 596400 489922 596496 489978
rect 596552 489922 596620 489978
rect 596676 489922 596744 489978
rect 596800 489922 596868 489978
rect 596924 489922 597020 489978
rect 596400 472350 597020 489922
rect 596400 472294 596496 472350
rect 596552 472294 596620 472350
rect 596676 472294 596744 472350
rect 596800 472294 596868 472350
rect 596924 472294 597020 472350
rect 596400 472226 597020 472294
rect 596400 472170 596496 472226
rect 596552 472170 596620 472226
rect 596676 472170 596744 472226
rect 596800 472170 596868 472226
rect 596924 472170 597020 472226
rect 596400 472102 597020 472170
rect 596400 472046 596496 472102
rect 596552 472046 596620 472102
rect 596676 472046 596744 472102
rect 596800 472046 596868 472102
rect 596924 472046 597020 472102
rect 596400 471978 597020 472046
rect 596400 471922 596496 471978
rect 596552 471922 596620 471978
rect 596676 471922 596744 471978
rect 596800 471922 596868 471978
rect 596924 471922 597020 471978
rect 596400 454350 597020 471922
rect 596400 454294 596496 454350
rect 596552 454294 596620 454350
rect 596676 454294 596744 454350
rect 596800 454294 596868 454350
rect 596924 454294 597020 454350
rect 596400 454226 597020 454294
rect 596400 454170 596496 454226
rect 596552 454170 596620 454226
rect 596676 454170 596744 454226
rect 596800 454170 596868 454226
rect 596924 454170 597020 454226
rect 596400 454102 597020 454170
rect 596400 454046 596496 454102
rect 596552 454046 596620 454102
rect 596676 454046 596744 454102
rect 596800 454046 596868 454102
rect 596924 454046 597020 454102
rect 596400 453978 597020 454046
rect 596400 453922 596496 453978
rect 596552 453922 596620 453978
rect 596676 453922 596744 453978
rect 596800 453922 596868 453978
rect 596924 453922 597020 453978
rect 596400 436350 597020 453922
rect 596400 436294 596496 436350
rect 596552 436294 596620 436350
rect 596676 436294 596744 436350
rect 596800 436294 596868 436350
rect 596924 436294 597020 436350
rect 596400 436226 597020 436294
rect 596400 436170 596496 436226
rect 596552 436170 596620 436226
rect 596676 436170 596744 436226
rect 596800 436170 596868 436226
rect 596924 436170 597020 436226
rect 596400 436102 597020 436170
rect 596400 436046 596496 436102
rect 596552 436046 596620 436102
rect 596676 436046 596744 436102
rect 596800 436046 596868 436102
rect 596924 436046 597020 436102
rect 596400 435978 597020 436046
rect 596400 435922 596496 435978
rect 596552 435922 596620 435978
rect 596676 435922 596744 435978
rect 596800 435922 596868 435978
rect 596924 435922 597020 435978
rect 596400 418350 597020 435922
rect 596400 418294 596496 418350
rect 596552 418294 596620 418350
rect 596676 418294 596744 418350
rect 596800 418294 596868 418350
rect 596924 418294 597020 418350
rect 596400 418226 597020 418294
rect 596400 418170 596496 418226
rect 596552 418170 596620 418226
rect 596676 418170 596744 418226
rect 596800 418170 596868 418226
rect 596924 418170 597020 418226
rect 596400 418102 597020 418170
rect 596400 418046 596496 418102
rect 596552 418046 596620 418102
rect 596676 418046 596744 418102
rect 596800 418046 596868 418102
rect 596924 418046 597020 418102
rect 596400 417978 597020 418046
rect 596400 417922 596496 417978
rect 596552 417922 596620 417978
rect 596676 417922 596744 417978
rect 596800 417922 596868 417978
rect 596924 417922 597020 417978
rect 596400 400350 597020 417922
rect 596400 400294 596496 400350
rect 596552 400294 596620 400350
rect 596676 400294 596744 400350
rect 596800 400294 596868 400350
rect 596924 400294 597020 400350
rect 596400 400226 597020 400294
rect 596400 400170 596496 400226
rect 596552 400170 596620 400226
rect 596676 400170 596744 400226
rect 596800 400170 596868 400226
rect 596924 400170 597020 400226
rect 596400 400102 597020 400170
rect 596400 400046 596496 400102
rect 596552 400046 596620 400102
rect 596676 400046 596744 400102
rect 596800 400046 596868 400102
rect 596924 400046 597020 400102
rect 596400 399978 597020 400046
rect 596400 399922 596496 399978
rect 596552 399922 596620 399978
rect 596676 399922 596744 399978
rect 596800 399922 596868 399978
rect 596924 399922 597020 399978
rect 596400 382350 597020 399922
rect 596400 382294 596496 382350
rect 596552 382294 596620 382350
rect 596676 382294 596744 382350
rect 596800 382294 596868 382350
rect 596924 382294 597020 382350
rect 596400 382226 597020 382294
rect 596400 382170 596496 382226
rect 596552 382170 596620 382226
rect 596676 382170 596744 382226
rect 596800 382170 596868 382226
rect 596924 382170 597020 382226
rect 596400 382102 597020 382170
rect 596400 382046 596496 382102
rect 596552 382046 596620 382102
rect 596676 382046 596744 382102
rect 596800 382046 596868 382102
rect 596924 382046 597020 382102
rect 596400 381978 597020 382046
rect 596400 381922 596496 381978
rect 596552 381922 596620 381978
rect 596676 381922 596744 381978
rect 596800 381922 596868 381978
rect 596924 381922 597020 381978
rect 596400 364350 597020 381922
rect 596400 364294 596496 364350
rect 596552 364294 596620 364350
rect 596676 364294 596744 364350
rect 596800 364294 596868 364350
rect 596924 364294 597020 364350
rect 596400 364226 597020 364294
rect 596400 364170 596496 364226
rect 596552 364170 596620 364226
rect 596676 364170 596744 364226
rect 596800 364170 596868 364226
rect 596924 364170 597020 364226
rect 596400 364102 597020 364170
rect 596400 364046 596496 364102
rect 596552 364046 596620 364102
rect 596676 364046 596744 364102
rect 596800 364046 596868 364102
rect 596924 364046 597020 364102
rect 596400 363978 597020 364046
rect 596400 363922 596496 363978
rect 596552 363922 596620 363978
rect 596676 363922 596744 363978
rect 596800 363922 596868 363978
rect 596924 363922 597020 363978
rect 596400 346350 597020 363922
rect 596400 346294 596496 346350
rect 596552 346294 596620 346350
rect 596676 346294 596744 346350
rect 596800 346294 596868 346350
rect 596924 346294 597020 346350
rect 596400 346226 597020 346294
rect 596400 346170 596496 346226
rect 596552 346170 596620 346226
rect 596676 346170 596744 346226
rect 596800 346170 596868 346226
rect 596924 346170 597020 346226
rect 596400 346102 597020 346170
rect 596400 346046 596496 346102
rect 596552 346046 596620 346102
rect 596676 346046 596744 346102
rect 596800 346046 596868 346102
rect 596924 346046 597020 346102
rect 596400 345978 597020 346046
rect 596400 345922 596496 345978
rect 596552 345922 596620 345978
rect 596676 345922 596744 345978
rect 596800 345922 596868 345978
rect 596924 345922 597020 345978
rect 596400 328350 597020 345922
rect 596400 328294 596496 328350
rect 596552 328294 596620 328350
rect 596676 328294 596744 328350
rect 596800 328294 596868 328350
rect 596924 328294 597020 328350
rect 596400 328226 597020 328294
rect 596400 328170 596496 328226
rect 596552 328170 596620 328226
rect 596676 328170 596744 328226
rect 596800 328170 596868 328226
rect 596924 328170 597020 328226
rect 596400 328102 597020 328170
rect 596400 328046 596496 328102
rect 596552 328046 596620 328102
rect 596676 328046 596744 328102
rect 596800 328046 596868 328102
rect 596924 328046 597020 328102
rect 596400 327978 597020 328046
rect 596400 327922 596496 327978
rect 596552 327922 596620 327978
rect 596676 327922 596744 327978
rect 596800 327922 596868 327978
rect 596924 327922 597020 327978
rect 596400 310350 597020 327922
rect 596400 310294 596496 310350
rect 596552 310294 596620 310350
rect 596676 310294 596744 310350
rect 596800 310294 596868 310350
rect 596924 310294 597020 310350
rect 596400 310226 597020 310294
rect 596400 310170 596496 310226
rect 596552 310170 596620 310226
rect 596676 310170 596744 310226
rect 596800 310170 596868 310226
rect 596924 310170 597020 310226
rect 596400 310102 597020 310170
rect 596400 310046 596496 310102
rect 596552 310046 596620 310102
rect 596676 310046 596744 310102
rect 596800 310046 596868 310102
rect 596924 310046 597020 310102
rect 596400 309978 597020 310046
rect 596400 309922 596496 309978
rect 596552 309922 596620 309978
rect 596676 309922 596744 309978
rect 596800 309922 596868 309978
rect 596924 309922 597020 309978
rect 596400 292350 597020 309922
rect 596400 292294 596496 292350
rect 596552 292294 596620 292350
rect 596676 292294 596744 292350
rect 596800 292294 596868 292350
rect 596924 292294 597020 292350
rect 596400 292226 597020 292294
rect 596400 292170 596496 292226
rect 596552 292170 596620 292226
rect 596676 292170 596744 292226
rect 596800 292170 596868 292226
rect 596924 292170 597020 292226
rect 596400 292102 597020 292170
rect 596400 292046 596496 292102
rect 596552 292046 596620 292102
rect 596676 292046 596744 292102
rect 596800 292046 596868 292102
rect 596924 292046 597020 292102
rect 596400 291978 597020 292046
rect 596400 291922 596496 291978
rect 596552 291922 596620 291978
rect 596676 291922 596744 291978
rect 596800 291922 596868 291978
rect 596924 291922 597020 291978
rect 596400 274350 597020 291922
rect 596400 274294 596496 274350
rect 596552 274294 596620 274350
rect 596676 274294 596744 274350
rect 596800 274294 596868 274350
rect 596924 274294 597020 274350
rect 596400 274226 597020 274294
rect 596400 274170 596496 274226
rect 596552 274170 596620 274226
rect 596676 274170 596744 274226
rect 596800 274170 596868 274226
rect 596924 274170 597020 274226
rect 596400 274102 597020 274170
rect 596400 274046 596496 274102
rect 596552 274046 596620 274102
rect 596676 274046 596744 274102
rect 596800 274046 596868 274102
rect 596924 274046 597020 274102
rect 596400 273978 597020 274046
rect 596400 273922 596496 273978
rect 596552 273922 596620 273978
rect 596676 273922 596744 273978
rect 596800 273922 596868 273978
rect 596924 273922 597020 273978
rect 596400 256350 597020 273922
rect 596400 256294 596496 256350
rect 596552 256294 596620 256350
rect 596676 256294 596744 256350
rect 596800 256294 596868 256350
rect 596924 256294 597020 256350
rect 596400 256226 597020 256294
rect 596400 256170 596496 256226
rect 596552 256170 596620 256226
rect 596676 256170 596744 256226
rect 596800 256170 596868 256226
rect 596924 256170 597020 256226
rect 596400 256102 597020 256170
rect 596400 256046 596496 256102
rect 596552 256046 596620 256102
rect 596676 256046 596744 256102
rect 596800 256046 596868 256102
rect 596924 256046 597020 256102
rect 596400 255978 597020 256046
rect 596400 255922 596496 255978
rect 596552 255922 596620 255978
rect 596676 255922 596744 255978
rect 596800 255922 596868 255978
rect 596924 255922 597020 255978
rect 596400 238350 597020 255922
rect 596400 238294 596496 238350
rect 596552 238294 596620 238350
rect 596676 238294 596744 238350
rect 596800 238294 596868 238350
rect 596924 238294 597020 238350
rect 596400 238226 597020 238294
rect 596400 238170 596496 238226
rect 596552 238170 596620 238226
rect 596676 238170 596744 238226
rect 596800 238170 596868 238226
rect 596924 238170 597020 238226
rect 596400 238102 597020 238170
rect 596400 238046 596496 238102
rect 596552 238046 596620 238102
rect 596676 238046 596744 238102
rect 596800 238046 596868 238102
rect 596924 238046 597020 238102
rect 596400 237978 597020 238046
rect 596400 237922 596496 237978
rect 596552 237922 596620 237978
rect 596676 237922 596744 237978
rect 596800 237922 596868 237978
rect 596924 237922 597020 237978
rect 596400 220350 597020 237922
rect 596400 220294 596496 220350
rect 596552 220294 596620 220350
rect 596676 220294 596744 220350
rect 596800 220294 596868 220350
rect 596924 220294 597020 220350
rect 596400 220226 597020 220294
rect 596400 220170 596496 220226
rect 596552 220170 596620 220226
rect 596676 220170 596744 220226
rect 596800 220170 596868 220226
rect 596924 220170 597020 220226
rect 596400 220102 597020 220170
rect 596400 220046 596496 220102
rect 596552 220046 596620 220102
rect 596676 220046 596744 220102
rect 596800 220046 596868 220102
rect 596924 220046 597020 220102
rect 596400 219978 597020 220046
rect 596400 219922 596496 219978
rect 596552 219922 596620 219978
rect 596676 219922 596744 219978
rect 596800 219922 596868 219978
rect 596924 219922 597020 219978
rect 596400 202350 597020 219922
rect 596400 202294 596496 202350
rect 596552 202294 596620 202350
rect 596676 202294 596744 202350
rect 596800 202294 596868 202350
rect 596924 202294 597020 202350
rect 596400 202226 597020 202294
rect 596400 202170 596496 202226
rect 596552 202170 596620 202226
rect 596676 202170 596744 202226
rect 596800 202170 596868 202226
rect 596924 202170 597020 202226
rect 596400 202102 597020 202170
rect 596400 202046 596496 202102
rect 596552 202046 596620 202102
rect 596676 202046 596744 202102
rect 596800 202046 596868 202102
rect 596924 202046 597020 202102
rect 596400 201978 597020 202046
rect 596400 201922 596496 201978
rect 596552 201922 596620 201978
rect 596676 201922 596744 201978
rect 596800 201922 596868 201978
rect 596924 201922 597020 201978
rect 596400 184350 597020 201922
rect 596400 184294 596496 184350
rect 596552 184294 596620 184350
rect 596676 184294 596744 184350
rect 596800 184294 596868 184350
rect 596924 184294 597020 184350
rect 596400 184226 597020 184294
rect 596400 184170 596496 184226
rect 596552 184170 596620 184226
rect 596676 184170 596744 184226
rect 596800 184170 596868 184226
rect 596924 184170 597020 184226
rect 596400 184102 597020 184170
rect 596400 184046 596496 184102
rect 596552 184046 596620 184102
rect 596676 184046 596744 184102
rect 596800 184046 596868 184102
rect 596924 184046 597020 184102
rect 596400 183978 597020 184046
rect 596400 183922 596496 183978
rect 596552 183922 596620 183978
rect 596676 183922 596744 183978
rect 596800 183922 596868 183978
rect 596924 183922 597020 183978
rect 596400 166350 597020 183922
rect 596400 166294 596496 166350
rect 596552 166294 596620 166350
rect 596676 166294 596744 166350
rect 596800 166294 596868 166350
rect 596924 166294 597020 166350
rect 596400 166226 597020 166294
rect 596400 166170 596496 166226
rect 596552 166170 596620 166226
rect 596676 166170 596744 166226
rect 596800 166170 596868 166226
rect 596924 166170 597020 166226
rect 596400 166102 597020 166170
rect 596400 166046 596496 166102
rect 596552 166046 596620 166102
rect 596676 166046 596744 166102
rect 596800 166046 596868 166102
rect 596924 166046 597020 166102
rect 596400 165978 597020 166046
rect 596400 165922 596496 165978
rect 596552 165922 596620 165978
rect 596676 165922 596744 165978
rect 596800 165922 596868 165978
rect 596924 165922 597020 165978
rect 596400 148350 597020 165922
rect 596400 148294 596496 148350
rect 596552 148294 596620 148350
rect 596676 148294 596744 148350
rect 596800 148294 596868 148350
rect 596924 148294 597020 148350
rect 596400 148226 597020 148294
rect 596400 148170 596496 148226
rect 596552 148170 596620 148226
rect 596676 148170 596744 148226
rect 596800 148170 596868 148226
rect 596924 148170 597020 148226
rect 596400 148102 597020 148170
rect 596400 148046 596496 148102
rect 596552 148046 596620 148102
rect 596676 148046 596744 148102
rect 596800 148046 596868 148102
rect 596924 148046 597020 148102
rect 596400 147978 597020 148046
rect 596400 147922 596496 147978
rect 596552 147922 596620 147978
rect 596676 147922 596744 147978
rect 596800 147922 596868 147978
rect 596924 147922 597020 147978
rect 596400 130350 597020 147922
rect 596400 130294 596496 130350
rect 596552 130294 596620 130350
rect 596676 130294 596744 130350
rect 596800 130294 596868 130350
rect 596924 130294 597020 130350
rect 596400 130226 597020 130294
rect 596400 130170 596496 130226
rect 596552 130170 596620 130226
rect 596676 130170 596744 130226
rect 596800 130170 596868 130226
rect 596924 130170 597020 130226
rect 596400 130102 597020 130170
rect 596400 130046 596496 130102
rect 596552 130046 596620 130102
rect 596676 130046 596744 130102
rect 596800 130046 596868 130102
rect 596924 130046 597020 130102
rect 596400 129978 597020 130046
rect 596400 129922 596496 129978
rect 596552 129922 596620 129978
rect 596676 129922 596744 129978
rect 596800 129922 596868 129978
rect 596924 129922 597020 129978
rect 596400 112350 597020 129922
rect 596400 112294 596496 112350
rect 596552 112294 596620 112350
rect 596676 112294 596744 112350
rect 596800 112294 596868 112350
rect 596924 112294 597020 112350
rect 596400 112226 597020 112294
rect 596400 112170 596496 112226
rect 596552 112170 596620 112226
rect 596676 112170 596744 112226
rect 596800 112170 596868 112226
rect 596924 112170 597020 112226
rect 596400 112102 597020 112170
rect 596400 112046 596496 112102
rect 596552 112046 596620 112102
rect 596676 112046 596744 112102
rect 596800 112046 596868 112102
rect 596924 112046 597020 112102
rect 596400 111978 597020 112046
rect 596400 111922 596496 111978
rect 596552 111922 596620 111978
rect 596676 111922 596744 111978
rect 596800 111922 596868 111978
rect 596924 111922 597020 111978
rect 596400 94350 597020 111922
rect 596400 94294 596496 94350
rect 596552 94294 596620 94350
rect 596676 94294 596744 94350
rect 596800 94294 596868 94350
rect 596924 94294 597020 94350
rect 596400 94226 597020 94294
rect 596400 94170 596496 94226
rect 596552 94170 596620 94226
rect 596676 94170 596744 94226
rect 596800 94170 596868 94226
rect 596924 94170 597020 94226
rect 596400 94102 597020 94170
rect 596400 94046 596496 94102
rect 596552 94046 596620 94102
rect 596676 94046 596744 94102
rect 596800 94046 596868 94102
rect 596924 94046 597020 94102
rect 596400 93978 597020 94046
rect 596400 93922 596496 93978
rect 596552 93922 596620 93978
rect 596676 93922 596744 93978
rect 596800 93922 596868 93978
rect 596924 93922 597020 93978
rect 596400 76350 597020 93922
rect 596400 76294 596496 76350
rect 596552 76294 596620 76350
rect 596676 76294 596744 76350
rect 596800 76294 596868 76350
rect 596924 76294 597020 76350
rect 596400 76226 597020 76294
rect 596400 76170 596496 76226
rect 596552 76170 596620 76226
rect 596676 76170 596744 76226
rect 596800 76170 596868 76226
rect 596924 76170 597020 76226
rect 596400 76102 597020 76170
rect 596400 76046 596496 76102
rect 596552 76046 596620 76102
rect 596676 76046 596744 76102
rect 596800 76046 596868 76102
rect 596924 76046 597020 76102
rect 596400 75978 597020 76046
rect 596400 75922 596496 75978
rect 596552 75922 596620 75978
rect 596676 75922 596744 75978
rect 596800 75922 596868 75978
rect 596924 75922 597020 75978
rect 596400 58350 597020 75922
rect 596400 58294 596496 58350
rect 596552 58294 596620 58350
rect 596676 58294 596744 58350
rect 596800 58294 596868 58350
rect 596924 58294 597020 58350
rect 596400 58226 597020 58294
rect 596400 58170 596496 58226
rect 596552 58170 596620 58226
rect 596676 58170 596744 58226
rect 596800 58170 596868 58226
rect 596924 58170 597020 58226
rect 596400 58102 597020 58170
rect 596400 58046 596496 58102
rect 596552 58046 596620 58102
rect 596676 58046 596744 58102
rect 596800 58046 596868 58102
rect 596924 58046 597020 58102
rect 596400 57978 597020 58046
rect 596400 57922 596496 57978
rect 596552 57922 596620 57978
rect 596676 57922 596744 57978
rect 596800 57922 596868 57978
rect 596924 57922 597020 57978
rect 596400 40350 597020 57922
rect 596400 40294 596496 40350
rect 596552 40294 596620 40350
rect 596676 40294 596744 40350
rect 596800 40294 596868 40350
rect 596924 40294 597020 40350
rect 596400 40226 597020 40294
rect 596400 40170 596496 40226
rect 596552 40170 596620 40226
rect 596676 40170 596744 40226
rect 596800 40170 596868 40226
rect 596924 40170 597020 40226
rect 596400 40102 597020 40170
rect 596400 40046 596496 40102
rect 596552 40046 596620 40102
rect 596676 40046 596744 40102
rect 596800 40046 596868 40102
rect 596924 40046 597020 40102
rect 596400 39978 597020 40046
rect 596400 39922 596496 39978
rect 596552 39922 596620 39978
rect 596676 39922 596744 39978
rect 596800 39922 596868 39978
rect 596924 39922 597020 39978
rect 596400 22350 597020 39922
rect 596400 22294 596496 22350
rect 596552 22294 596620 22350
rect 596676 22294 596744 22350
rect 596800 22294 596868 22350
rect 596924 22294 597020 22350
rect 596400 22226 597020 22294
rect 596400 22170 596496 22226
rect 596552 22170 596620 22226
rect 596676 22170 596744 22226
rect 596800 22170 596868 22226
rect 596924 22170 597020 22226
rect 596400 22102 597020 22170
rect 596400 22046 596496 22102
rect 596552 22046 596620 22102
rect 596676 22046 596744 22102
rect 596800 22046 596868 22102
rect 596924 22046 597020 22102
rect 596400 21978 597020 22046
rect 596400 21922 596496 21978
rect 596552 21922 596620 21978
rect 596676 21922 596744 21978
rect 596800 21922 596868 21978
rect 596924 21922 597020 21978
rect 596400 4350 597020 21922
rect 596400 4294 596496 4350
rect 596552 4294 596620 4350
rect 596676 4294 596744 4350
rect 596800 4294 596868 4350
rect 596924 4294 597020 4350
rect 596400 4226 597020 4294
rect 596400 4170 596496 4226
rect 596552 4170 596620 4226
rect 596676 4170 596744 4226
rect 596800 4170 596868 4226
rect 596924 4170 597020 4226
rect 596400 4102 597020 4170
rect 596400 4046 596496 4102
rect 596552 4046 596620 4102
rect 596676 4046 596744 4102
rect 596800 4046 596868 4102
rect 596924 4046 597020 4102
rect 596400 3978 597020 4046
rect 596400 3922 596496 3978
rect 596552 3922 596620 3978
rect 596676 3922 596744 3978
rect 596800 3922 596868 3978
rect 596924 3922 597020 3978
rect 596400 -160 597020 3922
rect 596400 -216 596496 -160
rect 596552 -216 596620 -160
rect 596676 -216 596744 -160
rect 596800 -216 596868 -160
rect 596924 -216 597020 -160
rect 596400 -284 597020 -216
rect 596400 -340 596496 -284
rect 596552 -340 596620 -284
rect 596676 -340 596744 -284
rect 596800 -340 596868 -284
rect 596924 -340 597020 -284
rect 596400 -408 597020 -340
rect 596400 -464 596496 -408
rect 596552 -464 596620 -408
rect 596676 -464 596744 -408
rect 596800 -464 596868 -408
rect 596924 -464 597020 -408
rect 596400 -532 597020 -464
rect 596400 -588 596496 -532
rect 596552 -588 596620 -532
rect 596676 -588 596744 -532
rect 596800 -588 596868 -532
rect 596924 -588 597020 -532
rect 596400 -684 597020 -588
rect 597360 586350 597980 597744
rect 597360 586294 597456 586350
rect 597512 586294 597580 586350
rect 597636 586294 597704 586350
rect 597760 586294 597828 586350
rect 597884 586294 597980 586350
rect 597360 586226 597980 586294
rect 597360 586170 597456 586226
rect 597512 586170 597580 586226
rect 597636 586170 597704 586226
rect 597760 586170 597828 586226
rect 597884 586170 597980 586226
rect 597360 586102 597980 586170
rect 597360 586046 597456 586102
rect 597512 586046 597580 586102
rect 597636 586046 597704 586102
rect 597760 586046 597828 586102
rect 597884 586046 597980 586102
rect 597360 585978 597980 586046
rect 597360 585922 597456 585978
rect 597512 585922 597580 585978
rect 597636 585922 597704 585978
rect 597760 585922 597828 585978
rect 597884 585922 597980 585978
rect 597360 568350 597980 585922
rect 597360 568294 597456 568350
rect 597512 568294 597580 568350
rect 597636 568294 597704 568350
rect 597760 568294 597828 568350
rect 597884 568294 597980 568350
rect 597360 568226 597980 568294
rect 597360 568170 597456 568226
rect 597512 568170 597580 568226
rect 597636 568170 597704 568226
rect 597760 568170 597828 568226
rect 597884 568170 597980 568226
rect 597360 568102 597980 568170
rect 597360 568046 597456 568102
rect 597512 568046 597580 568102
rect 597636 568046 597704 568102
rect 597760 568046 597828 568102
rect 597884 568046 597980 568102
rect 597360 567978 597980 568046
rect 597360 567922 597456 567978
rect 597512 567922 597580 567978
rect 597636 567922 597704 567978
rect 597760 567922 597828 567978
rect 597884 567922 597980 567978
rect 597360 550350 597980 567922
rect 597360 550294 597456 550350
rect 597512 550294 597580 550350
rect 597636 550294 597704 550350
rect 597760 550294 597828 550350
rect 597884 550294 597980 550350
rect 597360 550226 597980 550294
rect 597360 550170 597456 550226
rect 597512 550170 597580 550226
rect 597636 550170 597704 550226
rect 597760 550170 597828 550226
rect 597884 550170 597980 550226
rect 597360 550102 597980 550170
rect 597360 550046 597456 550102
rect 597512 550046 597580 550102
rect 597636 550046 597704 550102
rect 597760 550046 597828 550102
rect 597884 550046 597980 550102
rect 597360 549978 597980 550046
rect 597360 549922 597456 549978
rect 597512 549922 597580 549978
rect 597636 549922 597704 549978
rect 597760 549922 597828 549978
rect 597884 549922 597980 549978
rect 597360 532350 597980 549922
rect 597360 532294 597456 532350
rect 597512 532294 597580 532350
rect 597636 532294 597704 532350
rect 597760 532294 597828 532350
rect 597884 532294 597980 532350
rect 597360 532226 597980 532294
rect 597360 532170 597456 532226
rect 597512 532170 597580 532226
rect 597636 532170 597704 532226
rect 597760 532170 597828 532226
rect 597884 532170 597980 532226
rect 597360 532102 597980 532170
rect 597360 532046 597456 532102
rect 597512 532046 597580 532102
rect 597636 532046 597704 532102
rect 597760 532046 597828 532102
rect 597884 532046 597980 532102
rect 597360 531978 597980 532046
rect 597360 531922 597456 531978
rect 597512 531922 597580 531978
rect 597636 531922 597704 531978
rect 597760 531922 597828 531978
rect 597884 531922 597980 531978
rect 597360 514350 597980 531922
rect 597360 514294 597456 514350
rect 597512 514294 597580 514350
rect 597636 514294 597704 514350
rect 597760 514294 597828 514350
rect 597884 514294 597980 514350
rect 597360 514226 597980 514294
rect 597360 514170 597456 514226
rect 597512 514170 597580 514226
rect 597636 514170 597704 514226
rect 597760 514170 597828 514226
rect 597884 514170 597980 514226
rect 597360 514102 597980 514170
rect 597360 514046 597456 514102
rect 597512 514046 597580 514102
rect 597636 514046 597704 514102
rect 597760 514046 597828 514102
rect 597884 514046 597980 514102
rect 597360 513978 597980 514046
rect 597360 513922 597456 513978
rect 597512 513922 597580 513978
rect 597636 513922 597704 513978
rect 597760 513922 597828 513978
rect 597884 513922 597980 513978
rect 597360 496350 597980 513922
rect 597360 496294 597456 496350
rect 597512 496294 597580 496350
rect 597636 496294 597704 496350
rect 597760 496294 597828 496350
rect 597884 496294 597980 496350
rect 597360 496226 597980 496294
rect 597360 496170 597456 496226
rect 597512 496170 597580 496226
rect 597636 496170 597704 496226
rect 597760 496170 597828 496226
rect 597884 496170 597980 496226
rect 597360 496102 597980 496170
rect 597360 496046 597456 496102
rect 597512 496046 597580 496102
rect 597636 496046 597704 496102
rect 597760 496046 597828 496102
rect 597884 496046 597980 496102
rect 597360 495978 597980 496046
rect 597360 495922 597456 495978
rect 597512 495922 597580 495978
rect 597636 495922 597704 495978
rect 597760 495922 597828 495978
rect 597884 495922 597980 495978
rect 597360 478350 597980 495922
rect 597360 478294 597456 478350
rect 597512 478294 597580 478350
rect 597636 478294 597704 478350
rect 597760 478294 597828 478350
rect 597884 478294 597980 478350
rect 597360 478226 597980 478294
rect 597360 478170 597456 478226
rect 597512 478170 597580 478226
rect 597636 478170 597704 478226
rect 597760 478170 597828 478226
rect 597884 478170 597980 478226
rect 597360 478102 597980 478170
rect 597360 478046 597456 478102
rect 597512 478046 597580 478102
rect 597636 478046 597704 478102
rect 597760 478046 597828 478102
rect 597884 478046 597980 478102
rect 597360 477978 597980 478046
rect 597360 477922 597456 477978
rect 597512 477922 597580 477978
rect 597636 477922 597704 477978
rect 597760 477922 597828 477978
rect 597884 477922 597980 477978
rect 597360 460350 597980 477922
rect 597360 460294 597456 460350
rect 597512 460294 597580 460350
rect 597636 460294 597704 460350
rect 597760 460294 597828 460350
rect 597884 460294 597980 460350
rect 597360 460226 597980 460294
rect 597360 460170 597456 460226
rect 597512 460170 597580 460226
rect 597636 460170 597704 460226
rect 597760 460170 597828 460226
rect 597884 460170 597980 460226
rect 597360 460102 597980 460170
rect 597360 460046 597456 460102
rect 597512 460046 597580 460102
rect 597636 460046 597704 460102
rect 597760 460046 597828 460102
rect 597884 460046 597980 460102
rect 597360 459978 597980 460046
rect 597360 459922 597456 459978
rect 597512 459922 597580 459978
rect 597636 459922 597704 459978
rect 597760 459922 597828 459978
rect 597884 459922 597980 459978
rect 597360 442350 597980 459922
rect 597360 442294 597456 442350
rect 597512 442294 597580 442350
rect 597636 442294 597704 442350
rect 597760 442294 597828 442350
rect 597884 442294 597980 442350
rect 597360 442226 597980 442294
rect 597360 442170 597456 442226
rect 597512 442170 597580 442226
rect 597636 442170 597704 442226
rect 597760 442170 597828 442226
rect 597884 442170 597980 442226
rect 597360 442102 597980 442170
rect 597360 442046 597456 442102
rect 597512 442046 597580 442102
rect 597636 442046 597704 442102
rect 597760 442046 597828 442102
rect 597884 442046 597980 442102
rect 597360 441978 597980 442046
rect 597360 441922 597456 441978
rect 597512 441922 597580 441978
rect 597636 441922 597704 441978
rect 597760 441922 597828 441978
rect 597884 441922 597980 441978
rect 597360 424350 597980 441922
rect 597360 424294 597456 424350
rect 597512 424294 597580 424350
rect 597636 424294 597704 424350
rect 597760 424294 597828 424350
rect 597884 424294 597980 424350
rect 597360 424226 597980 424294
rect 597360 424170 597456 424226
rect 597512 424170 597580 424226
rect 597636 424170 597704 424226
rect 597760 424170 597828 424226
rect 597884 424170 597980 424226
rect 597360 424102 597980 424170
rect 597360 424046 597456 424102
rect 597512 424046 597580 424102
rect 597636 424046 597704 424102
rect 597760 424046 597828 424102
rect 597884 424046 597980 424102
rect 597360 423978 597980 424046
rect 597360 423922 597456 423978
rect 597512 423922 597580 423978
rect 597636 423922 597704 423978
rect 597760 423922 597828 423978
rect 597884 423922 597980 423978
rect 597360 406350 597980 423922
rect 597360 406294 597456 406350
rect 597512 406294 597580 406350
rect 597636 406294 597704 406350
rect 597760 406294 597828 406350
rect 597884 406294 597980 406350
rect 597360 406226 597980 406294
rect 597360 406170 597456 406226
rect 597512 406170 597580 406226
rect 597636 406170 597704 406226
rect 597760 406170 597828 406226
rect 597884 406170 597980 406226
rect 597360 406102 597980 406170
rect 597360 406046 597456 406102
rect 597512 406046 597580 406102
rect 597636 406046 597704 406102
rect 597760 406046 597828 406102
rect 597884 406046 597980 406102
rect 597360 405978 597980 406046
rect 597360 405922 597456 405978
rect 597512 405922 597580 405978
rect 597636 405922 597704 405978
rect 597760 405922 597828 405978
rect 597884 405922 597980 405978
rect 597360 388350 597980 405922
rect 597360 388294 597456 388350
rect 597512 388294 597580 388350
rect 597636 388294 597704 388350
rect 597760 388294 597828 388350
rect 597884 388294 597980 388350
rect 597360 388226 597980 388294
rect 597360 388170 597456 388226
rect 597512 388170 597580 388226
rect 597636 388170 597704 388226
rect 597760 388170 597828 388226
rect 597884 388170 597980 388226
rect 597360 388102 597980 388170
rect 597360 388046 597456 388102
rect 597512 388046 597580 388102
rect 597636 388046 597704 388102
rect 597760 388046 597828 388102
rect 597884 388046 597980 388102
rect 597360 387978 597980 388046
rect 597360 387922 597456 387978
rect 597512 387922 597580 387978
rect 597636 387922 597704 387978
rect 597760 387922 597828 387978
rect 597884 387922 597980 387978
rect 597360 370350 597980 387922
rect 597360 370294 597456 370350
rect 597512 370294 597580 370350
rect 597636 370294 597704 370350
rect 597760 370294 597828 370350
rect 597884 370294 597980 370350
rect 597360 370226 597980 370294
rect 597360 370170 597456 370226
rect 597512 370170 597580 370226
rect 597636 370170 597704 370226
rect 597760 370170 597828 370226
rect 597884 370170 597980 370226
rect 597360 370102 597980 370170
rect 597360 370046 597456 370102
rect 597512 370046 597580 370102
rect 597636 370046 597704 370102
rect 597760 370046 597828 370102
rect 597884 370046 597980 370102
rect 597360 369978 597980 370046
rect 597360 369922 597456 369978
rect 597512 369922 597580 369978
rect 597636 369922 597704 369978
rect 597760 369922 597828 369978
rect 597884 369922 597980 369978
rect 597360 352350 597980 369922
rect 597360 352294 597456 352350
rect 597512 352294 597580 352350
rect 597636 352294 597704 352350
rect 597760 352294 597828 352350
rect 597884 352294 597980 352350
rect 597360 352226 597980 352294
rect 597360 352170 597456 352226
rect 597512 352170 597580 352226
rect 597636 352170 597704 352226
rect 597760 352170 597828 352226
rect 597884 352170 597980 352226
rect 597360 352102 597980 352170
rect 597360 352046 597456 352102
rect 597512 352046 597580 352102
rect 597636 352046 597704 352102
rect 597760 352046 597828 352102
rect 597884 352046 597980 352102
rect 597360 351978 597980 352046
rect 597360 351922 597456 351978
rect 597512 351922 597580 351978
rect 597636 351922 597704 351978
rect 597760 351922 597828 351978
rect 597884 351922 597980 351978
rect 597360 334350 597980 351922
rect 597360 334294 597456 334350
rect 597512 334294 597580 334350
rect 597636 334294 597704 334350
rect 597760 334294 597828 334350
rect 597884 334294 597980 334350
rect 597360 334226 597980 334294
rect 597360 334170 597456 334226
rect 597512 334170 597580 334226
rect 597636 334170 597704 334226
rect 597760 334170 597828 334226
rect 597884 334170 597980 334226
rect 597360 334102 597980 334170
rect 597360 334046 597456 334102
rect 597512 334046 597580 334102
rect 597636 334046 597704 334102
rect 597760 334046 597828 334102
rect 597884 334046 597980 334102
rect 597360 333978 597980 334046
rect 597360 333922 597456 333978
rect 597512 333922 597580 333978
rect 597636 333922 597704 333978
rect 597760 333922 597828 333978
rect 597884 333922 597980 333978
rect 597360 316350 597980 333922
rect 597360 316294 597456 316350
rect 597512 316294 597580 316350
rect 597636 316294 597704 316350
rect 597760 316294 597828 316350
rect 597884 316294 597980 316350
rect 597360 316226 597980 316294
rect 597360 316170 597456 316226
rect 597512 316170 597580 316226
rect 597636 316170 597704 316226
rect 597760 316170 597828 316226
rect 597884 316170 597980 316226
rect 597360 316102 597980 316170
rect 597360 316046 597456 316102
rect 597512 316046 597580 316102
rect 597636 316046 597704 316102
rect 597760 316046 597828 316102
rect 597884 316046 597980 316102
rect 597360 315978 597980 316046
rect 597360 315922 597456 315978
rect 597512 315922 597580 315978
rect 597636 315922 597704 315978
rect 597760 315922 597828 315978
rect 597884 315922 597980 315978
rect 597360 298350 597980 315922
rect 597360 298294 597456 298350
rect 597512 298294 597580 298350
rect 597636 298294 597704 298350
rect 597760 298294 597828 298350
rect 597884 298294 597980 298350
rect 597360 298226 597980 298294
rect 597360 298170 597456 298226
rect 597512 298170 597580 298226
rect 597636 298170 597704 298226
rect 597760 298170 597828 298226
rect 597884 298170 597980 298226
rect 597360 298102 597980 298170
rect 597360 298046 597456 298102
rect 597512 298046 597580 298102
rect 597636 298046 597704 298102
rect 597760 298046 597828 298102
rect 597884 298046 597980 298102
rect 597360 297978 597980 298046
rect 597360 297922 597456 297978
rect 597512 297922 597580 297978
rect 597636 297922 597704 297978
rect 597760 297922 597828 297978
rect 597884 297922 597980 297978
rect 597360 280350 597980 297922
rect 597360 280294 597456 280350
rect 597512 280294 597580 280350
rect 597636 280294 597704 280350
rect 597760 280294 597828 280350
rect 597884 280294 597980 280350
rect 597360 280226 597980 280294
rect 597360 280170 597456 280226
rect 597512 280170 597580 280226
rect 597636 280170 597704 280226
rect 597760 280170 597828 280226
rect 597884 280170 597980 280226
rect 597360 280102 597980 280170
rect 597360 280046 597456 280102
rect 597512 280046 597580 280102
rect 597636 280046 597704 280102
rect 597760 280046 597828 280102
rect 597884 280046 597980 280102
rect 597360 279978 597980 280046
rect 597360 279922 597456 279978
rect 597512 279922 597580 279978
rect 597636 279922 597704 279978
rect 597760 279922 597828 279978
rect 597884 279922 597980 279978
rect 597360 262350 597980 279922
rect 597360 262294 597456 262350
rect 597512 262294 597580 262350
rect 597636 262294 597704 262350
rect 597760 262294 597828 262350
rect 597884 262294 597980 262350
rect 597360 262226 597980 262294
rect 597360 262170 597456 262226
rect 597512 262170 597580 262226
rect 597636 262170 597704 262226
rect 597760 262170 597828 262226
rect 597884 262170 597980 262226
rect 597360 262102 597980 262170
rect 597360 262046 597456 262102
rect 597512 262046 597580 262102
rect 597636 262046 597704 262102
rect 597760 262046 597828 262102
rect 597884 262046 597980 262102
rect 597360 261978 597980 262046
rect 597360 261922 597456 261978
rect 597512 261922 597580 261978
rect 597636 261922 597704 261978
rect 597760 261922 597828 261978
rect 597884 261922 597980 261978
rect 597360 244350 597980 261922
rect 597360 244294 597456 244350
rect 597512 244294 597580 244350
rect 597636 244294 597704 244350
rect 597760 244294 597828 244350
rect 597884 244294 597980 244350
rect 597360 244226 597980 244294
rect 597360 244170 597456 244226
rect 597512 244170 597580 244226
rect 597636 244170 597704 244226
rect 597760 244170 597828 244226
rect 597884 244170 597980 244226
rect 597360 244102 597980 244170
rect 597360 244046 597456 244102
rect 597512 244046 597580 244102
rect 597636 244046 597704 244102
rect 597760 244046 597828 244102
rect 597884 244046 597980 244102
rect 597360 243978 597980 244046
rect 597360 243922 597456 243978
rect 597512 243922 597580 243978
rect 597636 243922 597704 243978
rect 597760 243922 597828 243978
rect 597884 243922 597980 243978
rect 597360 226350 597980 243922
rect 597360 226294 597456 226350
rect 597512 226294 597580 226350
rect 597636 226294 597704 226350
rect 597760 226294 597828 226350
rect 597884 226294 597980 226350
rect 597360 226226 597980 226294
rect 597360 226170 597456 226226
rect 597512 226170 597580 226226
rect 597636 226170 597704 226226
rect 597760 226170 597828 226226
rect 597884 226170 597980 226226
rect 597360 226102 597980 226170
rect 597360 226046 597456 226102
rect 597512 226046 597580 226102
rect 597636 226046 597704 226102
rect 597760 226046 597828 226102
rect 597884 226046 597980 226102
rect 597360 225978 597980 226046
rect 597360 225922 597456 225978
rect 597512 225922 597580 225978
rect 597636 225922 597704 225978
rect 597760 225922 597828 225978
rect 597884 225922 597980 225978
rect 597360 208350 597980 225922
rect 597360 208294 597456 208350
rect 597512 208294 597580 208350
rect 597636 208294 597704 208350
rect 597760 208294 597828 208350
rect 597884 208294 597980 208350
rect 597360 208226 597980 208294
rect 597360 208170 597456 208226
rect 597512 208170 597580 208226
rect 597636 208170 597704 208226
rect 597760 208170 597828 208226
rect 597884 208170 597980 208226
rect 597360 208102 597980 208170
rect 597360 208046 597456 208102
rect 597512 208046 597580 208102
rect 597636 208046 597704 208102
rect 597760 208046 597828 208102
rect 597884 208046 597980 208102
rect 597360 207978 597980 208046
rect 597360 207922 597456 207978
rect 597512 207922 597580 207978
rect 597636 207922 597704 207978
rect 597760 207922 597828 207978
rect 597884 207922 597980 207978
rect 597360 190350 597980 207922
rect 597360 190294 597456 190350
rect 597512 190294 597580 190350
rect 597636 190294 597704 190350
rect 597760 190294 597828 190350
rect 597884 190294 597980 190350
rect 597360 190226 597980 190294
rect 597360 190170 597456 190226
rect 597512 190170 597580 190226
rect 597636 190170 597704 190226
rect 597760 190170 597828 190226
rect 597884 190170 597980 190226
rect 597360 190102 597980 190170
rect 597360 190046 597456 190102
rect 597512 190046 597580 190102
rect 597636 190046 597704 190102
rect 597760 190046 597828 190102
rect 597884 190046 597980 190102
rect 597360 189978 597980 190046
rect 597360 189922 597456 189978
rect 597512 189922 597580 189978
rect 597636 189922 597704 189978
rect 597760 189922 597828 189978
rect 597884 189922 597980 189978
rect 597360 172350 597980 189922
rect 597360 172294 597456 172350
rect 597512 172294 597580 172350
rect 597636 172294 597704 172350
rect 597760 172294 597828 172350
rect 597884 172294 597980 172350
rect 597360 172226 597980 172294
rect 597360 172170 597456 172226
rect 597512 172170 597580 172226
rect 597636 172170 597704 172226
rect 597760 172170 597828 172226
rect 597884 172170 597980 172226
rect 597360 172102 597980 172170
rect 597360 172046 597456 172102
rect 597512 172046 597580 172102
rect 597636 172046 597704 172102
rect 597760 172046 597828 172102
rect 597884 172046 597980 172102
rect 597360 171978 597980 172046
rect 597360 171922 597456 171978
rect 597512 171922 597580 171978
rect 597636 171922 597704 171978
rect 597760 171922 597828 171978
rect 597884 171922 597980 171978
rect 597360 154350 597980 171922
rect 597360 154294 597456 154350
rect 597512 154294 597580 154350
rect 597636 154294 597704 154350
rect 597760 154294 597828 154350
rect 597884 154294 597980 154350
rect 597360 154226 597980 154294
rect 597360 154170 597456 154226
rect 597512 154170 597580 154226
rect 597636 154170 597704 154226
rect 597760 154170 597828 154226
rect 597884 154170 597980 154226
rect 597360 154102 597980 154170
rect 597360 154046 597456 154102
rect 597512 154046 597580 154102
rect 597636 154046 597704 154102
rect 597760 154046 597828 154102
rect 597884 154046 597980 154102
rect 597360 153978 597980 154046
rect 597360 153922 597456 153978
rect 597512 153922 597580 153978
rect 597636 153922 597704 153978
rect 597760 153922 597828 153978
rect 597884 153922 597980 153978
rect 597360 136350 597980 153922
rect 597360 136294 597456 136350
rect 597512 136294 597580 136350
rect 597636 136294 597704 136350
rect 597760 136294 597828 136350
rect 597884 136294 597980 136350
rect 597360 136226 597980 136294
rect 597360 136170 597456 136226
rect 597512 136170 597580 136226
rect 597636 136170 597704 136226
rect 597760 136170 597828 136226
rect 597884 136170 597980 136226
rect 597360 136102 597980 136170
rect 597360 136046 597456 136102
rect 597512 136046 597580 136102
rect 597636 136046 597704 136102
rect 597760 136046 597828 136102
rect 597884 136046 597980 136102
rect 597360 135978 597980 136046
rect 597360 135922 597456 135978
rect 597512 135922 597580 135978
rect 597636 135922 597704 135978
rect 597760 135922 597828 135978
rect 597884 135922 597980 135978
rect 597360 118350 597980 135922
rect 597360 118294 597456 118350
rect 597512 118294 597580 118350
rect 597636 118294 597704 118350
rect 597760 118294 597828 118350
rect 597884 118294 597980 118350
rect 597360 118226 597980 118294
rect 597360 118170 597456 118226
rect 597512 118170 597580 118226
rect 597636 118170 597704 118226
rect 597760 118170 597828 118226
rect 597884 118170 597980 118226
rect 597360 118102 597980 118170
rect 597360 118046 597456 118102
rect 597512 118046 597580 118102
rect 597636 118046 597704 118102
rect 597760 118046 597828 118102
rect 597884 118046 597980 118102
rect 597360 117978 597980 118046
rect 597360 117922 597456 117978
rect 597512 117922 597580 117978
rect 597636 117922 597704 117978
rect 597760 117922 597828 117978
rect 597884 117922 597980 117978
rect 597360 100350 597980 117922
rect 597360 100294 597456 100350
rect 597512 100294 597580 100350
rect 597636 100294 597704 100350
rect 597760 100294 597828 100350
rect 597884 100294 597980 100350
rect 597360 100226 597980 100294
rect 597360 100170 597456 100226
rect 597512 100170 597580 100226
rect 597636 100170 597704 100226
rect 597760 100170 597828 100226
rect 597884 100170 597980 100226
rect 597360 100102 597980 100170
rect 597360 100046 597456 100102
rect 597512 100046 597580 100102
rect 597636 100046 597704 100102
rect 597760 100046 597828 100102
rect 597884 100046 597980 100102
rect 597360 99978 597980 100046
rect 597360 99922 597456 99978
rect 597512 99922 597580 99978
rect 597636 99922 597704 99978
rect 597760 99922 597828 99978
rect 597884 99922 597980 99978
rect 597360 82350 597980 99922
rect 597360 82294 597456 82350
rect 597512 82294 597580 82350
rect 597636 82294 597704 82350
rect 597760 82294 597828 82350
rect 597884 82294 597980 82350
rect 597360 82226 597980 82294
rect 597360 82170 597456 82226
rect 597512 82170 597580 82226
rect 597636 82170 597704 82226
rect 597760 82170 597828 82226
rect 597884 82170 597980 82226
rect 597360 82102 597980 82170
rect 597360 82046 597456 82102
rect 597512 82046 597580 82102
rect 597636 82046 597704 82102
rect 597760 82046 597828 82102
rect 597884 82046 597980 82102
rect 597360 81978 597980 82046
rect 597360 81922 597456 81978
rect 597512 81922 597580 81978
rect 597636 81922 597704 81978
rect 597760 81922 597828 81978
rect 597884 81922 597980 81978
rect 597360 64350 597980 81922
rect 597360 64294 597456 64350
rect 597512 64294 597580 64350
rect 597636 64294 597704 64350
rect 597760 64294 597828 64350
rect 597884 64294 597980 64350
rect 597360 64226 597980 64294
rect 597360 64170 597456 64226
rect 597512 64170 597580 64226
rect 597636 64170 597704 64226
rect 597760 64170 597828 64226
rect 597884 64170 597980 64226
rect 597360 64102 597980 64170
rect 597360 64046 597456 64102
rect 597512 64046 597580 64102
rect 597636 64046 597704 64102
rect 597760 64046 597828 64102
rect 597884 64046 597980 64102
rect 597360 63978 597980 64046
rect 597360 63922 597456 63978
rect 597512 63922 597580 63978
rect 597636 63922 597704 63978
rect 597760 63922 597828 63978
rect 597884 63922 597980 63978
rect 597360 46350 597980 63922
rect 597360 46294 597456 46350
rect 597512 46294 597580 46350
rect 597636 46294 597704 46350
rect 597760 46294 597828 46350
rect 597884 46294 597980 46350
rect 597360 46226 597980 46294
rect 597360 46170 597456 46226
rect 597512 46170 597580 46226
rect 597636 46170 597704 46226
rect 597760 46170 597828 46226
rect 597884 46170 597980 46226
rect 597360 46102 597980 46170
rect 597360 46046 597456 46102
rect 597512 46046 597580 46102
rect 597636 46046 597704 46102
rect 597760 46046 597828 46102
rect 597884 46046 597980 46102
rect 597360 45978 597980 46046
rect 597360 45922 597456 45978
rect 597512 45922 597580 45978
rect 597636 45922 597704 45978
rect 597760 45922 597828 45978
rect 597884 45922 597980 45978
rect 597360 28350 597980 45922
rect 597360 28294 597456 28350
rect 597512 28294 597580 28350
rect 597636 28294 597704 28350
rect 597760 28294 597828 28350
rect 597884 28294 597980 28350
rect 597360 28226 597980 28294
rect 597360 28170 597456 28226
rect 597512 28170 597580 28226
rect 597636 28170 597704 28226
rect 597760 28170 597828 28226
rect 597884 28170 597980 28226
rect 597360 28102 597980 28170
rect 597360 28046 597456 28102
rect 597512 28046 597580 28102
rect 597636 28046 597704 28102
rect 597760 28046 597828 28102
rect 597884 28046 597980 28102
rect 597360 27978 597980 28046
rect 597360 27922 597456 27978
rect 597512 27922 597580 27978
rect 597636 27922 597704 27978
rect 597760 27922 597828 27978
rect 597884 27922 597980 27978
rect 597360 10350 597980 27922
rect 597360 10294 597456 10350
rect 597512 10294 597580 10350
rect 597636 10294 597704 10350
rect 597760 10294 597828 10350
rect 597884 10294 597980 10350
rect 597360 10226 597980 10294
rect 597360 10170 597456 10226
rect 597512 10170 597580 10226
rect 597636 10170 597704 10226
rect 597760 10170 597828 10226
rect 597884 10170 597980 10226
rect 597360 10102 597980 10170
rect 597360 10046 597456 10102
rect 597512 10046 597580 10102
rect 597636 10046 597704 10102
rect 597760 10046 597828 10102
rect 597884 10046 597980 10102
rect 597360 9978 597980 10046
rect 597360 9922 597456 9978
rect 597512 9922 597580 9978
rect 597636 9922 597704 9978
rect 597760 9922 597828 9978
rect 597884 9922 597980 9978
rect 592818 -1176 592914 -1120
rect 592970 -1176 593038 -1120
rect 593094 -1176 593162 -1120
rect 593218 -1176 593286 -1120
rect 593342 -1176 593438 -1120
rect 592818 -1244 593438 -1176
rect 592818 -1300 592914 -1244
rect 592970 -1300 593038 -1244
rect 593094 -1300 593162 -1244
rect 593218 -1300 593286 -1244
rect 593342 -1300 593438 -1244
rect 592818 -1368 593438 -1300
rect 592818 -1424 592914 -1368
rect 592970 -1424 593038 -1368
rect 593094 -1424 593162 -1368
rect 593218 -1424 593286 -1368
rect 593342 -1424 593438 -1368
rect 592818 -1492 593438 -1424
rect 592818 -1548 592914 -1492
rect 592970 -1548 593038 -1492
rect 593094 -1548 593162 -1492
rect 593218 -1548 593286 -1492
rect 593342 -1548 593438 -1492
rect 592818 -1644 593438 -1548
rect 597360 -1120 597980 9922
rect 597360 -1176 597456 -1120
rect 597512 -1176 597580 -1120
rect 597636 -1176 597704 -1120
rect 597760 -1176 597828 -1120
rect 597884 -1176 597980 -1120
rect 597360 -1244 597980 -1176
rect 597360 -1300 597456 -1244
rect 597512 -1300 597580 -1244
rect 597636 -1300 597704 -1244
rect 597760 -1300 597828 -1244
rect 597884 -1300 597980 -1244
rect 597360 -1368 597980 -1300
rect 597360 -1424 597456 -1368
rect 597512 -1424 597580 -1368
rect 597636 -1424 597704 -1368
rect 597760 -1424 597828 -1368
rect 597884 -1424 597980 -1368
rect 597360 -1492 597980 -1424
rect 597360 -1548 597456 -1492
rect 597512 -1548 597580 -1492
rect 597636 -1548 597704 -1492
rect 597760 -1548 597828 -1492
rect 597884 -1548 597980 -1492
rect 597360 -1644 597980 -1548
<< via4 >>
rect -1820 598116 -1764 598172
rect -1696 598116 -1640 598172
rect -1572 598116 -1516 598172
rect -1448 598116 -1392 598172
rect -1820 597992 -1764 598048
rect -1696 597992 -1640 598048
rect -1572 597992 -1516 598048
rect -1448 597992 -1392 598048
rect -1820 597868 -1764 597924
rect -1696 597868 -1640 597924
rect -1572 597868 -1516 597924
rect -1448 597868 -1392 597924
rect -1820 597744 -1764 597800
rect -1696 597744 -1640 597800
rect -1572 597744 -1516 597800
rect -1448 597744 -1392 597800
rect -1820 586294 -1764 586350
rect -1696 586294 -1640 586350
rect -1572 586294 -1516 586350
rect -1448 586294 -1392 586350
rect -1820 586170 -1764 586226
rect -1696 586170 -1640 586226
rect -1572 586170 -1516 586226
rect -1448 586170 -1392 586226
rect -1820 586046 -1764 586102
rect -1696 586046 -1640 586102
rect -1572 586046 -1516 586102
rect -1448 586046 -1392 586102
rect -1820 585922 -1764 585978
rect -1696 585922 -1640 585978
rect -1572 585922 -1516 585978
rect -1448 585922 -1392 585978
rect -1820 568294 -1764 568350
rect -1696 568294 -1640 568350
rect -1572 568294 -1516 568350
rect -1448 568294 -1392 568350
rect -1820 568170 -1764 568226
rect -1696 568170 -1640 568226
rect -1572 568170 -1516 568226
rect -1448 568170 -1392 568226
rect -1820 568046 -1764 568102
rect -1696 568046 -1640 568102
rect -1572 568046 -1516 568102
rect -1448 568046 -1392 568102
rect -1820 567922 -1764 567978
rect -1696 567922 -1640 567978
rect -1572 567922 -1516 567978
rect -1448 567922 -1392 567978
rect -1820 550294 -1764 550350
rect -1696 550294 -1640 550350
rect -1572 550294 -1516 550350
rect -1448 550294 -1392 550350
rect -1820 550170 -1764 550226
rect -1696 550170 -1640 550226
rect -1572 550170 -1516 550226
rect -1448 550170 -1392 550226
rect -1820 550046 -1764 550102
rect -1696 550046 -1640 550102
rect -1572 550046 -1516 550102
rect -1448 550046 -1392 550102
rect -1820 549922 -1764 549978
rect -1696 549922 -1640 549978
rect -1572 549922 -1516 549978
rect -1448 549922 -1392 549978
rect -1820 532294 -1764 532350
rect -1696 532294 -1640 532350
rect -1572 532294 -1516 532350
rect -1448 532294 -1392 532350
rect -1820 532170 -1764 532226
rect -1696 532170 -1640 532226
rect -1572 532170 -1516 532226
rect -1448 532170 -1392 532226
rect -1820 532046 -1764 532102
rect -1696 532046 -1640 532102
rect -1572 532046 -1516 532102
rect -1448 532046 -1392 532102
rect -1820 531922 -1764 531978
rect -1696 531922 -1640 531978
rect -1572 531922 -1516 531978
rect -1448 531922 -1392 531978
rect -1820 514294 -1764 514350
rect -1696 514294 -1640 514350
rect -1572 514294 -1516 514350
rect -1448 514294 -1392 514350
rect -1820 514170 -1764 514226
rect -1696 514170 -1640 514226
rect -1572 514170 -1516 514226
rect -1448 514170 -1392 514226
rect -1820 514046 -1764 514102
rect -1696 514046 -1640 514102
rect -1572 514046 -1516 514102
rect -1448 514046 -1392 514102
rect -1820 513922 -1764 513978
rect -1696 513922 -1640 513978
rect -1572 513922 -1516 513978
rect -1448 513922 -1392 513978
rect -1820 496294 -1764 496350
rect -1696 496294 -1640 496350
rect -1572 496294 -1516 496350
rect -1448 496294 -1392 496350
rect -1820 496170 -1764 496226
rect -1696 496170 -1640 496226
rect -1572 496170 -1516 496226
rect -1448 496170 -1392 496226
rect -1820 496046 -1764 496102
rect -1696 496046 -1640 496102
rect -1572 496046 -1516 496102
rect -1448 496046 -1392 496102
rect -1820 495922 -1764 495978
rect -1696 495922 -1640 495978
rect -1572 495922 -1516 495978
rect -1448 495922 -1392 495978
rect -1820 478294 -1764 478350
rect -1696 478294 -1640 478350
rect -1572 478294 -1516 478350
rect -1448 478294 -1392 478350
rect -1820 478170 -1764 478226
rect -1696 478170 -1640 478226
rect -1572 478170 -1516 478226
rect -1448 478170 -1392 478226
rect -1820 478046 -1764 478102
rect -1696 478046 -1640 478102
rect -1572 478046 -1516 478102
rect -1448 478046 -1392 478102
rect -1820 477922 -1764 477978
rect -1696 477922 -1640 477978
rect -1572 477922 -1516 477978
rect -1448 477922 -1392 477978
rect -1820 460294 -1764 460350
rect -1696 460294 -1640 460350
rect -1572 460294 -1516 460350
rect -1448 460294 -1392 460350
rect -1820 460170 -1764 460226
rect -1696 460170 -1640 460226
rect -1572 460170 -1516 460226
rect -1448 460170 -1392 460226
rect -1820 460046 -1764 460102
rect -1696 460046 -1640 460102
rect -1572 460046 -1516 460102
rect -1448 460046 -1392 460102
rect -1820 459922 -1764 459978
rect -1696 459922 -1640 459978
rect -1572 459922 -1516 459978
rect -1448 459922 -1392 459978
rect -1820 442294 -1764 442350
rect -1696 442294 -1640 442350
rect -1572 442294 -1516 442350
rect -1448 442294 -1392 442350
rect -1820 442170 -1764 442226
rect -1696 442170 -1640 442226
rect -1572 442170 -1516 442226
rect -1448 442170 -1392 442226
rect -1820 442046 -1764 442102
rect -1696 442046 -1640 442102
rect -1572 442046 -1516 442102
rect -1448 442046 -1392 442102
rect -1820 441922 -1764 441978
rect -1696 441922 -1640 441978
rect -1572 441922 -1516 441978
rect -1448 441922 -1392 441978
rect -1820 424294 -1764 424350
rect -1696 424294 -1640 424350
rect -1572 424294 -1516 424350
rect -1448 424294 -1392 424350
rect -1820 424170 -1764 424226
rect -1696 424170 -1640 424226
rect -1572 424170 -1516 424226
rect -1448 424170 -1392 424226
rect -1820 424046 -1764 424102
rect -1696 424046 -1640 424102
rect -1572 424046 -1516 424102
rect -1448 424046 -1392 424102
rect -1820 423922 -1764 423978
rect -1696 423922 -1640 423978
rect -1572 423922 -1516 423978
rect -1448 423922 -1392 423978
rect -1820 406294 -1764 406350
rect -1696 406294 -1640 406350
rect -1572 406294 -1516 406350
rect -1448 406294 -1392 406350
rect -1820 406170 -1764 406226
rect -1696 406170 -1640 406226
rect -1572 406170 -1516 406226
rect -1448 406170 -1392 406226
rect -1820 406046 -1764 406102
rect -1696 406046 -1640 406102
rect -1572 406046 -1516 406102
rect -1448 406046 -1392 406102
rect -1820 405922 -1764 405978
rect -1696 405922 -1640 405978
rect -1572 405922 -1516 405978
rect -1448 405922 -1392 405978
rect -1820 388294 -1764 388350
rect -1696 388294 -1640 388350
rect -1572 388294 -1516 388350
rect -1448 388294 -1392 388350
rect -1820 388170 -1764 388226
rect -1696 388170 -1640 388226
rect -1572 388170 -1516 388226
rect -1448 388170 -1392 388226
rect -1820 388046 -1764 388102
rect -1696 388046 -1640 388102
rect -1572 388046 -1516 388102
rect -1448 388046 -1392 388102
rect -1820 387922 -1764 387978
rect -1696 387922 -1640 387978
rect -1572 387922 -1516 387978
rect -1448 387922 -1392 387978
rect -1820 370294 -1764 370350
rect -1696 370294 -1640 370350
rect -1572 370294 -1516 370350
rect -1448 370294 -1392 370350
rect -1820 370170 -1764 370226
rect -1696 370170 -1640 370226
rect -1572 370170 -1516 370226
rect -1448 370170 -1392 370226
rect -1820 370046 -1764 370102
rect -1696 370046 -1640 370102
rect -1572 370046 -1516 370102
rect -1448 370046 -1392 370102
rect -1820 369922 -1764 369978
rect -1696 369922 -1640 369978
rect -1572 369922 -1516 369978
rect -1448 369922 -1392 369978
rect -1820 352294 -1764 352350
rect -1696 352294 -1640 352350
rect -1572 352294 -1516 352350
rect -1448 352294 -1392 352350
rect -1820 352170 -1764 352226
rect -1696 352170 -1640 352226
rect -1572 352170 -1516 352226
rect -1448 352170 -1392 352226
rect -1820 352046 -1764 352102
rect -1696 352046 -1640 352102
rect -1572 352046 -1516 352102
rect -1448 352046 -1392 352102
rect -1820 351922 -1764 351978
rect -1696 351922 -1640 351978
rect -1572 351922 -1516 351978
rect -1448 351922 -1392 351978
rect -1820 334294 -1764 334350
rect -1696 334294 -1640 334350
rect -1572 334294 -1516 334350
rect -1448 334294 -1392 334350
rect -1820 334170 -1764 334226
rect -1696 334170 -1640 334226
rect -1572 334170 -1516 334226
rect -1448 334170 -1392 334226
rect -1820 334046 -1764 334102
rect -1696 334046 -1640 334102
rect -1572 334046 -1516 334102
rect -1448 334046 -1392 334102
rect -1820 333922 -1764 333978
rect -1696 333922 -1640 333978
rect -1572 333922 -1516 333978
rect -1448 333922 -1392 333978
rect -1820 316294 -1764 316350
rect -1696 316294 -1640 316350
rect -1572 316294 -1516 316350
rect -1448 316294 -1392 316350
rect -1820 316170 -1764 316226
rect -1696 316170 -1640 316226
rect -1572 316170 -1516 316226
rect -1448 316170 -1392 316226
rect -1820 316046 -1764 316102
rect -1696 316046 -1640 316102
rect -1572 316046 -1516 316102
rect -1448 316046 -1392 316102
rect -1820 315922 -1764 315978
rect -1696 315922 -1640 315978
rect -1572 315922 -1516 315978
rect -1448 315922 -1392 315978
rect -1820 298294 -1764 298350
rect -1696 298294 -1640 298350
rect -1572 298294 -1516 298350
rect -1448 298294 -1392 298350
rect -1820 298170 -1764 298226
rect -1696 298170 -1640 298226
rect -1572 298170 -1516 298226
rect -1448 298170 -1392 298226
rect -1820 298046 -1764 298102
rect -1696 298046 -1640 298102
rect -1572 298046 -1516 298102
rect -1448 298046 -1392 298102
rect -1820 297922 -1764 297978
rect -1696 297922 -1640 297978
rect -1572 297922 -1516 297978
rect -1448 297922 -1392 297978
rect -1820 280294 -1764 280350
rect -1696 280294 -1640 280350
rect -1572 280294 -1516 280350
rect -1448 280294 -1392 280350
rect -1820 280170 -1764 280226
rect -1696 280170 -1640 280226
rect -1572 280170 -1516 280226
rect -1448 280170 -1392 280226
rect -1820 280046 -1764 280102
rect -1696 280046 -1640 280102
rect -1572 280046 -1516 280102
rect -1448 280046 -1392 280102
rect -1820 279922 -1764 279978
rect -1696 279922 -1640 279978
rect -1572 279922 -1516 279978
rect -1448 279922 -1392 279978
rect -1820 262294 -1764 262350
rect -1696 262294 -1640 262350
rect -1572 262294 -1516 262350
rect -1448 262294 -1392 262350
rect -1820 262170 -1764 262226
rect -1696 262170 -1640 262226
rect -1572 262170 -1516 262226
rect -1448 262170 -1392 262226
rect -1820 262046 -1764 262102
rect -1696 262046 -1640 262102
rect -1572 262046 -1516 262102
rect -1448 262046 -1392 262102
rect -1820 261922 -1764 261978
rect -1696 261922 -1640 261978
rect -1572 261922 -1516 261978
rect -1448 261922 -1392 261978
rect -1820 244294 -1764 244350
rect -1696 244294 -1640 244350
rect -1572 244294 -1516 244350
rect -1448 244294 -1392 244350
rect -1820 244170 -1764 244226
rect -1696 244170 -1640 244226
rect -1572 244170 -1516 244226
rect -1448 244170 -1392 244226
rect -1820 244046 -1764 244102
rect -1696 244046 -1640 244102
rect -1572 244046 -1516 244102
rect -1448 244046 -1392 244102
rect -1820 243922 -1764 243978
rect -1696 243922 -1640 243978
rect -1572 243922 -1516 243978
rect -1448 243922 -1392 243978
rect -1820 226294 -1764 226350
rect -1696 226294 -1640 226350
rect -1572 226294 -1516 226350
rect -1448 226294 -1392 226350
rect -1820 226170 -1764 226226
rect -1696 226170 -1640 226226
rect -1572 226170 -1516 226226
rect -1448 226170 -1392 226226
rect -1820 226046 -1764 226102
rect -1696 226046 -1640 226102
rect -1572 226046 -1516 226102
rect -1448 226046 -1392 226102
rect -1820 225922 -1764 225978
rect -1696 225922 -1640 225978
rect -1572 225922 -1516 225978
rect -1448 225922 -1392 225978
rect -1820 208294 -1764 208350
rect -1696 208294 -1640 208350
rect -1572 208294 -1516 208350
rect -1448 208294 -1392 208350
rect -1820 208170 -1764 208226
rect -1696 208170 -1640 208226
rect -1572 208170 -1516 208226
rect -1448 208170 -1392 208226
rect -1820 208046 -1764 208102
rect -1696 208046 -1640 208102
rect -1572 208046 -1516 208102
rect -1448 208046 -1392 208102
rect -1820 207922 -1764 207978
rect -1696 207922 -1640 207978
rect -1572 207922 -1516 207978
rect -1448 207922 -1392 207978
rect -1820 190294 -1764 190350
rect -1696 190294 -1640 190350
rect -1572 190294 -1516 190350
rect -1448 190294 -1392 190350
rect -1820 190170 -1764 190226
rect -1696 190170 -1640 190226
rect -1572 190170 -1516 190226
rect -1448 190170 -1392 190226
rect -1820 190046 -1764 190102
rect -1696 190046 -1640 190102
rect -1572 190046 -1516 190102
rect -1448 190046 -1392 190102
rect -1820 189922 -1764 189978
rect -1696 189922 -1640 189978
rect -1572 189922 -1516 189978
rect -1448 189922 -1392 189978
rect -1820 172294 -1764 172350
rect -1696 172294 -1640 172350
rect -1572 172294 -1516 172350
rect -1448 172294 -1392 172350
rect -1820 172170 -1764 172226
rect -1696 172170 -1640 172226
rect -1572 172170 -1516 172226
rect -1448 172170 -1392 172226
rect -1820 172046 -1764 172102
rect -1696 172046 -1640 172102
rect -1572 172046 -1516 172102
rect -1448 172046 -1392 172102
rect -1820 171922 -1764 171978
rect -1696 171922 -1640 171978
rect -1572 171922 -1516 171978
rect -1448 171922 -1392 171978
rect -1820 154294 -1764 154350
rect -1696 154294 -1640 154350
rect -1572 154294 -1516 154350
rect -1448 154294 -1392 154350
rect -1820 154170 -1764 154226
rect -1696 154170 -1640 154226
rect -1572 154170 -1516 154226
rect -1448 154170 -1392 154226
rect -1820 154046 -1764 154102
rect -1696 154046 -1640 154102
rect -1572 154046 -1516 154102
rect -1448 154046 -1392 154102
rect -1820 153922 -1764 153978
rect -1696 153922 -1640 153978
rect -1572 153922 -1516 153978
rect -1448 153922 -1392 153978
rect -1820 136294 -1764 136350
rect -1696 136294 -1640 136350
rect -1572 136294 -1516 136350
rect -1448 136294 -1392 136350
rect -1820 136170 -1764 136226
rect -1696 136170 -1640 136226
rect -1572 136170 -1516 136226
rect -1448 136170 -1392 136226
rect -1820 136046 -1764 136102
rect -1696 136046 -1640 136102
rect -1572 136046 -1516 136102
rect -1448 136046 -1392 136102
rect -1820 135922 -1764 135978
rect -1696 135922 -1640 135978
rect -1572 135922 -1516 135978
rect -1448 135922 -1392 135978
rect -1820 118294 -1764 118350
rect -1696 118294 -1640 118350
rect -1572 118294 -1516 118350
rect -1448 118294 -1392 118350
rect -1820 118170 -1764 118226
rect -1696 118170 -1640 118226
rect -1572 118170 -1516 118226
rect -1448 118170 -1392 118226
rect -1820 118046 -1764 118102
rect -1696 118046 -1640 118102
rect -1572 118046 -1516 118102
rect -1448 118046 -1392 118102
rect -1820 117922 -1764 117978
rect -1696 117922 -1640 117978
rect -1572 117922 -1516 117978
rect -1448 117922 -1392 117978
rect -1820 100294 -1764 100350
rect -1696 100294 -1640 100350
rect -1572 100294 -1516 100350
rect -1448 100294 -1392 100350
rect -1820 100170 -1764 100226
rect -1696 100170 -1640 100226
rect -1572 100170 -1516 100226
rect -1448 100170 -1392 100226
rect -1820 100046 -1764 100102
rect -1696 100046 -1640 100102
rect -1572 100046 -1516 100102
rect -1448 100046 -1392 100102
rect -1820 99922 -1764 99978
rect -1696 99922 -1640 99978
rect -1572 99922 -1516 99978
rect -1448 99922 -1392 99978
rect -1820 82294 -1764 82350
rect -1696 82294 -1640 82350
rect -1572 82294 -1516 82350
rect -1448 82294 -1392 82350
rect -1820 82170 -1764 82226
rect -1696 82170 -1640 82226
rect -1572 82170 -1516 82226
rect -1448 82170 -1392 82226
rect -1820 82046 -1764 82102
rect -1696 82046 -1640 82102
rect -1572 82046 -1516 82102
rect -1448 82046 -1392 82102
rect -1820 81922 -1764 81978
rect -1696 81922 -1640 81978
rect -1572 81922 -1516 81978
rect -1448 81922 -1392 81978
rect -1820 64294 -1764 64350
rect -1696 64294 -1640 64350
rect -1572 64294 -1516 64350
rect -1448 64294 -1392 64350
rect -1820 64170 -1764 64226
rect -1696 64170 -1640 64226
rect -1572 64170 -1516 64226
rect -1448 64170 -1392 64226
rect -1820 64046 -1764 64102
rect -1696 64046 -1640 64102
rect -1572 64046 -1516 64102
rect -1448 64046 -1392 64102
rect -1820 63922 -1764 63978
rect -1696 63922 -1640 63978
rect -1572 63922 -1516 63978
rect -1448 63922 -1392 63978
rect -1820 46294 -1764 46350
rect -1696 46294 -1640 46350
rect -1572 46294 -1516 46350
rect -1448 46294 -1392 46350
rect -1820 46170 -1764 46226
rect -1696 46170 -1640 46226
rect -1572 46170 -1516 46226
rect -1448 46170 -1392 46226
rect -1820 46046 -1764 46102
rect -1696 46046 -1640 46102
rect -1572 46046 -1516 46102
rect -1448 46046 -1392 46102
rect -1820 45922 -1764 45978
rect -1696 45922 -1640 45978
rect -1572 45922 -1516 45978
rect -1448 45922 -1392 45978
rect -1820 28294 -1764 28350
rect -1696 28294 -1640 28350
rect -1572 28294 -1516 28350
rect -1448 28294 -1392 28350
rect -1820 28170 -1764 28226
rect -1696 28170 -1640 28226
rect -1572 28170 -1516 28226
rect -1448 28170 -1392 28226
rect -1820 28046 -1764 28102
rect -1696 28046 -1640 28102
rect -1572 28046 -1516 28102
rect -1448 28046 -1392 28102
rect -1820 27922 -1764 27978
rect -1696 27922 -1640 27978
rect -1572 27922 -1516 27978
rect -1448 27922 -1392 27978
rect -1820 10294 -1764 10350
rect -1696 10294 -1640 10350
rect -1572 10294 -1516 10350
rect -1448 10294 -1392 10350
rect -1820 10170 -1764 10226
rect -1696 10170 -1640 10226
rect -1572 10170 -1516 10226
rect -1448 10170 -1392 10226
rect -1820 10046 -1764 10102
rect -1696 10046 -1640 10102
rect -1572 10046 -1516 10102
rect -1448 10046 -1392 10102
rect -1820 9922 -1764 9978
rect -1696 9922 -1640 9978
rect -1572 9922 -1516 9978
rect -1448 9922 -1392 9978
rect -860 597156 -804 597212
rect -736 597156 -680 597212
rect -612 597156 -556 597212
rect -488 597156 -432 597212
rect -860 597032 -804 597088
rect -736 597032 -680 597088
rect -612 597032 -556 597088
rect -488 597032 -432 597088
rect -860 596908 -804 596964
rect -736 596908 -680 596964
rect -612 596908 -556 596964
rect -488 596908 -432 596964
rect -860 596784 -804 596840
rect -736 596784 -680 596840
rect -612 596784 -556 596840
rect -488 596784 -432 596840
rect 5514 597156 5570 597212
rect 5638 597156 5694 597212
rect 5762 597156 5818 597212
rect 5886 597156 5942 597212
rect 5514 597032 5570 597088
rect 5638 597032 5694 597088
rect 5762 597032 5818 597088
rect 5886 597032 5942 597088
rect 5514 596908 5570 596964
rect 5638 596908 5694 596964
rect 5762 596908 5818 596964
rect 5886 596908 5942 596964
rect 5514 596784 5570 596840
rect 5638 596784 5694 596840
rect 5762 596784 5818 596840
rect 5886 596784 5942 596840
rect -860 580294 -804 580350
rect -736 580294 -680 580350
rect -612 580294 -556 580350
rect -488 580294 -432 580350
rect -860 580170 -804 580226
rect -736 580170 -680 580226
rect -612 580170 -556 580226
rect -488 580170 -432 580226
rect -860 580046 -804 580102
rect -736 580046 -680 580102
rect -612 580046 -556 580102
rect -488 580046 -432 580102
rect -860 579922 -804 579978
rect -736 579922 -680 579978
rect -612 579922 -556 579978
rect -488 579922 -432 579978
rect -860 562294 -804 562350
rect -736 562294 -680 562350
rect -612 562294 -556 562350
rect -488 562294 -432 562350
rect -860 562170 -804 562226
rect -736 562170 -680 562226
rect -612 562170 -556 562226
rect -488 562170 -432 562226
rect -860 562046 -804 562102
rect -736 562046 -680 562102
rect -612 562046 -556 562102
rect -488 562046 -432 562102
rect -860 561922 -804 561978
rect -736 561922 -680 561978
rect -612 561922 -556 561978
rect -488 561922 -432 561978
rect 5514 580294 5570 580350
rect 5638 580294 5694 580350
rect 5762 580294 5818 580350
rect 5886 580294 5942 580350
rect 5514 580170 5570 580226
rect 5638 580170 5694 580226
rect 5762 580170 5818 580226
rect 5886 580170 5942 580226
rect 5514 580046 5570 580102
rect 5638 580046 5694 580102
rect 5762 580046 5818 580102
rect 5886 580046 5942 580102
rect 5514 579922 5570 579978
rect 5638 579922 5694 579978
rect 5762 579922 5818 579978
rect 5886 579922 5942 579978
rect -860 544294 -804 544350
rect -736 544294 -680 544350
rect -612 544294 -556 544350
rect -488 544294 -432 544350
rect -860 544170 -804 544226
rect -736 544170 -680 544226
rect -612 544170 -556 544226
rect -488 544170 -432 544226
rect -860 544046 -804 544102
rect -736 544046 -680 544102
rect -612 544046 -556 544102
rect -488 544046 -432 544102
rect -860 543922 -804 543978
rect -736 543922 -680 543978
rect -612 543922 -556 543978
rect -488 543922 -432 543978
rect -860 526294 -804 526350
rect -736 526294 -680 526350
rect -612 526294 -556 526350
rect -488 526294 -432 526350
rect -860 526170 -804 526226
rect -736 526170 -680 526226
rect -612 526170 -556 526226
rect -488 526170 -432 526226
rect -860 526046 -804 526102
rect -736 526046 -680 526102
rect -612 526046 -556 526102
rect -488 526046 -432 526102
rect -860 525922 -804 525978
rect -736 525922 -680 525978
rect -612 525922 -556 525978
rect -488 525922 -432 525978
rect -860 508294 -804 508350
rect -736 508294 -680 508350
rect -612 508294 -556 508350
rect -488 508294 -432 508350
rect -860 508170 -804 508226
rect -736 508170 -680 508226
rect -612 508170 -556 508226
rect -488 508170 -432 508226
rect -860 508046 -804 508102
rect -736 508046 -680 508102
rect -612 508046 -556 508102
rect -488 508046 -432 508102
rect -860 507922 -804 507978
rect -736 507922 -680 507978
rect -612 507922 -556 507978
rect -488 507922 -432 507978
rect -860 490294 -804 490350
rect -736 490294 -680 490350
rect -612 490294 -556 490350
rect -488 490294 -432 490350
rect -860 490170 -804 490226
rect -736 490170 -680 490226
rect -612 490170 -556 490226
rect -488 490170 -432 490226
rect -860 490046 -804 490102
rect -736 490046 -680 490102
rect -612 490046 -556 490102
rect -488 490046 -432 490102
rect -860 489922 -804 489978
rect -736 489922 -680 489978
rect -612 489922 -556 489978
rect -488 489922 -432 489978
rect -860 472294 -804 472350
rect -736 472294 -680 472350
rect -612 472294 -556 472350
rect -488 472294 -432 472350
rect -860 472170 -804 472226
rect -736 472170 -680 472226
rect -612 472170 -556 472226
rect -488 472170 -432 472226
rect -860 472046 -804 472102
rect -736 472046 -680 472102
rect -612 472046 -556 472102
rect -488 472046 -432 472102
rect -860 471922 -804 471978
rect -736 471922 -680 471978
rect -612 471922 -556 471978
rect -488 471922 -432 471978
rect -860 454294 -804 454350
rect -736 454294 -680 454350
rect -612 454294 -556 454350
rect -488 454294 -432 454350
rect -860 454170 -804 454226
rect -736 454170 -680 454226
rect -612 454170 -556 454226
rect -488 454170 -432 454226
rect -860 454046 -804 454102
rect -736 454046 -680 454102
rect -612 454046 -556 454102
rect -488 454046 -432 454102
rect -860 453922 -804 453978
rect -736 453922 -680 453978
rect -612 453922 -556 453978
rect -488 453922 -432 453978
rect -860 436294 -804 436350
rect -736 436294 -680 436350
rect -612 436294 -556 436350
rect -488 436294 -432 436350
rect -860 436170 -804 436226
rect -736 436170 -680 436226
rect -612 436170 -556 436226
rect -488 436170 -432 436226
rect -860 436046 -804 436102
rect -736 436046 -680 436102
rect -612 436046 -556 436102
rect -488 436046 -432 436102
rect -860 435922 -804 435978
rect -736 435922 -680 435978
rect -612 435922 -556 435978
rect -488 435922 -432 435978
rect -860 418294 -804 418350
rect -736 418294 -680 418350
rect -612 418294 -556 418350
rect -488 418294 -432 418350
rect -860 418170 -804 418226
rect -736 418170 -680 418226
rect -612 418170 -556 418226
rect -488 418170 -432 418226
rect -860 418046 -804 418102
rect -736 418046 -680 418102
rect -612 418046 -556 418102
rect -488 418046 -432 418102
rect -860 417922 -804 417978
rect -736 417922 -680 417978
rect -612 417922 -556 417978
rect -488 417922 -432 417978
rect -860 400294 -804 400350
rect -736 400294 -680 400350
rect -612 400294 -556 400350
rect -488 400294 -432 400350
rect -860 400170 -804 400226
rect -736 400170 -680 400226
rect -612 400170 -556 400226
rect -488 400170 -432 400226
rect -860 400046 -804 400102
rect -736 400046 -680 400102
rect -612 400046 -556 400102
rect -488 400046 -432 400102
rect -860 399922 -804 399978
rect -736 399922 -680 399978
rect -612 399922 -556 399978
rect -488 399922 -432 399978
rect -860 382294 -804 382350
rect -736 382294 -680 382350
rect -612 382294 -556 382350
rect -488 382294 -432 382350
rect -860 382170 -804 382226
rect -736 382170 -680 382226
rect -612 382170 -556 382226
rect -488 382170 -432 382226
rect -860 382046 -804 382102
rect -736 382046 -680 382102
rect -612 382046 -556 382102
rect -488 382046 -432 382102
rect -860 381922 -804 381978
rect -736 381922 -680 381978
rect -612 381922 -556 381978
rect -488 381922 -432 381978
rect -860 364294 -804 364350
rect -736 364294 -680 364350
rect -612 364294 -556 364350
rect -488 364294 -432 364350
rect -860 364170 -804 364226
rect -736 364170 -680 364226
rect -612 364170 -556 364226
rect -488 364170 -432 364226
rect -860 364046 -804 364102
rect -736 364046 -680 364102
rect -612 364046 -556 364102
rect -488 364046 -432 364102
rect -860 363922 -804 363978
rect -736 363922 -680 363978
rect -612 363922 -556 363978
rect -488 363922 -432 363978
rect -860 346294 -804 346350
rect -736 346294 -680 346350
rect -612 346294 -556 346350
rect -488 346294 -432 346350
rect -860 346170 -804 346226
rect -736 346170 -680 346226
rect -612 346170 -556 346226
rect -488 346170 -432 346226
rect -860 346046 -804 346102
rect -736 346046 -680 346102
rect -612 346046 -556 346102
rect -488 346046 -432 346102
rect -860 345922 -804 345978
rect -736 345922 -680 345978
rect -612 345922 -556 345978
rect -488 345922 -432 345978
rect -860 328294 -804 328350
rect -736 328294 -680 328350
rect -612 328294 -556 328350
rect -488 328294 -432 328350
rect -860 328170 -804 328226
rect -736 328170 -680 328226
rect -612 328170 -556 328226
rect -488 328170 -432 328226
rect -860 328046 -804 328102
rect -736 328046 -680 328102
rect -612 328046 -556 328102
rect -488 328046 -432 328102
rect -860 327922 -804 327978
rect -736 327922 -680 327978
rect -612 327922 -556 327978
rect -488 327922 -432 327978
rect -860 310294 -804 310350
rect -736 310294 -680 310350
rect -612 310294 -556 310350
rect -488 310294 -432 310350
rect -860 310170 -804 310226
rect -736 310170 -680 310226
rect -612 310170 -556 310226
rect -488 310170 -432 310226
rect -860 310046 -804 310102
rect -736 310046 -680 310102
rect -612 310046 -556 310102
rect -488 310046 -432 310102
rect -860 309922 -804 309978
rect -736 309922 -680 309978
rect -612 309922 -556 309978
rect -488 309922 -432 309978
rect -860 292294 -804 292350
rect -736 292294 -680 292350
rect -612 292294 -556 292350
rect -488 292294 -432 292350
rect -860 292170 -804 292226
rect -736 292170 -680 292226
rect -612 292170 -556 292226
rect -488 292170 -432 292226
rect -860 292046 -804 292102
rect -736 292046 -680 292102
rect -612 292046 -556 292102
rect -488 292046 -432 292102
rect -860 291922 -804 291978
rect -736 291922 -680 291978
rect -612 291922 -556 291978
rect -488 291922 -432 291978
rect -860 274294 -804 274350
rect -736 274294 -680 274350
rect -612 274294 -556 274350
rect -488 274294 -432 274350
rect -860 274170 -804 274226
rect -736 274170 -680 274226
rect -612 274170 -556 274226
rect -488 274170 -432 274226
rect -860 274046 -804 274102
rect -736 274046 -680 274102
rect -612 274046 -556 274102
rect -488 274046 -432 274102
rect -860 273922 -804 273978
rect -736 273922 -680 273978
rect -612 273922 -556 273978
rect -488 273922 -432 273978
rect -860 256294 -804 256350
rect -736 256294 -680 256350
rect -612 256294 -556 256350
rect -488 256294 -432 256350
rect -860 256170 -804 256226
rect -736 256170 -680 256226
rect -612 256170 -556 256226
rect -488 256170 -432 256226
rect -860 256046 -804 256102
rect -736 256046 -680 256102
rect -612 256046 -556 256102
rect -488 256046 -432 256102
rect -860 255922 -804 255978
rect -736 255922 -680 255978
rect -612 255922 -556 255978
rect -488 255922 -432 255978
rect -860 238294 -804 238350
rect -736 238294 -680 238350
rect -612 238294 -556 238350
rect -488 238294 -432 238350
rect -860 238170 -804 238226
rect -736 238170 -680 238226
rect -612 238170 -556 238226
rect -488 238170 -432 238226
rect -860 238046 -804 238102
rect -736 238046 -680 238102
rect -612 238046 -556 238102
rect -488 238046 -432 238102
rect -860 237922 -804 237978
rect -736 237922 -680 237978
rect -612 237922 -556 237978
rect -488 237922 -432 237978
rect -860 220294 -804 220350
rect -736 220294 -680 220350
rect -612 220294 -556 220350
rect -488 220294 -432 220350
rect -860 220170 -804 220226
rect -736 220170 -680 220226
rect -612 220170 -556 220226
rect -488 220170 -432 220226
rect -860 220046 -804 220102
rect -736 220046 -680 220102
rect -612 220046 -556 220102
rect -488 220046 -432 220102
rect -860 219922 -804 219978
rect -736 219922 -680 219978
rect -612 219922 -556 219978
rect -488 219922 -432 219978
rect -860 202294 -804 202350
rect -736 202294 -680 202350
rect -612 202294 -556 202350
rect -488 202294 -432 202350
rect -860 202170 -804 202226
rect -736 202170 -680 202226
rect -612 202170 -556 202226
rect -488 202170 -432 202226
rect -860 202046 -804 202102
rect -736 202046 -680 202102
rect -612 202046 -556 202102
rect -488 202046 -432 202102
rect -860 201922 -804 201978
rect -736 201922 -680 201978
rect -612 201922 -556 201978
rect -488 201922 -432 201978
rect -860 184294 -804 184350
rect -736 184294 -680 184350
rect -612 184294 -556 184350
rect -488 184294 -432 184350
rect -860 184170 -804 184226
rect -736 184170 -680 184226
rect -612 184170 -556 184226
rect -488 184170 -432 184226
rect -860 184046 -804 184102
rect -736 184046 -680 184102
rect -612 184046 -556 184102
rect -488 184046 -432 184102
rect -860 183922 -804 183978
rect -736 183922 -680 183978
rect -612 183922 -556 183978
rect -488 183922 -432 183978
rect -860 166294 -804 166350
rect -736 166294 -680 166350
rect -612 166294 -556 166350
rect -488 166294 -432 166350
rect -860 166170 -804 166226
rect -736 166170 -680 166226
rect -612 166170 -556 166226
rect -488 166170 -432 166226
rect -860 166046 -804 166102
rect -736 166046 -680 166102
rect -612 166046 -556 166102
rect -488 166046 -432 166102
rect -860 165922 -804 165978
rect -736 165922 -680 165978
rect -612 165922 -556 165978
rect -488 165922 -432 165978
rect -860 148294 -804 148350
rect -736 148294 -680 148350
rect -612 148294 -556 148350
rect -488 148294 -432 148350
rect -860 148170 -804 148226
rect -736 148170 -680 148226
rect -612 148170 -556 148226
rect -488 148170 -432 148226
rect -860 148046 -804 148102
rect -736 148046 -680 148102
rect -612 148046 -556 148102
rect -488 148046 -432 148102
rect -860 147922 -804 147978
rect -736 147922 -680 147978
rect -612 147922 -556 147978
rect -488 147922 -432 147978
rect -860 130294 -804 130350
rect -736 130294 -680 130350
rect -612 130294 -556 130350
rect -488 130294 -432 130350
rect -860 130170 -804 130226
rect -736 130170 -680 130226
rect -612 130170 -556 130226
rect -488 130170 -432 130226
rect -860 130046 -804 130102
rect -736 130046 -680 130102
rect -612 130046 -556 130102
rect -488 130046 -432 130102
rect -860 129922 -804 129978
rect -736 129922 -680 129978
rect -612 129922 -556 129978
rect -488 129922 -432 129978
rect -860 112294 -804 112350
rect -736 112294 -680 112350
rect -612 112294 -556 112350
rect -488 112294 -432 112350
rect -860 112170 -804 112226
rect -736 112170 -680 112226
rect -612 112170 -556 112226
rect -488 112170 -432 112226
rect -860 112046 -804 112102
rect -736 112046 -680 112102
rect -612 112046 -556 112102
rect -488 112046 -432 112102
rect -860 111922 -804 111978
rect -736 111922 -680 111978
rect -612 111922 -556 111978
rect -488 111922 -432 111978
rect -860 94294 -804 94350
rect -736 94294 -680 94350
rect -612 94294 -556 94350
rect -488 94294 -432 94350
rect -860 94170 -804 94226
rect -736 94170 -680 94226
rect -612 94170 -556 94226
rect -488 94170 -432 94226
rect -860 94046 -804 94102
rect -736 94046 -680 94102
rect -612 94046 -556 94102
rect -488 94046 -432 94102
rect -860 93922 -804 93978
rect -736 93922 -680 93978
rect -612 93922 -556 93978
rect -488 93922 -432 93978
rect -860 76294 -804 76350
rect -736 76294 -680 76350
rect -612 76294 -556 76350
rect -488 76294 -432 76350
rect -860 76170 -804 76226
rect -736 76170 -680 76226
rect -612 76170 -556 76226
rect -488 76170 -432 76226
rect -860 76046 -804 76102
rect -736 76046 -680 76102
rect -612 76046 -556 76102
rect -488 76046 -432 76102
rect -860 75922 -804 75978
rect -736 75922 -680 75978
rect -612 75922 -556 75978
rect -488 75922 -432 75978
rect -860 58294 -804 58350
rect -736 58294 -680 58350
rect -612 58294 -556 58350
rect -488 58294 -432 58350
rect -860 58170 -804 58226
rect -736 58170 -680 58226
rect -612 58170 -556 58226
rect -488 58170 -432 58226
rect -860 58046 -804 58102
rect -736 58046 -680 58102
rect -612 58046 -556 58102
rect -488 58046 -432 58102
rect -860 57922 -804 57978
rect -736 57922 -680 57978
rect -612 57922 -556 57978
rect -488 57922 -432 57978
rect -860 40294 -804 40350
rect -736 40294 -680 40350
rect -612 40294 -556 40350
rect -488 40294 -432 40350
rect -860 40170 -804 40226
rect -736 40170 -680 40226
rect -612 40170 -556 40226
rect -488 40170 -432 40226
rect -860 40046 -804 40102
rect -736 40046 -680 40102
rect -612 40046 -556 40102
rect -488 40046 -432 40102
rect -860 39922 -804 39978
rect -736 39922 -680 39978
rect -612 39922 -556 39978
rect -488 39922 -432 39978
rect -860 22294 -804 22350
rect -736 22294 -680 22350
rect -612 22294 -556 22350
rect -488 22294 -432 22350
rect -860 22170 -804 22226
rect -736 22170 -680 22226
rect -612 22170 -556 22226
rect -488 22170 -432 22226
rect -860 22046 -804 22102
rect -736 22046 -680 22102
rect -612 22046 -556 22102
rect -488 22046 -432 22102
rect -860 21922 -804 21978
rect -736 21922 -680 21978
rect -612 21922 -556 21978
rect -488 21922 -432 21978
rect 3052 79982 3108 80038
rect 5514 562294 5570 562350
rect 5638 562294 5694 562350
rect 5762 562294 5818 562350
rect 5886 562294 5942 562350
rect 5514 562170 5570 562226
rect 5638 562170 5694 562226
rect 5762 562170 5818 562226
rect 5886 562170 5942 562226
rect 5514 562046 5570 562102
rect 5638 562046 5694 562102
rect 5762 562046 5818 562102
rect 5886 562046 5942 562102
rect 5514 561922 5570 561978
rect 5638 561922 5694 561978
rect 5762 561922 5818 561978
rect 5886 561922 5942 561978
rect 5514 544294 5570 544350
rect 5638 544294 5694 544350
rect 5762 544294 5818 544350
rect 5886 544294 5942 544350
rect 5514 544170 5570 544226
rect 5638 544170 5694 544226
rect 5762 544170 5818 544226
rect 5886 544170 5942 544226
rect 5514 544046 5570 544102
rect 5638 544046 5694 544102
rect 5762 544046 5818 544102
rect 5886 544046 5942 544102
rect 5514 543922 5570 543978
rect 5638 543922 5694 543978
rect 5762 543922 5818 543978
rect 5886 543922 5942 543978
rect 5514 526294 5570 526350
rect 5638 526294 5694 526350
rect 5762 526294 5818 526350
rect 5886 526294 5942 526350
rect 5514 526170 5570 526226
rect 5638 526170 5694 526226
rect 5762 526170 5818 526226
rect 5886 526170 5942 526226
rect 5514 526046 5570 526102
rect 5638 526046 5694 526102
rect 5762 526046 5818 526102
rect 5886 526046 5942 526102
rect 5514 525922 5570 525978
rect 5638 525922 5694 525978
rect 5762 525922 5818 525978
rect 5886 525922 5942 525978
rect 5514 508294 5570 508350
rect 5638 508294 5694 508350
rect 5762 508294 5818 508350
rect 5886 508294 5942 508350
rect 5514 508170 5570 508226
rect 5638 508170 5694 508226
rect 5762 508170 5818 508226
rect 5886 508170 5942 508226
rect 5514 508046 5570 508102
rect 5638 508046 5694 508102
rect 5762 508046 5818 508102
rect 5886 508046 5942 508102
rect 5514 507922 5570 507978
rect 5638 507922 5694 507978
rect 5762 507922 5818 507978
rect 5886 507922 5942 507978
rect 5514 490294 5570 490350
rect 5638 490294 5694 490350
rect 5762 490294 5818 490350
rect 5886 490294 5942 490350
rect 5514 490170 5570 490226
rect 5638 490170 5694 490226
rect 5762 490170 5818 490226
rect 5886 490170 5942 490226
rect 5514 490046 5570 490102
rect 5638 490046 5694 490102
rect 5762 490046 5818 490102
rect 5886 490046 5942 490102
rect 5514 489922 5570 489978
rect 5638 489922 5694 489978
rect 5762 489922 5818 489978
rect 5886 489922 5942 489978
rect 9234 598116 9290 598172
rect 9358 598116 9414 598172
rect 9482 598116 9538 598172
rect 9606 598116 9662 598172
rect 9234 597992 9290 598048
rect 9358 597992 9414 598048
rect 9482 597992 9538 598048
rect 9606 597992 9662 598048
rect 9234 597868 9290 597924
rect 9358 597868 9414 597924
rect 9482 597868 9538 597924
rect 9606 597868 9662 597924
rect 9234 597744 9290 597800
rect 9358 597744 9414 597800
rect 9482 597744 9538 597800
rect 9606 597744 9662 597800
rect 36234 597156 36290 597212
rect 36358 597156 36414 597212
rect 36482 597156 36538 597212
rect 36606 597156 36662 597212
rect 36234 597032 36290 597088
rect 36358 597032 36414 597088
rect 36482 597032 36538 597088
rect 36606 597032 36662 597088
rect 36234 596908 36290 596964
rect 36358 596908 36414 596964
rect 36482 596908 36538 596964
rect 36606 596908 36662 596964
rect 36234 596784 36290 596840
rect 36358 596784 36414 596840
rect 36482 596784 36538 596840
rect 36606 596784 36662 596840
rect 9234 586294 9290 586350
rect 9358 586294 9414 586350
rect 9482 586294 9538 586350
rect 9606 586294 9662 586350
rect 9234 586170 9290 586226
rect 9358 586170 9414 586226
rect 9482 586170 9538 586226
rect 9606 586170 9662 586226
rect 9234 586046 9290 586102
rect 9358 586046 9414 586102
rect 9482 586046 9538 586102
rect 9606 586046 9662 586102
rect 9234 585922 9290 585978
rect 9358 585922 9414 585978
rect 9482 585922 9538 585978
rect 9606 585922 9662 585978
rect 9234 568294 9290 568350
rect 9358 568294 9414 568350
rect 9482 568294 9538 568350
rect 9606 568294 9662 568350
rect 9234 568170 9290 568226
rect 9358 568170 9414 568226
rect 9482 568170 9538 568226
rect 9606 568170 9662 568226
rect 9234 568046 9290 568102
rect 9358 568046 9414 568102
rect 9482 568046 9538 568102
rect 9606 568046 9662 568102
rect 9234 567922 9290 567978
rect 9358 567922 9414 567978
rect 9482 567922 9538 567978
rect 9606 567922 9662 567978
rect 9234 550294 9290 550350
rect 9358 550294 9414 550350
rect 9482 550294 9538 550350
rect 9606 550294 9662 550350
rect 9234 550170 9290 550226
rect 9358 550170 9414 550226
rect 9482 550170 9538 550226
rect 9606 550170 9662 550226
rect 9234 550046 9290 550102
rect 9358 550046 9414 550102
rect 9482 550046 9538 550102
rect 9606 550046 9662 550102
rect 9234 549922 9290 549978
rect 9358 549922 9414 549978
rect 9482 549922 9538 549978
rect 9606 549922 9662 549978
rect 9234 532294 9290 532350
rect 9358 532294 9414 532350
rect 9482 532294 9538 532350
rect 9606 532294 9662 532350
rect 9234 532170 9290 532226
rect 9358 532170 9414 532226
rect 9482 532170 9538 532226
rect 9606 532170 9662 532226
rect 9234 532046 9290 532102
rect 9358 532046 9414 532102
rect 9482 532046 9538 532102
rect 9606 532046 9662 532102
rect 9234 531922 9290 531978
rect 9358 531922 9414 531978
rect 9482 531922 9538 531978
rect 9606 531922 9662 531978
rect 9234 514294 9290 514350
rect 9358 514294 9414 514350
rect 9482 514294 9538 514350
rect 9606 514294 9662 514350
rect 9234 514170 9290 514226
rect 9358 514170 9414 514226
rect 9482 514170 9538 514226
rect 9606 514170 9662 514226
rect 9234 514046 9290 514102
rect 9358 514046 9414 514102
rect 9482 514046 9538 514102
rect 9606 514046 9662 514102
rect 9234 513922 9290 513978
rect 9358 513922 9414 513978
rect 9482 513922 9538 513978
rect 9606 513922 9662 513978
rect 9234 496294 9290 496350
rect 9358 496294 9414 496350
rect 9482 496294 9538 496350
rect 9606 496294 9662 496350
rect 9234 496170 9290 496226
rect 9358 496170 9414 496226
rect 9482 496170 9538 496226
rect 9606 496170 9662 496226
rect 9234 496046 9290 496102
rect 9358 496046 9414 496102
rect 9482 496046 9538 496102
rect 9606 496046 9662 496102
rect 9234 495922 9290 495978
rect 9358 495922 9414 495978
rect 9482 495922 9538 495978
rect 9606 495922 9662 495978
rect 5514 472294 5570 472350
rect 5638 472294 5694 472350
rect 5762 472294 5818 472350
rect 5886 472294 5942 472350
rect 5514 472170 5570 472226
rect 5638 472170 5694 472226
rect 5762 472170 5818 472226
rect 5886 472170 5942 472226
rect 5514 472046 5570 472102
rect 5638 472046 5694 472102
rect 5762 472046 5818 472102
rect 5886 472046 5942 472102
rect 5514 471922 5570 471978
rect 5638 471922 5694 471978
rect 5762 471922 5818 471978
rect 5886 471922 5942 471978
rect 5514 454294 5570 454350
rect 5638 454294 5694 454350
rect 5762 454294 5818 454350
rect 5886 454294 5942 454350
rect 5514 454170 5570 454226
rect 5638 454170 5694 454226
rect 5762 454170 5818 454226
rect 5886 454170 5942 454226
rect 5514 454046 5570 454102
rect 5638 454046 5694 454102
rect 5762 454046 5818 454102
rect 5886 454046 5942 454102
rect 5514 453922 5570 453978
rect 5638 453922 5694 453978
rect 5762 453922 5818 453978
rect 5886 453922 5942 453978
rect 5514 436294 5570 436350
rect 5638 436294 5694 436350
rect 5762 436294 5818 436350
rect 5886 436294 5942 436350
rect 5514 436170 5570 436226
rect 5638 436170 5694 436226
rect 5762 436170 5818 436226
rect 5886 436170 5942 436226
rect 5514 436046 5570 436102
rect 5638 436046 5694 436102
rect 5762 436046 5818 436102
rect 5886 436046 5942 436102
rect 5514 435922 5570 435978
rect 5638 435922 5694 435978
rect 5762 435922 5818 435978
rect 5886 435922 5942 435978
rect 5514 418294 5570 418350
rect 5638 418294 5694 418350
rect 5762 418294 5818 418350
rect 5886 418294 5942 418350
rect 5514 418170 5570 418226
rect 5638 418170 5694 418226
rect 5762 418170 5818 418226
rect 5886 418170 5942 418226
rect 5514 418046 5570 418102
rect 5638 418046 5694 418102
rect 5762 418046 5818 418102
rect 5886 418046 5942 418102
rect 5514 417922 5570 417978
rect 5638 417922 5694 417978
rect 5762 417922 5818 417978
rect 5886 417922 5942 417978
rect 5514 400294 5570 400350
rect 5638 400294 5694 400350
rect 5762 400294 5818 400350
rect 5886 400294 5942 400350
rect 5514 400170 5570 400226
rect 5638 400170 5694 400226
rect 5762 400170 5818 400226
rect 5886 400170 5942 400226
rect 5514 400046 5570 400102
rect 5638 400046 5694 400102
rect 5762 400046 5818 400102
rect 5886 400046 5942 400102
rect 5514 399922 5570 399978
rect 5638 399922 5694 399978
rect 5762 399922 5818 399978
rect 5886 399922 5942 399978
rect 5514 382294 5570 382350
rect 5638 382294 5694 382350
rect 5762 382294 5818 382350
rect 5886 382294 5942 382350
rect 5514 382170 5570 382226
rect 5638 382170 5694 382226
rect 5762 382170 5818 382226
rect 5886 382170 5942 382226
rect 5514 382046 5570 382102
rect 5638 382046 5694 382102
rect 5762 382046 5818 382102
rect 5886 382046 5942 382102
rect 5514 381922 5570 381978
rect 5638 381922 5694 381978
rect 5762 381922 5818 381978
rect 5886 381922 5942 381978
rect 5514 364294 5570 364350
rect 5638 364294 5694 364350
rect 5762 364294 5818 364350
rect 5886 364294 5942 364350
rect 5514 364170 5570 364226
rect 5638 364170 5694 364226
rect 5762 364170 5818 364226
rect 5886 364170 5942 364226
rect 5514 364046 5570 364102
rect 5638 364046 5694 364102
rect 5762 364046 5818 364102
rect 5886 364046 5942 364102
rect 5514 363922 5570 363978
rect 5638 363922 5694 363978
rect 5762 363922 5818 363978
rect 5886 363922 5942 363978
rect 5514 346294 5570 346350
rect 5638 346294 5694 346350
rect 5762 346294 5818 346350
rect 5886 346294 5942 346350
rect 5514 346170 5570 346226
rect 5638 346170 5694 346226
rect 5762 346170 5818 346226
rect 5886 346170 5942 346226
rect 5514 346046 5570 346102
rect 5638 346046 5694 346102
rect 5762 346046 5818 346102
rect 5886 346046 5942 346102
rect 5514 345922 5570 345978
rect 5638 345922 5694 345978
rect 5762 345922 5818 345978
rect 5886 345922 5942 345978
rect 5514 328294 5570 328350
rect 5638 328294 5694 328350
rect 5762 328294 5818 328350
rect 5886 328294 5942 328350
rect 5514 328170 5570 328226
rect 5638 328170 5694 328226
rect 5762 328170 5818 328226
rect 5886 328170 5942 328226
rect 5514 328046 5570 328102
rect 5638 328046 5694 328102
rect 5762 328046 5818 328102
rect 5886 328046 5942 328102
rect 5514 327922 5570 327978
rect 5638 327922 5694 327978
rect 5762 327922 5818 327978
rect 5886 327922 5942 327978
rect 5514 310294 5570 310350
rect 5638 310294 5694 310350
rect 5762 310294 5818 310350
rect 5886 310294 5942 310350
rect 5514 310170 5570 310226
rect 5638 310170 5694 310226
rect 5762 310170 5818 310226
rect 5886 310170 5942 310226
rect 5514 310046 5570 310102
rect 5638 310046 5694 310102
rect 5762 310046 5818 310102
rect 5886 310046 5942 310102
rect 5514 309922 5570 309978
rect 5638 309922 5694 309978
rect 5762 309922 5818 309978
rect 5886 309922 5942 309978
rect 5514 292294 5570 292350
rect 5638 292294 5694 292350
rect 5762 292294 5818 292350
rect 5886 292294 5942 292350
rect 5514 292170 5570 292226
rect 5638 292170 5694 292226
rect 5762 292170 5818 292226
rect 5886 292170 5942 292226
rect 5514 292046 5570 292102
rect 5638 292046 5694 292102
rect 5762 292046 5818 292102
rect 5886 292046 5942 292102
rect 5514 291922 5570 291978
rect 5638 291922 5694 291978
rect 5762 291922 5818 291978
rect 5886 291922 5942 291978
rect 5514 274294 5570 274350
rect 5638 274294 5694 274350
rect 5762 274294 5818 274350
rect 5886 274294 5942 274350
rect 5514 274170 5570 274226
rect 5638 274170 5694 274226
rect 5762 274170 5818 274226
rect 5886 274170 5942 274226
rect 5514 274046 5570 274102
rect 5638 274046 5694 274102
rect 5762 274046 5818 274102
rect 5886 274046 5942 274102
rect 5514 273922 5570 273978
rect 5638 273922 5694 273978
rect 5762 273922 5818 273978
rect 5886 273922 5942 273978
rect 5514 256294 5570 256350
rect 5638 256294 5694 256350
rect 5762 256294 5818 256350
rect 5886 256294 5942 256350
rect 5514 256170 5570 256226
rect 5638 256170 5694 256226
rect 5762 256170 5818 256226
rect 5886 256170 5942 256226
rect 5514 256046 5570 256102
rect 5638 256046 5694 256102
rect 5762 256046 5818 256102
rect 5886 256046 5942 256102
rect 5514 255922 5570 255978
rect 5638 255922 5694 255978
rect 5762 255922 5818 255978
rect 5886 255922 5942 255978
rect 5514 238294 5570 238350
rect 5638 238294 5694 238350
rect 5762 238294 5818 238350
rect 5886 238294 5942 238350
rect 5514 238170 5570 238226
rect 5638 238170 5694 238226
rect 5762 238170 5818 238226
rect 5886 238170 5942 238226
rect 5514 238046 5570 238102
rect 5638 238046 5694 238102
rect 5762 238046 5818 238102
rect 5886 238046 5942 238102
rect 5514 237922 5570 237978
rect 5638 237922 5694 237978
rect 5762 237922 5818 237978
rect 5886 237922 5942 237978
rect 5514 220294 5570 220350
rect 5638 220294 5694 220350
rect 5762 220294 5818 220350
rect 5886 220294 5942 220350
rect 5514 220170 5570 220226
rect 5638 220170 5694 220226
rect 5762 220170 5818 220226
rect 5886 220170 5942 220226
rect 5514 220046 5570 220102
rect 5638 220046 5694 220102
rect 5762 220046 5818 220102
rect 5886 220046 5942 220102
rect 5514 219922 5570 219978
rect 5638 219922 5694 219978
rect 5762 219922 5818 219978
rect 5886 219922 5942 219978
rect 5514 202294 5570 202350
rect 5638 202294 5694 202350
rect 5762 202294 5818 202350
rect 5886 202294 5942 202350
rect 5514 202170 5570 202226
rect 5638 202170 5694 202226
rect 5762 202170 5818 202226
rect 5886 202170 5942 202226
rect 5514 202046 5570 202102
rect 5638 202046 5694 202102
rect 5762 202046 5818 202102
rect 5886 202046 5942 202102
rect 5514 201922 5570 201978
rect 5638 201922 5694 201978
rect 5762 201922 5818 201978
rect 5886 201922 5942 201978
rect 5514 184294 5570 184350
rect 5638 184294 5694 184350
rect 5762 184294 5818 184350
rect 5886 184294 5942 184350
rect 5514 184170 5570 184226
rect 5638 184170 5694 184226
rect 5762 184170 5818 184226
rect 5886 184170 5942 184226
rect 5514 184046 5570 184102
rect 5638 184046 5694 184102
rect 5762 184046 5818 184102
rect 5886 184046 5942 184102
rect 5514 183922 5570 183978
rect 5638 183922 5694 183978
rect 5762 183922 5818 183978
rect 5886 183922 5942 183978
rect 5514 166294 5570 166350
rect 5638 166294 5694 166350
rect 5762 166294 5818 166350
rect 5886 166294 5942 166350
rect 5514 166170 5570 166226
rect 5638 166170 5694 166226
rect 5762 166170 5818 166226
rect 5886 166170 5942 166226
rect 5514 166046 5570 166102
rect 5638 166046 5694 166102
rect 5762 166046 5818 166102
rect 5886 166046 5942 166102
rect 5514 165922 5570 165978
rect 5638 165922 5694 165978
rect 5762 165922 5818 165978
rect 5886 165922 5942 165978
rect 5514 148294 5570 148350
rect 5638 148294 5694 148350
rect 5762 148294 5818 148350
rect 5886 148294 5942 148350
rect 5514 148170 5570 148226
rect 5638 148170 5694 148226
rect 5762 148170 5818 148226
rect 5886 148170 5942 148226
rect 5514 148046 5570 148102
rect 5638 148046 5694 148102
rect 5762 148046 5818 148102
rect 5886 148046 5942 148102
rect 5514 147922 5570 147978
rect 5638 147922 5694 147978
rect 5762 147922 5818 147978
rect 5886 147922 5942 147978
rect 5514 130294 5570 130350
rect 5638 130294 5694 130350
rect 5762 130294 5818 130350
rect 5886 130294 5942 130350
rect 5514 130170 5570 130226
rect 5638 130170 5694 130226
rect 5762 130170 5818 130226
rect 5886 130170 5942 130226
rect 5514 130046 5570 130102
rect 5638 130046 5694 130102
rect 5762 130046 5818 130102
rect 5886 130046 5942 130102
rect 5514 129922 5570 129978
rect 5638 129922 5694 129978
rect 5762 129922 5818 129978
rect 5886 129922 5942 129978
rect 5514 112294 5570 112350
rect 5638 112294 5694 112350
rect 5762 112294 5818 112350
rect 5886 112294 5942 112350
rect 5514 112170 5570 112226
rect 5638 112170 5694 112226
rect 5762 112170 5818 112226
rect 5886 112170 5942 112226
rect 5514 112046 5570 112102
rect 5638 112046 5694 112102
rect 5762 112046 5818 112102
rect 5886 112046 5942 112102
rect 5514 111922 5570 111978
rect 5638 111922 5694 111978
rect 5762 111922 5818 111978
rect 5886 111922 5942 111978
rect 5514 94294 5570 94350
rect 5638 94294 5694 94350
rect 5762 94294 5818 94350
rect 5886 94294 5942 94350
rect 5514 94170 5570 94226
rect 5638 94170 5694 94226
rect 5762 94170 5818 94226
rect 5886 94170 5942 94226
rect 5514 94046 5570 94102
rect 5638 94046 5694 94102
rect 5762 94046 5818 94102
rect 5886 94046 5942 94102
rect 5514 93922 5570 93978
rect 5638 93922 5694 93978
rect 5762 93922 5818 93978
rect 5886 93922 5942 93978
rect 5514 76294 5570 76350
rect 5638 76294 5694 76350
rect 5762 76294 5818 76350
rect 5886 76294 5942 76350
rect 5514 76170 5570 76226
rect 5638 76170 5694 76226
rect 5762 76170 5818 76226
rect 5886 76170 5942 76226
rect 5514 76046 5570 76102
rect 5638 76046 5694 76102
rect 5762 76046 5818 76102
rect 5886 76046 5942 76102
rect 5514 75922 5570 75978
rect 5638 75922 5694 75978
rect 5762 75922 5818 75978
rect 5886 75922 5942 75978
rect 5514 58294 5570 58350
rect 5638 58294 5694 58350
rect 5762 58294 5818 58350
rect 5886 58294 5942 58350
rect 5514 58170 5570 58226
rect 5638 58170 5694 58226
rect 5762 58170 5818 58226
rect 5886 58170 5942 58226
rect 5514 58046 5570 58102
rect 5638 58046 5694 58102
rect 5762 58046 5818 58102
rect 5886 58046 5942 58102
rect 5514 57922 5570 57978
rect 5638 57922 5694 57978
rect 5762 57922 5818 57978
rect 5886 57922 5942 57978
rect 5514 40294 5570 40350
rect 5638 40294 5694 40350
rect 5762 40294 5818 40350
rect 5886 40294 5942 40350
rect 5514 40170 5570 40226
rect 5638 40170 5694 40226
rect 5762 40170 5818 40226
rect 5886 40170 5942 40226
rect 5514 40046 5570 40102
rect 5638 40046 5694 40102
rect 5762 40046 5818 40102
rect 5886 40046 5942 40102
rect 5514 39922 5570 39978
rect 5638 39922 5694 39978
rect 5762 39922 5818 39978
rect 5886 39922 5942 39978
rect 5514 22294 5570 22350
rect 5638 22294 5694 22350
rect 5762 22294 5818 22350
rect 5886 22294 5942 22350
rect 5514 22170 5570 22226
rect 5638 22170 5694 22226
rect 5762 22170 5818 22226
rect 5886 22170 5942 22226
rect 5514 22046 5570 22102
rect 5638 22046 5694 22102
rect 5762 22046 5818 22102
rect 5886 22046 5942 22102
rect 5514 21922 5570 21978
rect 5638 21922 5694 21978
rect 5762 21922 5818 21978
rect 5886 21922 5942 21978
rect -860 4294 -804 4350
rect -736 4294 -680 4350
rect -612 4294 -556 4350
rect -488 4294 -432 4350
rect -860 4170 -804 4226
rect -736 4170 -680 4226
rect -612 4170 -556 4226
rect -488 4170 -432 4226
rect -860 4046 -804 4102
rect -736 4046 -680 4102
rect -612 4046 -556 4102
rect -488 4046 -432 4102
rect -860 3922 -804 3978
rect -736 3922 -680 3978
rect -612 3922 -556 3978
rect -488 3922 -432 3978
rect -860 -216 -804 -160
rect -736 -216 -680 -160
rect -612 -216 -556 -160
rect -488 -216 -432 -160
rect -860 -340 -804 -284
rect -736 -340 -680 -284
rect -612 -340 -556 -284
rect -488 -340 -432 -284
rect -860 -464 -804 -408
rect -736 -464 -680 -408
rect -612 -464 -556 -408
rect -488 -464 -432 -408
rect -860 -588 -804 -532
rect -736 -588 -680 -532
rect -612 -588 -556 -532
rect -488 -588 -432 -532
rect 6524 79802 6580 79858
rect 6636 78182 6692 78238
rect 8092 78362 8148 78418
rect 7980 74942 8036 74998
rect 9234 478294 9290 478350
rect 9358 478294 9414 478350
rect 9482 478294 9538 478350
rect 9606 478294 9662 478350
rect 9234 478170 9290 478226
rect 9358 478170 9414 478226
rect 9482 478170 9538 478226
rect 9606 478170 9662 478226
rect 9234 478046 9290 478102
rect 9358 478046 9414 478102
rect 9482 478046 9538 478102
rect 9606 478046 9662 478102
rect 9234 477922 9290 477978
rect 9358 477922 9414 477978
rect 9482 477922 9538 477978
rect 9606 477922 9662 477978
rect 9234 460294 9290 460350
rect 9358 460294 9414 460350
rect 9482 460294 9538 460350
rect 9606 460294 9662 460350
rect 9234 460170 9290 460226
rect 9358 460170 9414 460226
rect 9482 460170 9538 460226
rect 9606 460170 9662 460226
rect 9234 460046 9290 460102
rect 9358 460046 9414 460102
rect 9482 460046 9538 460102
rect 9606 460046 9662 460102
rect 9234 459922 9290 459978
rect 9358 459922 9414 459978
rect 9482 459922 9538 459978
rect 9606 459922 9662 459978
rect 9234 442294 9290 442350
rect 9358 442294 9414 442350
rect 9482 442294 9538 442350
rect 9606 442294 9662 442350
rect 9234 442170 9290 442226
rect 9358 442170 9414 442226
rect 9482 442170 9538 442226
rect 9606 442170 9662 442226
rect 9234 442046 9290 442102
rect 9358 442046 9414 442102
rect 9482 442046 9538 442102
rect 9606 442046 9662 442102
rect 9234 441922 9290 441978
rect 9358 441922 9414 441978
rect 9482 441922 9538 441978
rect 9606 441922 9662 441978
rect 9234 424294 9290 424350
rect 9358 424294 9414 424350
rect 9482 424294 9538 424350
rect 9606 424294 9662 424350
rect 9234 424170 9290 424226
rect 9358 424170 9414 424226
rect 9482 424170 9538 424226
rect 9606 424170 9662 424226
rect 9234 424046 9290 424102
rect 9358 424046 9414 424102
rect 9482 424046 9538 424102
rect 9606 424046 9662 424102
rect 9234 423922 9290 423978
rect 9358 423922 9414 423978
rect 9482 423922 9538 423978
rect 9606 423922 9662 423978
rect 9234 406294 9290 406350
rect 9358 406294 9414 406350
rect 9482 406294 9538 406350
rect 9606 406294 9662 406350
rect 9234 406170 9290 406226
rect 9358 406170 9414 406226
rect 9482 406170 9538 406226
rect 9606 406170 9662 406226
rect 9234 406046 9290 406102
rect 9358 406046 9414 406102
rect 9482 406046 9538 406102
rect 9606 406046 9662 406102
rect 9234 405922 9290 405978
rect 9358 405922 9414 405978
rect 9482 405922 9538 405978
rect 9606 405922 9662 405978
rect 9234 388294 9290 388350
rect 9358 388294 9414 388350
rect 9482 388294 9538 388350
rect 9606 388294 9662 388350
rect 9234 388170 9290 388226
rect 9358 388170 9414 388226
rect 9482 388170 9538 388226
rect 9606 388170 9662 388226
rect 9234 388046 9290 388102
rect 9358 388046 9414 388102
rect 9482 388046 9538 388102
rect 9606 388046 9662 388102
rect 9234 387922 9290 387978
rect 9358 387922 9414 387978
rect 9482 387922 9538 387978
rect 9606 387922 9662 387978
rect 9234 370294 9290 370350
rect 9358 370294 9414 370350
rect 9482 370294 9538 370350
rect 9606 370294 9662 370350
rect 9234 370170 9290 370226
rect 9358 370170 9414 370226
rect 9482 370170 9538 370226
rect 9606 370170 9662 370226
rect 9234 370046 9290 370102
rect 9358 370046 9414 370102
rect 9482 370046 9538 370102
rect 9606 370046 9662 370102
rect 9234 369922 9290 369978
rect 9358 369922 9414 369978
rect 9482 369922 9538 369978
rect 9606 369922 9662 369978
rect 9234 352294 9290 352350
rect 9358 352294 9414 352350
rect 9482 352294 9538 352350
rect 9606 352294 9662 352350
rect 9234 352170 9290 352226
rect 9358 352170 9414 352226
rect 9482 352170 9538 352226
rect 9606 352170 9662 352226
rect 9234 352046 9290 352102
rect 9358 352046 9414 352102
rect 9482 352046 9538 352102
rect 9606 352046 9662 352102
rect 9234 351922 9290 351978
rect 9358 351922 9414 351978
rect 9482 351922 9538 351978
rect 9606 351922 9662 351978
rect 9234 334294 9290 334350
rect 9358 334294 9414 334350
rect 9482 334294 9538 334350
rect 9606 334294 9662 334350
rect 9234 334170 9290 334226
rect 9358 334170 9414 334226
rect 9482 334170 9538 334226
rect 9606 334170 9662 334226
rect 9234 334046 9290 334102
rect 9358 334046 9414 334102
rect 9482 334046 9538 334102
rect 9606 334046 9662 334102
rect 9234 333922 9290 333978
rect 9358 333922 9414 333978
rect 9482 333922 9538 333978
rect 9606 333922 9662 333978
rect 9234 316294 9290 316350
rect 9358 316294 9414 316350
rect 9482 316294 9538 316350
rect 9606 316294 9662 316350
rect 9234 316170 9290 316226
rect 9358 316170 9414 316226
rect 9482 316170 9538 316226
rect 9606 316170 9662 316226
rect 9234 316046 9290 316102
rect 9358 316046 9414 316102
rect 9482 316046 9538 316102
rect 9606 316046 9662 316102
rect 9234 315922 9290 315978
rect 9358 315922 9414 315978
rect 9482 315922 9538 315978
rect 9606 315922 9662 315978
rect 9234 298294 9290 298350
rect 9358 298294 9414 298350
rect 9482 298294 9538 298350
rect 9606 298294 9662 298350
rect 9234 298170 9290 298226
rect 9358 298170 9414 298226
rect 9482 298170 9538 298226
rect 9606 298170 9662 298226
rect 9234 298046 9290 298102
rect 9358 298046 9414 298102
rect 9482 298046 9538 298102
rect 9606 298046 9662 298102
rect 9234 297922 9290 297978
rect 9358 297922 9414 297978
rect 9482 297922 9538 297978
rect 9606 297922 9662 297978
rect 9234 280294 9290 280350
rect 9358 280294 9414 280350
rect 9482 280294 9538 280350
rect 9606 280294 9662 280350
rect 9234 280170 9290 280226
rect 9358 280170 9414 280226
rect 9482 280170 9538 280226
rect 9606 280170 9662 280226
rect 9234 280046 9290 280102
rect 9358 280046 9414 280102
rect 9482 280046 9538 280102
rect 9606 280046 9662 280102
rect 9234 279922 9290 279978
rect 9358 279922 9414 279978
rect 9482 279922 9538 279978
rect 9606 279922 9662 279978
rect 9234 262294 9290 262350
rect 9358 262294 9414 262350
rect 9482 262294 9538 262350
rect 9606 262294 9662 262350
rect 9234 262170 9290 262226
rect 9358 262170 9414 262226
rect 9482 262170 9538 262226
rect 9606 262170 9662 262226
rect 9234 262046 9290 262102
rect 9358 262046 9414 262102
rect 9482 262046 9538 262102
rect 9606 262046 9662 262102
rect 9234 261922 9290 261978
rect 9358 261922 9414 261978
rect 9482 261922 9538 261978
rect 9606 261922 9662 261978
rect 9234 244294 9290 244350
rect 9358 244294 9414 244350
rect 9482 244294 9538 244350
rect 9606 244294 9662 244350
rect 9234 244170 9290 244226
rect 9358 244170 9414 244226
rect 9482 244170 9538 244226
rect 9606 244170 9662 244226
rect 9234 244046 9290 244102
rect 9358 244046 9414 244102
rect 9482 244046 9538 244102
rect 9606 244046 9662 244102
rect 9234 243922 9290 243978
rect 9358 243922 9414 243978
rect 9482 243922 9538 243978
rect 9606 243922 9662 243978
rect 9234 226294 9290 226350
rect 9358 226294 9414 226350
rect 9482 226294 9538 226350
rect 9606 226294 9662 226350
rect 9234 226170 9290 226226
rect 9358 226170 9414 226226
rect 9482 226170 9538 226226
rect 9606 226170 9662 226226
rect 9234 226046 9290 226102
rect 9358 226046 9414 226102
rect 9482 226046 9538 226102
rect 9606 226046 9662 226102
rect 9234 225922 9290 225978
rect 9358 225922 9414 225978
rect 9482 225922 9538 225978
rect 9606 225922 9662 225978
rect 9234 208294 9290 208350
rect 9358 208294 9414 208350
rect 9482 208294 9538 208350
rect 9606 208294 9662 208350
rect 9234 208170 9290 208226
rect 9358 208170 9414 208226
rect 9482 208170 9538 208226
rect 9606 208170 9662 208226
rect 9234 208046 9290 208102
rect 9358 208046 9414 208102
rect 9482 208046 9538 208102
rect 9606 208046 9662 208102
rect 9234 207922 9290 207978
rect 9358 207922 9414 207978
rect 9482 207922 9538 207978
rect 9606 207922 9662 207978
rect 9234 190294 9290 190350
rect 9358 190294 9414 190350
rect 9482 190294 9538 190350
rect 9606 190294 9662 190350
rect 9234 190170 9290 190226
rect 9358 190170 9414 190226
rect 9482 190170 9538 190226
rect 9606 190170 9662 190226
rect 9234 190046 9290 190102
rect 9358 190046 9414 190102
rect 9482 190046 9538 190102
rect 9606 190046 9662 190102
rect 9234 189922 9290 189978
rect 9358 189922 9414 189978
rect 9482 189922 9538 189978
rect 9606 189922 9662 189978
rect 9234 172294 9290 172350
rect 9358 172294 9414 172350
rect 9482 172294 9538 172350
rect 9606 172294 9662 172350
rect 9234 172170 9290 172226
rect 9358 172170 9414 172226
rect 9482 172170 9538 172226
rect 9606 172170 9662 172226
rect 9234 172046 9290 172102
rect 9358 172046 9414 172102
rect 9482 172046 9538 172102
rect 9606 172046 9662 172102
rect 9234 171922 9290 171978
rect 9358 171922 9414 171978
rect 9482 171922 9538 171978
rect 9606 171922 9662 171978
rect 9234 154294 9290 154350
rect 9358 154294 9414 154350
rect 9482 154294 9538 154350
rect 9606 154294 9662 154350
rect 9234 154170 9290 154226
rect 9358 154170 9414 154226
rect 9482 154170 9538 154226
rect 9606 154170 9662 154226
rect 9234 154046 9290 154102
rect 9358 154046 9414 154102
rect 9482 154046 9538 154102
rect 9606 154046 9662 154102
rect 9234 153922 9290 153978
rect 9358 153922 9414 153978
rect 9482 153922 9538 153978
rect 9606 153922 9662 153978
rect 9234 136294 9290 136350
rect 9358 136294 9414 136350
rect 9482 136294 9538 136350
rect 9606 136294 9662 136350
rect 9234 136170 9290 136226
rect 9358 136170 9414 136226
rect 9482 136170 9538 136226
rect 9606 136170 9662 136226
rect 9234 136046 9290 136102
rect 9358 136046 9414 136102
rect 9482 136046 9538 136102
rect 9606 136046 9662 136102
rect 9234 135922 9290 135978
rect 9358 135922 9414 135978
rect 9482 135922 9538 135978
rect 9606 135922 9662 135978
rect 9234 118294 9290 118350
rect 9358 118294 9414 118350
rect 9482 118294 9538 118350
rect 9606 118294 9662 118350
rect 9234 118170 9290 118226
rect 9358 118170 9414 118226
rect 9482 118170 9538 118226
rect 9606 118170 9662 118226
rect 9234 118046 9290 118102
rect 9358 118046 9414 118102
rect 9482 118046 9538 118102
rect 9606 118046 9662 118102
rect 9234 117922 9290 117978
rect 9358 117922 9414 117978
rect 9482 117922 9538 117978
rect 9606 117922 9662 117978
rect 9234 100294 9290 100350
rect 9358 100294 9414 100350
rect 9482 100294 9538 100350
rect 9606 100294 9662 100350
rect 9234 100170 9290 100226
rect 9358 100170 9414 100226
rect 9482 100170 9538 100226
rect 9606 100170 9662 100226
rect 9234 100046 9290 100102
rect 9358 100046 9414 100102
rect 9482 100046 9538 100102
rect 9606 100046 9662 100102
rect 9234 99922 9290 99978
rect 9358 99922 9414 99978
rect 9482 99922 9538 99978
rect 9606 99922 9662 99978
rect 9234 82294 9290 82350
rect 9358 82294 9414 82350
rect 9482 82294 9538 82350
rect 9606 82294 9662 82350
rect 9234 82170 9290 82226
rect 9358 82170 9414 82226
rect 9482 82170 9538 82226
rect 9606 82170 9662 82226
rect 9234 82046 9290 82102
rect 9358 82046 9414 82102
rect 9482 82046 9538 82102
rect 9606 82046 9662 82102
rect 9234 81922 9290 81978
rect 9358 81922 9414 81978
rect 9482 81922 9538 81978
rect 9606 81922 9662 81978
rect 8988 72062 9044 72118
rect 8876 68822 8932 68878
rect 9234 64294 9290 64350
rect 9358 64294 9414 64350
rect 9482 64294 9538 64350
rect 9606 64294 9662 64350
rect 9234 64170 9290 64226
rect 9358 64170 9414 64226
rect 9482 64170 9538 64226
rect 9606 64170 9662 64226
rect 9234 64046 9290 64102
rect 9358 64046 9414 64102
rect 9482 64046 9538 64102
rect 9606 64046 9662 64102
rect 9234 63922 9290 63978
rect 9358 63922 9414 63978
rect 9482 63922 9538 63978
rect 9606 63922 9662 63978
rect 9234 46294 9290 46350
rect 9358 46294 9414 46350
rect 9482 46294 9538 46350
rect 9606 46294 9662 46350
rect 9234 46170 9290 46226
rect 9358 46170 9414 46226
rect 9482 46170 9538 46226
rect 9606 46170 9662 46226
rect 9234 46046 9290 46102
rect 9358 46046 9414 46102
rect 9482 46046 9538 46102
rect 9606 46046 9662 46102
rect 9234 45922 9290 45978
rect 9358 45922 9414 45978
rect 9482 45922 9538 45978
rect 9606 45922 9662 45978
rect 9996 49562 10052 49618
rect 9234 28294 9290 28350
rect 9358 28294 9414 28350
rect 9482 28294 9538 28350
rect 9606 28294 9662 28350
rect 9234 28170 9290 28226
rect 9358 28170 9414 28226
rect 9482 28170 9538 28226
rect 9606 28170 9662 28226
rect 9234 28046 9290 28102
rect 9358 28046 9414 28102
rect 9482 28046 9538 28102
rect 9606 28046 9662 28102
rect 9234 27922 9290 27978
rect 9358 27922 9414 27978
rect 9482 27922 9538 27978
rect 9606 27922 9662 27978
rect 11452 78002 11508 78058
rect 11564 74762 11620 74818
rect 12684 69002 12740 69058
rect 13468 68822 13524 68878
rect 12684 67022 12740 67078
rect 12460 65402 12516 65458
rect 12460 63602 12516 63658
rect 12684 61982 12740 62038
rect 12684 60722 12740 60778
rect 12460 60362 12516 60418
rect 15148 72062 15204 72118
rect 15932 69002 15988 69058
rect 14252 60722 14308 60778
rect 16518 58294 16574 58350
rect 16642 58294 16698 58350
rect 16518 58170 16574 58226
rect 16642 58170 16698 58226
rect 16518 58046 16574 58102
rect 16642 58046 16698 58102
rect 16518 57922 16574 57978
rect 16642 57922 16698 57978
rect 12348 56942 12404 56998
rect 12348 54602 12404 54658
rect 12684 53732 12740 53758
rect 12684 53702 12740 53732
rect 17612 53702 17668 53758
rect 12348 51902 12404 51958
rect 12684 48662 12740 48718
rect 20972 61982 21028 62038
rect 24332 56942 24388 56998
rect 26012 54602 26068 54658
rect 22652 51902 22708 51958
rect 36234 580294 36290 580350
rect 36358 580294 36414 580350
rect 36482 580294 36538 580350
rect 36606 580294 36662 580350
rect 36234 580170 36290 580226
rect 36358 580170 36414 580226
rect 36482 580170 36538 580226
rect 36606 580170 36662 580226
rect 36234 580046 36290 580102
rect 36358 580046 36414 580102
rect 36482 580046 36538 580102
rect 36606 580046 36662 580102
rect 36234 579922 36290 579978
rect 36358 579922 36414 579978
rect 36482 579922 36538 579978
rect 36606 579922 36662 579978
rect 36234 562294 36290 562350
rect 36358 562294 36414 562350
rect 36482 562294 36538 562350
rect 36606 562294 36662 562350
rect 36234 562170 36290 562226
rect 36358 562170 36414 562226
rect 36482 562170 36538 562226
rect 36606 562170 36662 562226
rect 36234 562046 36290 562102
rect 36358 562046 36414 562102
rect 36482 562046 36538 562102
rect 36606 562046 36662 562102
rect 36234 561922 36290 561978
rect 36358 561922 36414 561978
rect 36482 561922 36538 561978
rect 36606 561922 36662 561978
rect 36234 544294 36290 544350
rect 36358 544294 36414 544350
rect 36482 544294 36538 544350
rect 36606 544294 36662 544350
rect 36234 544170 36290 544226
rect 36358 544170 36414 544226
rect 36482 544170 36538 544226
rect 36606 544170 36662 544226
rect 36234 544046 36290 544102
rect 36358 544046 36414 544102
rect 36482 544046 36538 544102
rect 36606 544046 36662 544102
rect 36234 543922 36290 543978
rect 36358 543922 36414 543978
rect 36482 543922 36538 543978
rect 36606 543922 36662 543978
rect 36234 526294 36290 526350
rect 36358 526294 36414 526350
rect 36482 526294 36538 526350
rect 36606 526294 36662 526350
rect 36234 526170 36290 526226
rect 36358 526170 36414 526226
rect 36482 526170 36538 526226
rect 36606 526170 36662 526226
rect 36234 526046 36290 526102
rect 36358 526046 36414 526102
rect 36482 526046 36538 526102
rect 36606 526046 36662 526102
rect 36234 525922 36290 525978
rect 36358 525922 36414 525978
rect 36482 525922 36538 525978
rect 36606 525922 36662 525978
rect 36234 508294 36290 508350
rect 36358 508294 36414 508350
rect 36482 508294 36538 508350
rect 36606 508294 36662 508350
rect 36234 508170 36290 508226
rect 36358 508170 36414 508226
rect 36482 508170 36538 508226
rect 36606 508170 36662 508226
rect 36234 508046 36290 508102
rect 36358 508046 36414 508102
rect 36482 508046 36538 508102
rect 36606 508046 36662 508102
rect 36234 507922 36290 507978
rect 36358 507922 36414 507978
rect 36482 507922 36538 507978
rect 36606 507922 36662 507978
rect 29372 67022 29428 67078
rect 36234 490294 36290 490350
rect 36358 490294 36414 490350
rect 36482 490294 36538 490350
rect 36606 490294 36662 490350
rect 36234 490170 36290 490226
rect 36358 490170 36414 490226
rect 36482 490170 36538 490226
rect 36606 490170 36662 490226
rect 36234 490046 36290 490102
rect 36358 490046 36414 490102
rect 36482 490046 36538 490102
rect 36606 490046 36662 490102
rect 36234 489922 36290 489978
rect 36358 489922 36414 489978
rect 36482 489922 36538 489978
rect 36606 489922 36662 489978
rect 36234 472294 36290 472350
rect 36358 472294 36414 472350
rect 36482 472294 36538 472350
rect 36606 472294 36662 472350
rect 36234 472170 36290 472226
rect 36358 472170 36414 472226
rect 36482 472170 36538 472226
rect 36606 472170 36662 472226
rect 36234 472046 36290 472102
rect 36358 472046 36414 472102
rect 36482 472046 36538 472102
rect 36606 472046 36662 472102
rect 36234 471922 36290 471978
rect 36358 471922 36414 471978
rect 36482 471922 36538 471978
rect 36606 471922 36662 471978
rect 36234 454294 36290 454350
rect 36358 454294 36414 454350
rect 36482 454294 36538 454350
rect 36606 454294 36662 454350
rect 36234 454170 36290 454226
rect 36358 454170 36414 454226
rect 36482 454170 36538 454226
rect 36606 454170 36662 454226
rect 36234 454046 36290 454102
rect 36358 454046 36414 454102
rect 36482 454046 36538 454102
rect 36606 454046 36662 454102
rect 36234 453922 36290 453978
rect 36358 453922 36414 453978
rect 36482 453922 36538 453978
rect 36606 453922 36662 453978
rect 36234 436294 36290 436350
rect 36358 436294 36414 436350
rect 36482 436294 36538 436350
rect 36606 436294 36662 436350
rect 36234 436170 36290 436226
rect 36358 436170 36414 436226
rect 36482 436170 36538 436226
rect 36606 436170 36662 436226
rect 36234 436046 36290 436102
rect 36358 436046 36414 436102
rect 36482 436046 36538 436102
rect 36606 436046 36662 436102
rect 36234 435922 36290 435978
rect 36358 435922 36414 435978
rect 36482 435922 36538 435978
rect 36606 435922 36662 435978
rect 36234 418294 36290 418350
rect 36358 418294 36414 418350
rect 36482 418294 36538 418350
rect 36606 418294 36662 418350
rect 36234 418170 36290 418226
rect 36358 418170 36414 418226
rect 36482 418170 36538 418226
rect 36606 418170 36662 418226
rect 36234 418046 36290 418102
rect 36358 418046 36414 418102
rect 36482 418046 36538 418102
rect 36606 418046 36662 418102
rect 36234 417922 36290 417978
rect 36358 417922 36414 417978
rect 36482 417922 36538 417978
rect 36606 417922 36662 417978
rect 36234 400294 36290 400350
rect 36358 400294 36414 400350
rect 36482 400294 36538 400350
rect 36606 400294 36662 400350
rect 36234 400170 36290 400226
rect 36358 400170 36414 400226
rect 36482 400170 36538 400226
rect 36606 400170 36662 400226
rect 36234 400046 36290 400102
rect 36358 400046 36414 400102
rect 36482 400046 36538 400102
rect 36606 400046 36662 400102
rect 36234 399922 36290 399978
rect 36358 399922 36414 399978
rect 36482 399922 36538 399978
rect 36606 399922 36662 399978
rect 36234 382294 36290 382350
rect 36358 382294 36414 382350
rect 36482 382294 36538 382350
rect 36606 382294 36662 382350
rect 36234 382170 36290 382226
rect 36358 382170 36414 382226
rect 36482 382170 36538 382226
rect 36606 382170 36662 382226
rect 36234 382046 36290 382102
rect 36358 382046 36414 382102
rect 36482 382046 36538 382102
rect 36606 382046 36662 382102
rect 36234 381922 36290 381978
rect 36358 381922 36414 381978
rect 36482 381922 36538 381978
rect 36606 381922 36662 381978
rect 36234 364294 36290 364350
rect 36358 364294 36414 364350
rect 36482 364294 36538 364350
rect 36606 364294 36662 364350
rect 36234 364170 36290 364226
rect 36358 364170 36414 364226
rect 36482 364170 36538 364226
rect 36606 364170 36662 364226
rect 36234 364046 36290 364102
rect 36358 364046 36414 364102
rect 36482 364046 36538 364102
rect 36606 364046 36662 364102
rect 36234 363922 36290 363978
rect 36358 363922 36414 363978
rect 36482 363922 36538 363978
rect 36606 363922 36662 363978
rect 36234 346294 36290 346350
rect 36358 346294 36414 346350
rect 36482 346294 36538 346350
rect 36606 346294 36662 346350
rect 36234 346170 36290 346226
rect 36358 346170 36414 346226
rect 36482 346170 36538 346226
rect 36606 346170 36662 346226
rect 36234 346046 36290 346102
rect 36358 346046 36414 346102
rect 36482 346046 36538 346102
rect 36606 346046 36662 346102
rect 36234 345922 36290 345978
rect 36358 345922 36414 345978
rect 36482 345922 36538 345978
rect 36606 345922 36662 345978
rect 36234 328294 36290 328350
rect 36358 328294 36414 328350
rect 36482 328294 36538 328350
rect 36606 328294 36662 328350
rect 36234 328170 36290 328226
rect 36358 328170 36414 328226
rect 36482 328170 36538 328226
rect 36606 328170 36662 328226
rect 36234 328046 36290 328102
rect 36358 328046 36414 328102
rect 36482 328046 36538 328102
rect 36606 328046 36662 328102
rect 36234 327922 36290 327978
rect 36358 327922 36414 327978
rect 36482 327922 36538 327978
rect 36606 327922 36662 327978
rect 36234 310294 36290 310350
rect 36358 310294 36414 310350
rect 36482 310294 36538 310350
rect 36606 310294 36662 310350
rect 36234 310170 36290 310226
rect 36358 310170 36414 310226
rect 36482 310170 36538 310226
rect 36606 310170 36662 310226
rect 36234 310046 36290 310102
rect 36358 310046 36414 310102
rect 36482 310046 36538 310102
rect 36606 310046 36662 310102
rect 36234 309922 36290 309978
rect 36358 309922 36414 309978
rect 36482 309922 36538 309978
rect 36606 309922 36662 309978
rect 36234 292294 36290 292350
rect 36358 292294 36414 292350
rect 36482 292294 36538 292350
rect 36606 292294 36662 292350
rect 36234 292170 36290 292226
rect 36358 292170 36414 292226
rect 36482 292170 36538 292226
rect 36606 292170 36662 292226
rect 36234 292046 36290 292102
rect 36358 292046 36414 292102
rect 36482 292046 36538 292102
rect 36606 292046 36662 292102
rect 36234 291922 36290 291978
rect 36358 291922 36414 291978
rect 36482 291922 36538 291978
rect 36606 291922 36662 291978
rect 36234 274294 36290 274350
rect 36358 274294 36414 274350
rect 36482 274294 36538 274350
rect 36606 274294 36662 274350
rect 36234 274170 36290 274226
rect 36358 274170 36414 274226
rect 36482 274170 36538 274226
rect 36606 274170 36662 274226
rect 36234 274046 36290 274102
rect 36358 274046 36414 274102
rect 36482 274046 36538 274102
rect 36606 274046 36662 274102
rect 36234 273922 36290 273978
rect 36358 273922 36414 273978
rect 36482 273922 36538 273978
rect 36606 273922 36662 273978
rect 36234 256294 36290 256350
rect 36358 256294 36414 256350
rect 36482 256294 36538 256350
rect 36606 256294 36662 256350
rect 36234 256170 36290 256226
rect 36358 256170 36414 256226
rect 36482 256170 36538 256226
rect 36606 256170 36662 256226
rect 36234 256046 36290 256102
rect 36358 256046 36414 256102
rect 36482 256046 36538 256102
rect 36606 256046 36662 256102
rect 36234 255922 36290 255978
rect 36358 255922 36414 255978
rect 36482 255922 36538 255978
rect 36606 255922 36662 255978
rect 36234 238294 36290 238350
rect 36358 238294 36414 238350
rect 36482 238294 36538 238350
rect 36606 238294 36662 238350
rect 36234 238170 36290 238226
rect 36358 238170 36414 238226
rect 36482 238170 36538 238226
rect 36606 238170 36662 238226
rect 36234 238046 36290 238102
rect 36358 238046 36414 238102
rect 36482 238046 36538 238102
rect 36606 238046 36662 238102
rect 36234 237922 36290 237978
rect 36358 237922 36414 237978
rect 36482 237922 36538 237978
rect 36606 237922 36662 237978
rect 36234 220294 36290 220350
rect 36358 220294 36414 220350
rect 36482 220294 36538 220350
rect 36606 220294 36662 220350
rect 36234 220170 36290 220226
rect 36358 220170 36414 220226
rect 36482 220170 36538 220226
rect 36606 220170 36662 220226
rect 36234 220046 36290 220102
rect 36358 220046 36414 220102
rect 36482 220046 36538 220102
rect 36606 220046 36662 220102
rect 36234 219922 36290 219978
rect 36358 219922 36414 219978
rect 36482 219922 36538 219978
rect 36606 219922 36662 219978
rect 36234 202294 36290 202350
rect 36358 202294 36414 202350
rect 36482 202294 36538 202350
rect 36606 202294 36662 202350
rect 36234 202170 36290 202226
rect 36358 202170 36414 202226
rect 36482 202170 36538 202226
rect 36606 202170 36662 202226
rect 36234 202046 36290 202102
rect 36358 202046 36414 202102
rect 36482 202046 36538 202102
rect 36606 202046 36662 202102
rect 36234 201922 36290 201978
rect 36358 201922 36414 201978
rect 36482 201922 36538 201978
rect 36606 201922 36662 201978
rect 36234 184294 36290 184350
rect 36358 184294 36414 184350
rect 36482 184294 36538 184350
rect 36606 184294 36662 184350
rect 36234 184170 36290 184226
rect 36358 184170 36414 184226
rect 36482 184170 36538 184226
rect 36606 184170 36662 184226
rect 36234 184046 36290 184102
rect 36358 184046 36414 184102
rect 36482 184046 36538 184102
rect 36606 184046 36662 184102
rect 36234 183922 36290 183978
rect 36358 183922 36414 183978
rect 36482 183922 36538 183978
rect 36606 183922 36662 183978
rect 36234 166294 36290 166350
rect 36358 166294 36414 166350
rect 36482 166294 36538 166350
rect 36606 166294 36662 166350
rect 36234 166170 36290 166226
rect 36358 166170 36414 166226
rect 36482 166170 36538 166226
rect 36606 166170 36662 166226
rect 36234 166046 36290 166102
rect 36358 166046 36414 166102
rect 36482 166046 36538 166102
rect 36606 166046 36662 166102
rect 36234 165922 36290 165978
rect 36358 165922 36414 165978
rect 36482 165922 36538 165978
rect 36606 165922 36662 165978
rect 36234 148294 36290 148350
rect 36358 148294 36414 148350
rect 36482 148294 36538 148350
rect 36606 148294 36662 148350
rect 36234 148170 36290 148226
rect 36358 148170 36414 148226
rect 36482 148170 36538 148226
rect 36606 148170 36662 148226
rect 36234 148046 36290 148102
rect 36358 148046 36414 148102
rect 36482 148046 36538 148102
rect 36606 148046 36662 148102
rect 36234 147922 36290 147978
rect 36358 147922 36414 147978
rect 36482 147922 36538 147978
rect 36606 147922 36662 147978
rect 36234 130294 36290 130350
rect 36358 130294 36414 130350
rect 36482 130294 36538 130350
rect 36606 130294 36662 130350
rect 36234 130170 36290 130226
rect 36358 130170 36414 130226
rect 36482 130170 36538 130226
rect 36606 130170 36662 130226
rect 36234 130046 36290 130102
rect 36358 130046 36414 130102
rect 36482 130046 36538 130102
rect 36606 130046 36662 130102
rect 36234 129922 36290 129978
rect 36358 129922 36414 129978
rect 36482 129922 36538 129978
rect 36606 129922 36662 129978
rect 36234 112294 36290 112350
rect 36358 112294 36414 112350
rect 36482 112294 36538 112350
rect 36606 112294 36662 112350
rect 36234 112170 36290 112226
rect 36358 112170 36414 112226
rect 36482 112170 36538 112226
rect 36606 112170 36662 112226
rect 36234 112046 36290 112102
rect 36358 112046 36414 112102
rect 36482 112046 36538 112102
rect 36606 112046 36662 112102
rect 36234 111922 36290 111978
rect 36358 111922 36414 111978
rect 36482 111922 36538 111978
rect 36606 111922 36662 111978
rect 36234 94294 36290 94350
rect 36358 94294 36414 94350
rect 36482 94294 36538 94350
rect 36606 94294 36662 94350
rect 36234 94170 36290 94226
rect 36358 94170 36414 94226
rect 36482 94170 36538 94226
rect 36606 94170 36662 94226
rect 36234 94046 36290 94102
rect 36358 94046 36414 94102
rect 36482 94046 36538 94102
rect 36606 94046 36662 94102
rect 36234 93922 36290 93978
rect 36358 93922 36414 93978
rect 36482 93922 36538 93978
rect 36606 93922 36662 93978
rect 36234 76294 36290 76350
rect 36358 76294 36414 76350
rect 36482 76294 36538 76350
rect 36606 76294 36662 76350
rect 36234 76170 36290 76226
rect 36358 76170 36414 76226
rect 36482 76170 36538 76226
rect 36606 76170 36662 76226
rect 36234 76046 36290 76102
rect 36358 76046 36414 76102
rect 36482 76046 36538 76102
rect 36606 76046 36662 76102
rect 36234 75922 36290 75978
rect 36358 75922 36414 75978
rect 36482 75922 36538 75978
rect 36606 75922 36662 75978
rect 31878 64294 31934 64350
rect 32002 64294 32058 64350
rect 31878 64170 31934 64226
rect 32002 64170 32058 64226
rect 31878 64046 31934 64102
rect 32002 64046 32058 64102
rect 31878 63922 31934 63978
rect 32002 63922 32058 63978
rect 31052 60362 31108 60418
rect 27692 49562 27748 49618
rect 36234 58294 36290 58350
rect 36358 58294 36414 58350
rect 36482 58294 36538 58350
rect 36606 58294 36662 58350
rect 36234 58170 36290 58226
rect 36358 58170 36414 58226
rect 36482 58170 36538 58226
rect 36606 58170 36662 58226
rect 36234 58046 36290 58102
rect 36358 58046 36414 58102
rect 36482 58046 36538 58102
rect 36606 58046 36662 58102
rect 36234 57922 36290 57978
rect 36358 57922 36414 57978
rect 36482 57922 36538 57978
rect 36606 57922 36662 57978
rect 19292 48662 19348 48718
rect 31878 46294 31934 46350
rect 32002 46294 32058 46350
rect 31878 46170 31934 46226
rect 32002 46170 32058 46226
rect 31878 46046 31934 46102
rect 32002 46046 32058 46102
rect 31878 45922 31934 45978
rect 32002 45922 32058 45978
rect 16518 40294 16574 40350
rect 16642 40294 16698 40350
rect 16518 40170 16574 40226
rect 16642 40170 16698 40226
rect 16518 40046 16574 40102
rect 16642 40046 16698 40102
rect 16518 39922 16574 39978
rect 16642 39922 16698 39978
rect 36234 40294 36290 40350
rect 36358 40294 36414 40350
rect 36482 40294 36538 40350
rect 36606 40294 36662 40350
rect 36234 40170 36290 40226
rect 36358 40170 36414 40226
rect 36482 40170 36538 40226
rect 36606 40170 36662 40226
rect 36234 40046 36290 40102
rect 36358 40046 36414 40102
rect 36482 40046 36538 40102
rect 36606 40046 36662 40102
rect 36234 39922 36290 39978
rect 36358 39922 36414 39978
rect 36482 39922 36538 39978
rect 36606 39922 36662 39978
rect 31878 28294 31934 28350
rect 32002 28294 32058 28350
rect 31878 28170 31934 28226
rect 32002 28170 32058 28226
rect 31878 28046 31934 28102
rect 32002 28046 32058 28102
rect 31878 27922 31934 27978
rect 32002 27922 32058 27978
rect 16518 22294 16574 22350
rect 16642 22294 16698 22350
rect 16518 22170 16574 22226
rect 16642 22170 16698 22226
rect 16518 22046 16574 22102
rect 16642 22046 16698 22102
rect 16518 21922 16574 21978
rect 16642 21922 16698 21978
rect 36234 22294 36290 22350
rect 36358 22294 36414 22350
rect 36482 22294 36538 22350
rect 36606 22294 36662 22350
rect 36234 22170 36290 22226
rect 36358 22170 36414 22226
rect 36482 22170 36538 22226
rect 36606 22170 36662 22226
rect 36234 22046 36290 22102
rect 36358 22046 36414 22102
rect 36482 22046 36538 22102
rect 36606 22046 36662 22102
rect 36234 21922 36290 21978
rect 36358 21922 36414 21978
rect 36482 21922 36538 21978
rect 36606 21922 36662 21978
rect 9234 10294 9290 10350
rect 9358 10294 9414 10350
rect 9482 10294 9538 10350
rect 9606 10294 9662 10350
rect 9234 10170 9290 10226
rect 9358 10170 9414 10226
rect 9482 10170 9538 10226
rect 9606 10170 9662 10226
rect 9234 10046 9290 10102
rect 9358 10046 9414 10102
rect 9482 10046 9538 10102
rect 9606 10046 9662 10102
rect 9234 9922 9290 9978
rect 9358 9922 9414 9978
rect 9482 9922 9538 9978
rect 9606 9922 9662 9978
rect 5514 4294 5570 4350
rect 5638 4294 5694 4350
rect 5762 4294 5818 4350
rect 5886 4294 5942 4350
rect 5514 4170 5570 4226
rect 5638 4170 5694 4226
rect 5762 4170 5818 4226
rect 5886 4170 5942 4226
rect 5514 4046 5570 4102
rect 5638 4046 5694 4102
rect 5762 4046 5818 4102
rect 5886 4046 5942 4102
rect 5514 3922 5570 3978
rect 5638 3922 5694 3978
rect 5762 3922 5818 3978
rect 5886 3922 5942 3978
rect 5514 -216 5570 -160
rect 5638 -216 5694 -160
rect 5762 -216 5818 -160
rect 5886 -216 5942 -160
rect 5514 -340 5570 -284
rect 5638 -340 5694 -284
rect 5762 -340 5818 -284
rect 5886 -340 5942 -284
rect 5514 -464 5570 -408
rect 5638 -464 5694 -408
rect 5762 -464 5818 -408
rect 5886 -464 5942 -408
rect 5514 -588 5570 -532
rect 5638 -588 5694 -532
rect 5762 -588 5818 -532
rect 5886 -588 5942 -532
rect -1820 -1176 -1764 -1120
rect -1696 -1176 -1640 -1120
rect -1572 -1176 -1516 -1120
rect -1448 -1176 -1392 -1120
rect -1820 -1300 -1764 -1244
rect -1696 -1300 -1640 -1244
rect -1572 -1300 -1516 -1244
rect -1448 -1300 -1392 -1244
rect -1820 -1424 -1764 -1368
rect -1696 -1424 -1640 -1368
rect -1572 -1424 -1516 -1368
rect -1448 -1424 -1392 -1368
rect -1820 -1548 -1764 -1492
rect -1696 -1548 -1640 -1492
rect -1572 -1548 -1516 -1492
rect -1448 -1548 -1392 -1492
rect 31878 10294 31934 10350
rect 32002 10294 32058 10350
rect 31878 10170 31934 10226
rect 32002 10170 32058 10226
rect 31878 10046 31934 10102
rect 32002 10046 32058 10102
rect 31878 9922 31934 9978
rect 32002 9922 32058 9978
rect 36234 4294 36290 4350
rect 36358 4294 36414 4350
rect 36482 4294 36538 4350
rect 36606 4294 36662 4350
rect 36234 4170 36290 4226
rect 36358 4170 36414 4226
rect 36482 4170 36538 4226
rect 36606 4170 36662 4226
rect 36234 4046 36290 4102
rect 36358 4046 36414 4102
rect 36482 4046 36538 4102
rect 36606 4046 36662 4102
rect 36234 3922 36290 3978
rect 36358 3922 36414 3978
rect 36482 3922 36538 3978
rect 36606 3922 36662 3978
rect 9234 -1176 9290 -1120
rect 9358 -1176 9414 -1120
rect 9482 -1176 9538 -1120
rect 9606 -1176 9662 -1120
rect 9234 -1300 9290 -1244
rect 9358 -1300 9414 -1244
rect 9482 -1300 9538 -1244
rect 9606 -1300 9662 -1244
rect 9234 -1424 9290 -1368
rect 9358 -1424 9414 -1368
rect 9482 -1424 9538 -1368
rect 9606 -1424 9662 -1368
rect 9234 -1548 9290 -1492
rect 9358 -1548 9414 -1492
rect 9482 -1548 9538 -1492
rect 9606 -1548 9662 -1492
rect 36234 -216 36290 -160
rect 36358 -216 36414 -160
rect 36482 -216 36538 -160
rect 36606 -216 36662 -160
rect 36234 -340 36290 -284
rect 36358 -340 36414 -284
rect 36482 -340 36538 -284
rect 36606 -340 36662 -284
rect 36234 -464 36290 -408
rect 36358 -464 36414 -408
rect 36482 -464 36538 -408
rect 36606 -464 36662 -408
rect 36234 -588 36290 -532
rect 36358 -588 36414 -532
rect 36482 -588 36538 -532
rect 36606 -588 36662 -532
rect 39954 598116 40010 598172
rect 40078 598116 40134 598172
rect 40202 598116 40258 598172
rect 40326 598116 40382 598172
rect 39954 597992 40010 598048
rect 40078 597992 40134 598048
rect 40202 597992 40258 598048
rect 40326 597992 40382 598048
rect 39954 597868 40010 597924
rect 40078 597868 40134 597924
rect 40202 597868 40258 597924
rect 40326 597868 40382 597924
rect 39954 597744 40010 597800
rect 40078 597744 40134 597800
rect 40202 597744 40258 597800
rect 40326 597744 40382 597800
rect 39954 586294 40010 586350
rect 40078 586294 40134 586350
rect 40202 586294 40258 586350
rect 40326 586294 40382 586350
rect 39954 586170 40010 586226
rect 40078 586170 40134 586226
rect 40202 586170 40258 586226
rect 40326 586170 40382 586226
rect 39954 586046 40010 586102
rect 40078 586046 40134 586102
rect 40202 586046 40258 586102
rect 40326 586046 40382 586102
rect 39954 585922 40010 585978
rect 40078 585922 40134 585978
rect 40202 585922 40258 585978
rect 40326 585922 40382 585978
rect 39954 568294 40010 568350
rect 40078 568294 40134 568350
rect 40202 568294 40258 568350
rect 40326 568294 40382 568350
rect 39954 568170 40010 568226
rect 40078 568170 40134 568226
rect 40202 568170 40258 568226
rect 40326 568170 40382 568226
rect 39954 568046 40010 568102
rect 40078 568046 40134 568102
rect 40202 568046 40258 568102
rect 40326 568046 40382 568102
rect 39954 567922 40010 567978
rect 40078 567922 40134 567978
rect 40202 567922 40258 567978
rect 40326 567922 40382 567978
rect 39954 550294 40010 550350
rect 40078 550294 40134 550350
rect 40202 550294 40258 550350
rect 40326 550294 40382 550350
rect 39954 550170 40010 550226
rect 40078 550170 40134 550226
rect 40202 550170 40258 550226
rect 40326 550170 40382 550226
rect 39954 550046 40010 550102
rect 40078 550046 40134 550102
rect 40202 550046 40258 550102
rect 40326 550046 40382 550102
rect 39954 549922 40010 549978
rect 40078 549922 40134 549978
rect 40202 549922 40258 549978
rect 40326 549922 40382 549978
rect 39954 532294 40010 532350
rect 40078 532294 40134 532350
rect 40202 532294 40258 532350
rect 40326 532294 40382 532350
rect 39954 532170 40010 532226
rect 40078 532170 40134 532226
rect 40202 532170 40258 532226
rect 40326 532170 40382 532226
rect 39954 532046 40010 532102
rect 40078 532046 40134 532102
rect 40202 532046 40258 532102
rect 40326 532046 40382 532102
rect 39954 531922 40010 531978
rect 40078 531922 40134 531978
rect 40202 531922 40258 531978
rect 40326 531922 40382 531978
rect 39954 514294 40010 514350
rect 40078 514294 40134 514350
rect 40202 514294 40258 514350
rect 40326 514294 40382 514350
rect 39954 514170 40010 514226
rect 40078 514170 40134 514226
rect 40202 514170 40258 514226
rect 40326 514170 40382 514226
rect 39954 514046 40010 514102
rect 40078 514046 40134 514102
rect 40202 514046 40258 514102
rect 40326 514046 40382 514102
rect 39954 513922 40010 513978
rect 40078 513922 40134 513978
rect 40202 513922 40258 513978
rect 40326 513922 40382 513978
rect 39954 496294 40010 496350
rect 40078 496294 40134 496350
rect 40202 496294 40258 496350
rect 40326 496294 40382 496350
rect 39954 496170 40010 496226
rect 40078 496170 40134 496226
rect 40202 496170 40258 496226
rect 40326 496170 40382 496226
rect 39954 496046 40010 496102
rect 40078 496046 40134 496102
rect 40202 496046 40258 496102
rect 40326 496046 40382 496102
rect 39954 495922 40010 495978
rect 40078 495922 40134 495978
rect 40202 495922 40258 495978
rect 40326 495922 40382 495978
rect 39954 478294 40010 478350
rect 40078 478294 40134 478350
rect 40202 478294 40258 478350
rect 40326 478294 40382 478350
rect 39954 478170 40010 478226
rect 40078 478170 40134 478226
rect 40202 478170 40258 478226
rect 40326 478170 40382 478226
rect 39954 478046 40010 478102
rect 40078 478046 40134 478102
rect 40202 478046 40258 478102
rect 40326 478046 40382 478102
rect 39954 477922 40010 477978
rect 40078 477922 40134 477978
rect 40202 477922 40258 477978
rect 40326 477922 40382 477978
rect 39954 460294 40010 460350
rect 40078 460294 40134 460350
rect 40202 460294 40258 460350
rect 40326 460294 40382 460350
rect 39954 460170 40010 460226
rect 40078 460170 40134 460226
rect 40202 460170 40258 460226
rect 40326 460170 40382 460226
rect 39954 460046 40010 460102
rect 40078 460046 40134 460102
rect 40202 460046 40258 460102
rect 40326 460046 40382 460102
rect 39954 459922 40010 459978
rect 40078 459922 40134 459978
rect 40202 459922 40258 459978
rect 40326 459922 40382 459978
rect 39954 442294 40010 442350
rect 40078 442294 40134 442350
rect 40202 442294 40258 442350
rect 40326 442294 40382 442350
rect 39954 442170 40010 442226
rect 40078 442170 40134 442226
rect 40202 442170 40258 442226
rect 40326 442170 40382 442226
rect 39954 442046 40010 442102
rect 40078 442046 40134 442102
rect 40202 442046 40258 442102
rect 40326 442046 40382 442102
rect 39954 441922 40010 441978
rect 40078 441922 40134 441978
rect 40202 441922 40258 441978
rect 40326 441922 40382 441978
rect 39954 424294 40010 424350
rect 40078 424294 40134 424350
rect 40202 424294 40258 424350
rect 40326 424294 40382 424350
rect 39954 424170 40010 424226
rect 40078 424170 40134 424226
rect 40202 424170 40258 424226
rect 40326 424170 40382 424226
rect 39954 424046 40010 424102
rect 40078 424046 40134 424102
rect 40202 424046 40258 424102
rect 40326 424046 40382 424102
rect 39954 423922 40010 423978
rect 40078 423922 40134 423978
rect 40202 423922 40258 423978
rect 40326 423922 40382 423978
rect 39954 406294 40010 406350
rect 40078 406294 40134 406350
rect 40202 406294 40258 406350
rect 40326 406294 40382 406350
rect 39954 406170 40010 406226
rect 40078 406170 40134 406226
rect 40202 406170 40258 406226
rect 40326 406170 40382 406226
rect 39954 406046 40010 406102
rect 40078 406046 40134 406102
rect 40202 406046 40258 406102
rect 40326 406046 40382 406102
rect 39954 405922 40010 405978
rect 40078 405922 40134 405978
rect 40202 405922 40258 405978
rect 40326 405922 40382 405978
rect 39954 388294 40010 388350
rect 40078 388294 40134 388350
rect 40202 388294 40258 388350
rect 40326 388294 40382 388350
rect 39954 388170 40010 388226
rect 40078 388170 40134 388226
rect 40202 388170 40258 388226
rect 40326 388170 40382 388226
rect 39954 388046 40010 388102
rect 40078 388046 40134 388102
rect 40202 388046 40258 388102
rect 40326 388046 40382 388102
rect 39954 387922 40010 387978
rect 40078 387922 40134 387978
rect 40202 387922 40258 387978
rect 40326 387922 40382 387978
rect 39954 370294 40010 370350
rect 40078 370294 40134 370350
rect 40202 370294 40258 370350
rect 40326 370294 40382 370350
rect 39954 370170 40010 370226
rect 40078 370170 40134 370226
rect 40202 370170 40258 370226
rect 40326 370170 40382 370226
rect 39954 370046 40010 370102
rect 40078 370046 40134 370102
rect 40202 370046 40258 370102
rect 40326 370046 40382 370102
rect 39954 369922 40010 369978
rect 40078 369922 40134 369978
rect 40202 369922 40258 369978
rect 40326 369922 40382 369978
rect 39954 352294 40010 352350
rect 40078 352294 40134 352350
rect 40202 352294 40258 352350
rect 40326 352294 40382 352350
rect 39954 352170 40010 352226
rect 40078 352170 40134 352226
rect 40202 352170 40258 352226
rect 40326 352170 40382 352226
rect 39954 352046 40010 352102
rect 40078 352046 40134 352102
rect 40202 352046 40258 352102
rect 40326 352046 40382 352102
rect 39954 351922 40010 351978
rect 40078 351922 40134 351978
rect 40202 351922 40258 351978
rect 40326 351922 40382 351978
rect 39954 334294 40010 334350
rect 40078 334294 40134 334350
rect 40202 334294 40258 334350
rect 40326 334294 40382 334350
rect 39954 334170 40010 334226
rect 40078 334170 40134 334226
rect 40202 334170 40258 334226
rect 40326 334170 40382 334226
rect 39954 334046 40010 334102
rect 40078 334046 40134 334102
rect 40202 334046 40258 334102
rect 40326 334046 40382 334102
rect 39954 333922 40010 333978
rect 40078 333922 40134 333978
rect 40202 333922 40258 333978
rect 40326 333922 40382 333978
rect 66954 597156 67010 597212
rect 67078 597156 67134 597212
rect 67202 597156 67258 597212
rect 67326 597156 67382 597212
rect 66954 597032 67010 597088
rect 67078 597032 67134 597088
rect 67202 597032 67258 597088
rect 67326 597032 67382 597088
rect 66954 596908 67010 596964
rect 67078 596908 67134 596964
rect 67202 596908 67258 596964
rect 67326 596908 67382 596964
rect 66954 596784 67010 596840
rect 67078 596784 67134 596840
rect 67202 596784 67258 596840
rect 67326 596784 67382 596840
rect 66954 580294 67010 580350
rect 67078 580294 67134 580350
rect 67202 580294 67258 580350
rect 67326 580294 67382 580350
rect 66954 580170 67010 580226
rect 67078 580170 67134 580226
rect 67202 580170 67258 580226
rect 67326 580170 67382 580226
rect 66954 580046 67010 580102
rect 67078 580046 67134 580102
rect 67202 580046 67258 580102
rect 67326 580046 67382 580102
rect 66954 579922 67010 579978
rect 67078 579922 67134 579978
rect 67202 579922 67258 579978
rect 67326 579922 67382 579978
rect 66954 562294 67010 562350
rect 67078 562294 67134 562350
rect 67202 562294 67258 562350
rect 67326 562294 67382 562350
rect 66954 562170 67010 562226
rect 67078 562170 67134 562226
rect 67202 562170 67258 562226
rect 67326 562170 67382 562226
rect 66954 562046 67010 562102
rect 67078 562046 67134 562102
rect 67202 562046 67258 562102
rect 67326 562046 67382 562102
rect 66954 561922 67010 561978
rect 67078 561922 67134 561978
rect 67202 561922 67258 561978
rect 67326 561922 67382 561978
rect 66954 544294 67010 544350
rect 67078 544294 67134 544350
rect 67202 544294 67258 544350
rect 67326 544294 67382 544350
rect 66954 544170 67010 544226
rect 67078 544170 67134 544226
rect 67202 544170 67258 544226
rect 67326 544170 67382 544226
rect 66954 544046 67010 544102
rect 67078 544046 67134 544102
rect 67202 544046 67258 544102
rect 67326 544046 67382 544102
rect 66954 543922 67010 543978
rect 67078 543922 67134 543978
rect 67202 543922 67258 543978
rect 67326 543922 67382 543978
rect 66954 526294 67010 526350
rect 67078 526294 67134 526350
rect 67202 526294 67258 526350
rect 67326 526294 67382 526350
rect 66954 526170 67010 526226
rect 67078 526170 67134 526226
rect 67202 526170 67258 526226
rect 67326 526170 67382 526226
rect 66954 526046 67010 526102
rect 67078 526046 67134 526102
rect 67202 526046 67258 526102
rect 67326 526046 67382 526102
rect 66954 525922 67010 525978
rect 67078 525922 67134 525978
rect 67202 525922 67258 525978
rect 67326 525922 67382 525978
rect 66954 508294 67010 508350
rect 67078 508294 67134 508350
rect 67202 508294 67258 508350
rect 67326 508294 67382 508350
rect 66954 508170 67010 508226
rect 67078 508170 67134 508226
rect 67202 508170 67258 508226
rect 67326 508170 67382 508226
rect 66954 508046 67010 508102
rect 67078 508046 67134 508102
rect 67202 508046 67258 508102
rect 67326 508046 67382 508102
rect 66954 507922 67010 507978
rect 67078 507922 67134 507978
rect 67202 507922 67258 507978
rect 67326 507922 67382 507978
rect 66954 490294 67010 490350
rect 67078 490294 67134 490350
rect 67202 490294 67258 490350
rect 67326 490294 67382 490350
rect 66954 490170 67010 490226
rect 67078 490170 67134 490226
rect 67202 490170 67258 490226
rect 67326 490170 67382 490226
rect 66954 490046 67010 490102
rect 67078 490046 67134 490102
rect 67202 490046 67258 490102
rect 67326 490046 67382 490102
rect 66954 489922 67010 489978
rect 67078 489922 67134 489978
rect 67202 489922 67258 489978
rect 67326 489922 67382 489978
rect 66954 472294 67010 472350
rect 67078 472294 67134 472350
rect 67202 472294 67258 472350
rect 67326 472294 67382 472350
rect 66954 472170 67010 472226
rect 67078 472170 67134 472226
rect 67202 472170 67258 472226
rect 67326 472170 67382 472226
rect 66954 472046 67010 472102
rect 67078 472046 67134 472102
rect 67202 472046 67258 472102
rect 67326 472046 67382 472102
rect 66954 471922 67010 471978
rect 67078 471922 67134 471978
rect 67202 471922 67258 471978
rect 67326 471922 67382 471978
rect 66954 454294 67010 454350
rect 67078 454294 67134 454350
rect 67202 454294 67258 454350
rect 67326 454294 67382 454350
rect 66954 454170 67010 454226
rect 67078 454170 67134 454226
rect 67202 454170 67258 454226
rect 67326 454170 67382 454226
rect 66954 454046 67010 454102
rect 67078 454046 67134 454102
rect 67202 454046 67258 454102
rect 67326 454046 67382 454102
rect 66954 453922 67010 453978
rect 67078 453922 67134 453978
rect 67202 453922 67258 453978
rect 67326 453922 67382 453978
rect 66954 436294 67010 436350
rect 67078 436294 67134 436350
rect 67202 436294 67258 436350
rect 67326 436294 67382 436350
rect 66954 436170 67010 436226
rect 67078 436170 67134 436226
rect 67202 436170 67258 436226
rect 67326 436170 67382 436226
rect 66954 436046 67010 436102
rect 67078 436046 67134 436102
rect 67202 436046 67258 436102
rect 67326 436046 67382 436102
rect 66954 435922 67010 435978
rect 67078 435922 67134 435978
rect 67202 435922 67258 435978
rect 67326 435922 67382 435978
rect 66954 418294 67010 418350
rect 67078 418294 67134 418350
rect 67202 418294 67258 418350
rect 67326 418294 67382 418350
rect 66954 418170 67010 418226
rect 67078 418170 67134 418226
rect 67202 418170 67258 418226
rect 67326 418170 67382 418226
rect 66954 418046 67010 418102
rect 67078 418046 67134 418102
rect 67202 418046 67258 418102
rect 67326 418046 67382 418102
rect 66954 417922 67010 417978
rect 67078 417922 67134 417978
rect 67202 417922 67258 417978
rect 67326 417922 67382 417978
rect 66954 400294 67010 400350
rect 67078 400294 67134 400350
rect 67202 400294 67258 400350
rect 67326 400294 67382 400350
rect 66954 400170 67010 400226
rect 67078 400170 67134 400226
rect 67202 400170 67258 400226
rect 67326 400170 67382 400226
rect 66954 400046 67010 400102
rect 67078 400046 67134 400102
rect 67202 400046 67258 400102
rect 67326 400046 67382 400102
rect 66954 399922 67010 399978
rect 67078 399922 67134 399978
rect 67202 399922 67258 399978
rect 67326 399922 67382 399978
rect 66954 382294 67010 382350
rect 67078 382294 67134 382350
rect 67202 382294 67258 382350
rect 67326 382294 67382 382350
rect 66954 382170 67010 382226
rect 67078 382170 67134 382226
rect 67202 382170 67258 382226
rect 67326 382170 67382 382226
rect 66954 382046 67010 382102
rect 67078 382046 67134 382102
rect 67202 382046 67258 382102
rect 67326 382046 67382 382102
rect 66954 381922 67010 381978
rect 67078 381922 67134 381978
rect 67202 381922 67258 381978
rect 67326 381922 67382 381978
rect 66954 364294 67010 364350
rect 67078 364294 67134 364350
rect 67202 364294 67258 364350
rect 67326 364294 67382 364350
rect 66954 364170 67010 364226
rect 67078 364170 67134 364226
rect 67202 364170 67258 364226
rect 67326 364170 67382 364226
rect 66954 364046 67010 364102
rect 67078 364046 67134 364102
rect 67202 364046 67258 364102
rect 67326 364046 67382 364102
rect 66954 363922 67010 363978
rect 67078 363922 67134 363978
rect 67202 363922 67258 363978
rect 67326 363922 67382 363978
rect 66954 346294 67010 346350
rect 67078 346294 67134 346350
rect 67202 346294 67258 346350
rect 67326 346294 67382 346350
rect 66954 346170 67010 346226
rect 67078 346170 67134 346226
rect 67202 346170 67258 346226
rect 67326 346170 67382 346226
rect 66954 346046 67010 346102
rect 67078 346046 67134 346102
rect 67202 346046 67258 346102
rect 67326 346046 67382 346102
rect 66954 345922 67010 345978
rect 67078 345922 67134 345978
rect 67202 345922 67258 345978
rect 67326 345922 67382 345978
rect 66954 328294 67010 328350
rect 67078 328294 67134 328350
rect 67202 328294 67258 328350
rect 67326 328294 67382 328350
rect 66954 328170 67010 328226
rect 67078 328170 67134 328226
rect 67202 328170 67258 328226
rect 67326 328170 67382 328226
rect 66954 328046 67010 328102
rect 67078 328046 67134 328102
rect 67202 328046 67258 328102
rect 67326 328046 67382 328102
rect 66954 327922 67010 327978
rect 67078 327922 67134 327978
rect 67202 327922 67258 327978
rect 67326 327922 67382 327978
rect 39954 316294 40010 316350
rect 40078 316294 40134 316350
rect 40202 316294 40258 316350
rect 40326 316294 40382 316350
rect 39954 316170 40010 316226
rect 40078 316170 40134 316226
rect 40202 316170 40258 316226
rect 40326 316170 40382 316226
rect 39954 316046 40010 316102
rect 40078 316046 40134 316102
rect 40202 316046 40258 316102
rect 40326 316046 40382 316102
rect 39954 315922 40010 315978
rect 40078 315922 40134 315978
rect 40202 315922 40258 315978
rect 40326 315922 40382 315978
rect 39954 298294 40010 298350
rect 40078 298294 40134 298350
rect 40202 298294 40258 298350
rect 40326 298294 40382 298350
rect 39954 298170 40010 298226
rect 40078 298170 40134 298226
rect 40202 298170 40258 298226
rect 40326 298170 40382 298226
rect 39954 298046 40010 298102
rect 40078 298046 40134 298102
rect 40202 298046 40258 298102
rect 40326 298046 40382 298102
rect 39954 297922 40010 297978
rect 40078 297922 40134 297978
rect 40202 297922 40258 297978
rect 40326 297922 40382 297978
rect 39954 280294 40010 280350
rect 40078 280294 40134 280350
rect 40202 280294 40258 280350
rect 40326 280294 40382 280350
rect 39954 280170 40010 280226
rect 40078 280170 40134 280226
rect 40202 280170 40258 280226
rect 40326 280170 40382 280226
rect 39954 280046 40010 280102
rect 40078 280046 40134 280102
rect 40202 280046 40258 280102
rect 40326 280046 40382 280102
rect 39954 279922 40010 279978
rect 40078 279922 40134 279978
rect 40202 279922 40258 279978
rect 40326 279922 40382 279978
rect 39954 262294 40010 262350
rect 40078 262294 40134 262350
rect 40202 262294 40258 262350
rect 40326 262294 40382 262350
rect 39954 262170 40010 262226
rect 40078 262170 40134 262226
rect 40202 262170 40258 262226
rect 40326 262170 40382 262226
rect 39954 262046 40010 262102
rect 40078 262046 40134 262102
rect 40202 262046 40258 262102
rect 40326 262046 40382 262102
rect 39954 261922 40010 261978
rect 40078 261922 40134 261978
rect 40202 261922 40258 261978
rect 40326 261922 40382 261978
rect 39954 244294 40010 244350
rect 40078 244294 40134 244350
rect 40202 244294 40258 244350
rect 40326 244294 40382 244350
rect 39954 244170 40010 244226
rect 40078 244170 40134 244226
rect 40202 244170 40258 244226
rect 40326 244170 40382 244226
rect 39954 244046 40010 244102
rect 40078 244046 40134 244102
rect 40202 244046 40258 244102
rect 40326 244046 40382 244102
rect 39954 243922 40010 243978
rect 40078 243922 40134 243978
rect 40202 243922 40258 243978
rect 40326 243922 40382 243978
rect 39954 226294 40010 226350
rect 40078 226294 40134 226350
rect 40202 226294 40258 226350
rect 40326 226294 40382 226350
rect 39954 226170 40010 226226
rect 40078 226170 40134 226226
rect 40202 226170 40258 226226
rect 40326 226170 40382 226226
rect 39954 226046 40010 226102
rect 40078 226046 40134 226102
rect 40202 226046 40258 226102
rect 40326 226046 40382 226102
rect 39954 225922 40010 225978
rect 40078 225922 40134 225978
rect 40202 225922 40258 225978
rect 40326 225922 40382 225978
rect 39954 208294 40010 208350
rect 40078 208294 40134 208350
rect 40202 208294 40258 208350
rect 40326 208294 40382 208350
rect 39954 208170 40010 208226
rect 40078 208170 40134 208226
rect 40202 208170 40258 208226
rect 40326 208170 40382 208226
rect 39954 208046 40010 208102
rect 40078 208046 40134 208102
rect 40202 208046 40258 208102
rect 40326 208046 40382 208102
rect 39954 207922 40010 207978
rect 40078 207922 40134 207978
rect 40202 207922 40258 207978
rect 40326 207922 40382 207978
rect 39954 190294 40010 190350
rect 40078 190294 40134 190350
rect 40202 190294 40258 190350
rect 40326 190294 40382 190350
rect 39954 190170 40010 190226
rect 40078 190170 40134 190226
rect 40202 190170 40258 190226
rect 40326 190170 40382 190226
rect 39954 190046 40010 190102
rect 40078 190046 40134 190102
rect 40202 190046 40258 190102
rect 40326 190046 40382 190102
rect 39954 189922 40010 189978
rect 40078 189922 40134 189978
rect 40202 189922 40258 189978
rect 40326 189922 40382 189978
rect 39954 172294 40010 172350
rect 40078 172294 40134 172350
rect 40202 172294 40258 172350
rect 40326 172294 40382 172350
rect 39954 172170 40010 172226
rect 40078 172170 40134 172226
rect 40202 172170 40258 172226
rect 40326 172170 40382 172226
rect 39954 172046 40010 172102
rect 40078 172046 40134 172102
rect 40202 172046 40258 172102
rect 40326 172046 40382 172102
rect 39954 171922 40010 171978
rect 40078 171922 40134 171978
rect 40202 171922 40258 171978
rect 40326 171922 40382 171978
rect 39954 154294 40010 154350
rect 40078 154294 40134 154350
rect 40202 154294 40258 154350
rect 40326 154294 40382 154350
rect 39954 154170 40010 154226
rect 40078 154170 40134 154226
rect 40202 154170 40258 154226
rect 40326 154170 40382 154226
rect 39954 154046 40010 154102
rect 40078 154046 40134 154102
rect 40202 154046 40258 154102
rect 40326 154046 40382 154102
rect 39954 153922 40010 153978
rect 40078 153922 40134 153978
rect 40202 153922 40258 153978
rect 40326 153922 40382 153978
rect 39954 136294 40010 136350
rect 40078 136294 40134 136350
rect 40202 136294 40258 136350
rect 40326 136294 40382 136350
rect 39954 136170 40010 136226
rect 40078 136170 40134 136226
rect 40202 136170 40258 136226
rect 40326 136170 40382 136226
rect 39954 136046 40010 136102
rect 40078 136046 40134 136102
rect 40202 136046 40258 136102
rect 40326 136046 40382 136102
rect 39954 135922 40010 135978
rect 40078 135922 40134 135978
rect 40202 135922 40258 135978
rect 40326 135922 40382 135978
rect 39954 118294 40010 118350
rect 40078 118294 40134 118350
rect 40202 118294 40258 118350
rect 40326 118294 40382 118350
rect 39954 118170 40010 118226
rect 40078 118170 40134 118226
rect 40202 118170 40258 118226
rect 40326 118170 40382 118226
rect 39954 118046 40010 118102
rect 40078 118046 40134 118102
rect 40202 118046 40258 118102
rect 40326 118046 40382 118102
rect 39954 117922 40010 117978
rect 40078 117922 40134 117978
rect 40202 117922 40258 117978
rect 40326 117922 40382 117978
rect 39954 100294 40010 100350
rect 40078 100294 40134 100350
rect 40202 100294 40258 100350
rect 40326 100294 40382 100350
rect 39954 100170 40010 100226
rect 40078 100170 40134 100226
rect 40202 100170 40258 100226
rect 40326 100170 40382 100226
rect 39954 100046 40010 100102
rect 40078 100046 40134 100102
rect 40202 100046 40258 100102
rect 40326 100046 40382 100102
rect 39954 99922 40010 99978
rect 40078 99922 40134 99978
rect 40202 99922 40258 99978
rect 40326 99922 40382 99978
rect 39954 82294 40010 82350
rect 40078 82294 40134 82350
rect 40202 82294 40258 82350
rect 40326 82294 40382 82350
rect 39954 82170 40010 82226
rect 40078 82170 40134 82226
rect 40202 82170 40258 82226
rect 40326 82170 40382 82226
rect 39954 82046 40010 82102
rect 40078 82046 40134 82102
rect 40202 82046 40258 82102
rect 40326 82046 40382 82102
rect 39954 81922 40010 81978
rect 40078 81922 40134 81978
rect 40202 81922 40258 81978
rect 40326 81922 40382 81978
rect 39954 64294 40010 64350
rect 40078 64294 40134 64350
rect 40202 64294 40258 64350
rect 40326 64294 40382 64350
rect 39954 64170 40010 64226
rect 40078 64170 40134 64226
rect 40202 64170 40258 64226
rect 40326 64170 40382 64226
rect 39954 64046 40010 64102
rect 40078 64046 40134 64102
rect 40202 64046 40258 64102
rect 40326 64046 40382 64102
rect 39954 63922 40010 63978
rect 40078 63922 40134 63978
rect 40202 63922 40258 63978
rect 40326 63922 40382 63978
rect 39954 46294 40010 46350
rect 40078 46294 40134 46350
rect 40202 46294 40258 46350
rect 40326 46294 40382 46350
rect 39954 46170 40010 46226
rect 40078 46170 40134 46226
rect 40202 46170 40258 46226
rect 40326 46170 40382 46226
rect 39954 46046 40010 46102
rect 40078 46046 40134 46102
rect 40202 46046 40258 46102
rect 40326 46046 40382 46102
rect 39954 45922 40010 45978
rect 40078 45922 40134 45978
rect 40202 45922 40258 45978
rect 40326 45922 40382 45978
rect 39954 28294 40010 28350
rect 40078 28294 40134 28350
rect 40202 28294 40258 28350
rect 40326 28294 40382 28350
rect 39954 28170 40010 28226
rect 40078 28170 40134 28226
rect 40202 28170 40258 28226
rect 40326 28170 40382 28226
rect 39954 28046 40010 28102
rect 40078 28046 40134 28102
rect 40202 28046 40258 28102
rect 40326 28046 40382 28102
rect 39954 27922 40010 27978
rect 40078 27922 40134 27978
rect 40202 27922 40258 27978
rect 40326 27922 40382 27978
rect 39954 10294 40010 10350
rect 40078 10294 40134 10350
rect 40202 10294 40258 10350
rect 40326 10294 40382 10350
rect 39954 10170 40010 10226
rect 40078 10170 40134 10226
rect 40202 10170 40258 10226
rect 40326 10170 40382 10226
rect 39954 10046 40010 10102
rect 40078 10046 40134 10102
rect 40202 10046 40258 10102
rect 40326 10046 40382 10102
rect 39954 9922 40010 9978
rect 40078 9922 40134 9978
rect 40202 9922 40258 9978
rect 40326 9922 40382 9978
rect 42476 16802 42532 16858
rect 40908 5462 40964 5518
rect 43148 8522 43204 8578
rect 46732 34622 46788 34678
rect 46620 31202 46676 31258
rect 46508 25262 46564 25318
rect 44716 15182 44772 15238
rect 44268 5102 44324 5158
rect 45612 11942 45668 11998
rect 44940 7802 44996 7858
rect 46620 3662 46676 3718
rect 45836 3332 45892 3358
rect 45836 3302 45892 3332
rect 43820 2762 43876 2818
rect 43596 1502 43652 1558
rect 46844 14462 46900 14518
rect 47238 58294 47294 58350
rect 47362 58294 47418 58350
rect 47238 58170 47294 58226
rect 47362 58170 47418 58226
rect 47238 58046 47294 58102
rect 47362 58046 47418 58102
rect 47238 57922 47294 57978
rect 47362 57922 47418 57978
rect 47238 40294 47294 40350
rect 47362 40294 47418 40350
rect 47238 40170 47294 40226
rect 47362 40170 47418 40226
rect 47238 40046 47294 40102
rect 47362 40046 47418 40102
rect 47238 39922 47294 39978
rect 47362 39922 47418 39978
rect 47238 22294 47294 22350
rect 47362 22294 47418 22350
rect 47238 22170 47294 22226
rect 47362 22170 47418 22226
rect 47238 22046 47294 22102
rect 47362 22046 47418 22102
rect 47238 21922 47294 21978
rect 47362 21922 47418 21978
rect 46956 14102 47012 14158
rect 66954 310294 67010 310350
rect 67078 310294 67134 310350
rect 67202 310294 67258 310350
rect 67326 310294 67382 310350
rect 66954 310170 67010 310226
rect 67078 310170 67134 310226
rect 67202 310170 67258 310226
rect 67326 310170 67382 310226
rect 66954 310046 67010 310102
rect 67078 310046 67134 310102
rect 67202 310046 67258 310102
rect 67326 310046 67382 310102
rect 66954 309922 67010 309978
rect 67078 309922 67134 309978
rect 67202 309922 67258 309978
rect 67326 309922 67382 309978
rect 66954 292294 67010 292350
rect 67078 292294 67134 292350
rect 67202 292294 67258 292350
rect 67326 292294 67382 292350
rect 66954 292170 67010 292226
rect 67078 292170 67134 292226
rect 67202 292170 67258 292226
rect 67326 292170 67382 292226
rect 66954 292046 67010 292102
rect 67078 292046 67134 292102
rect 67202 292046 67258 292102
rect 67326 292046 67382 292102
rect 66954 291922 67010 291978
rect 67078 291922 67134 291978
rect 67202 291922 67258 291978
rect 67326 291922 67382 291978
rect 66954 274294 67010 274350
rect 67078 274294 67134 274350
rect 67202 274294 67258 274350
rect 67326 274294 67382 274350
rect 66954 274170 67010 274226
rect 67078 274170 67134 274226
rect 67202 274170 67258 274226
rect 67326 274170 67382 274226
rect 66954 274046 67010 274102
rect 67078 274046 67134 274102
rect 67202 274046 67258 274102
rect 67326 274046 67382 274102
rect 66954 273922 67010 273978
rect 67078 273922 67134 273978
rect 67202 273922 67258 273978
rect 67326 273922 67382 273978
rect 66954 256294 67010 256350
rect 67078 256294 67134 256350
rect 67202 256294 67258 256350
rect 67326 256294 67382 256350
rect 66954 256170 67010 256226
rect 67078 256170 67134 256226
rect 67202 256170 67258 256226
rect 67326 256170 67382 256226
rect 66954 256046 67010 256102
rect 67078 256046 67134 256102
rect 67202 256046 67258 256102
rect 67326 256046 67382 256102
rect 66954 255922 67010 255978
rect 67078 255922 67134 255978
rect 67202 255922 67258 255978
rect 67326 255922 67382 255978
rect 66954 238294 67010 238350
rect 67078 238294 67134 238350
rect 67202 238294 67258 238350
rect 67326 238294 67382 238350
rect 66954 238170 67010 238226
rect 67078 238170 67134 238226
rect 67202 238170 67258 238226
rect 67326 238170 67382 238226
rect 66954 238046 67010 238102
rect 67078 238046 67134 238102
rect 67202 238046 67258 238102
rect 67326 238046 67382 238102
rect 66954 237922 67010 237978
rect 67078 237922 67134 237978
rect 67202 237922 67258 237978
rect 67326 237922 67382 237978
rect 66954 220294 67010 220350
rect 67078 220294 67134 220350
rect 67202 220294 67258 220350
rect 67326 220294 67382 220350
rect 66954 220170 67010 220226
rect 67078 220170 67134 220226
rect 67202 220170 67258 220226
rect 67326 220170 67382 220226
rect 66954 220046 67010 220102
rect 67078 220046 67134 220102
rect 67202 220046 67258 220102
rect 67326 220046 67382 220102
rect 66954 219922 67010 219978
rect 67078 219922 67134 219978
rect 67202 219922 67258 219978
rect 67326 219922 67382 219978
rect 66954 202294 67010 202350
rect 67078 202294 67134 202350
rect 67202 202294 67258 202350
rect 67326 202294 67382 202350
rect 66954 202170 67010 202226
rect 67078 202170 67134 202226
rect 67202 202170 67258 202226
rect 67326 202170 67382 202226
rect 66954 202046 67010 202102
rect 67078 202046 67134 202102
rect 67202 202046 67258 202102
rect 67326 202046 67382 202102
rect 66954 201922 67010 201978
rect 67078 201922 67134 201978
rect 67202 201922 67258 201978
rect 67326 201922 67382 201978
rect 66954 184294 67010 184350
rect 67078 184294 67134 184350
rect 67202 184294 67258 184350
rect 67326 184294 67382 184350
rect 66954 184170 67010 184226
rect 67078 184170 67134 184226
rect 67202 184170 67258 184226
rect 67326 184170 67382 184226
rect 66954 184046 67010 184102
rect 67078 184046 67134 184102
rect 67202 184046 67258 184102
rect 67326 184046 67382 184102
rect 66954 183922 67010 183978
rect 67078 183922 67134 183978
rect 67202 183922 67258 183978
rect 67326 183922 67382 183978
rect 66954 166294 67010 166350
rect 67078 166294 67134 166350
rect 67202 166294 67258 166350
rect 67326 166294 67382 166350
rect 66954 166170 67010 166226
rect 67078 166170 67134 166226
rect 67202 166170 67258 166226
rect 67326 166170 67382 166226
rect 66954 166046 67010 166102
rect 67078 166046 67134 166102
rect 67202 166046 67258 166102
rect 67326 166046 67382 166102
rect 66954 165922 67010 165978
rect 67078 165922 67134 165978
rect 67202 165922 67258 165978
rect 67326 165922 67382 165978
rect 66954 148294 67010 148350
rect 67078 148294 67134 148350
rect 67202 148294 67258 148350
rect 67326 148294 67382 148350
rect 66954 148170 67010 148226
rect 67078 148170 67134 148226
rect 67202 148170 67258 148226
rect 67326 148170 67382 148226
rect 66954 148046 67010 148102
rect 67078 148046 67134 148102
rect 67202 148046 67258 148102
rect 67326 148046 67382 148102
rect 66954 147922 67010 147978
rect 67078 147922 67134 147978
rect 67202 147922 67258 147978
rect 67326 147922 67382 147978
rect 66954 130294 67010 130350
rect 67078 130294 67134 130350
rect 67202 130294 67258 130350
rect 67326 130294 67382 130350
rect 66954 130170 67010 130226
rect 67078 130170 67134 130226
rect 67202 130170 67258 130226
rect 67326 130170 67382 130226
rect 66954 130046 67010 130102
rect 67078 130046 67134 130102
rect 67202 130046 67258 130102
rect 67326 130046 67382 130102
rect 66954 129922 67010 129978
rect 67078 129922 67134 129978
rect 67202 129922 67258 129978
rect 67326 129922 67382 129978
rect 66954 112294 67010 112350
rect 67078 112294 67134 112350
rect 67202 112294 67258 112350
rect 67326 112294 67382 112350
rect 66954 112170 67010 112226
rect 67078 112170 67134 112226
rect 67202 112170 67258 112226
rect 67326 112170 67382 112226
rect 66954 112046 67010 112102
rect 67078 112046 67134 112102
rect 67202 112046 67258 112102
rect 67326 112046 67382 112102
rect 66954 111922 67010 111978
rect 67078 111922 67134 111978
rect 67202 111922 67258 111978
rect 67326 111922 67382 111978
rect 66954 94294 67010 94350
rect 67078 94294 67134 94350
rect 67202 94294 67258 94350
rect 67326 94294 67382 94350
rect 66954 94170 67010 94226
rect 67078 94170 67134 94226
rect 67202 94170 67258 94226
rect 67326 94170 67382 94226
rect 66954 94046 67010 94102
rect 67078 94046 67134 94102
rect 67202 94046 67258 94102
rect 67326 94046 67382 94102
rect 66954 93922 67010 93978
rect 67078 93922 67134 93978
rect 67202 93922 67258 93978
rect 67326 93922 67382 93978
rect 48188 36242 48244 36298
rect 49196 47762 49252 47818
rect 48972 44522 49028 44578
rect 51212 37682 51268 37738
rect 50316 24362 50372 24418
rect 50204 19142 50260 19198
rect 50092 14282 50148 14338
rect 49868 12482 49924 12538
rect 50988 17522 51044 17578
rect 50540 15902 50596 15958
rect 51996 30842 52052 30898
rect 51884 24182 51940 24238
rect 51772 18962 51828 19018
rect 52556 29222 52612 29278
rect 52332 14102 52388 14158
rect 48076 1502 48132 1558
rect 48636 1502 48692 1558
rect 56140 69362 56196 69418
rect 54572 59822 54628 59878
rect 53676 56222 53732 56278
rect 53452 29042 53508 29098
rect 53340 24542 53396 24598
rect 53228 8882 53284 8938
rect 54124 41102 54180 41158
rect 53676 7622 53732 7678
rect 53900 20582 53956 20638
rect 53788 5282 53844 5338
rect 52780 1322 52836 1378
rect 53452 962 53508 1018
rect 54348 32462 54404 32518
rect 55692 42722 55748 42778
rect 55468 20402 55524 20458
rect 55244 17342 55300 17398
rect 55356 13922 55412 13978
rect 56140 3482 56196 3538
rect 57036 51362 57092 51418
rect 56364 13382 56420 13438
rect 56700 18782 56756 18838
rect 56924 15722 56980 15778
rect 57036 6722 57092 6778
rect 57260 10862 57316 10918
rect 56588 2942 56644 2998
rect 57708 54602 57764 54658
rect 57932 7262 57988 7318
rect 56252 1502 56308 1558
rect 58380 37502 58436 37558
rect 58716 61082 58772 61138
rect 59500 47582 59556 47638
rect 59276 40922 59332 40978
rect 58940 3662 58996 3718
rect 60172 36062 60228 36118
rect 59724 7622 59780 7678
rect 61068 52802 61124 52858
rect 60844 32282 60900 32338
rect 61852 37322 61908 37378
rect 61740 35882 61796 35938
rect 61292 25802 61348 25858
rect 58044 1142 58100 1198
rect 65212 70622 65268 70678
rect 62598 64294 62654 64350
rect 62722 64294 62778 64350
rect 62598 64170 62654 64226
rect 62722 64170 62778 64226
rect 62598 64046 62654 64102
rect 62722 64046 62778 64102
rect 62598 63922 62654 63978
rect 62722 63922 62778 63978
rect 63196 62882 63252 62938
rect 62598 46294 62654 46350
rect 62722 46294 62778 46350
rect 62598 46170 62654 46226
rect 62722 46170 62778 46226
rect 62598 46046 62654 46102
rect 62722 46046 62778 46102
rect 62598 45922 62654 45978
rect 62722 45922 62778 45978
rect 62598 28294 62654 28350
rect 62722 28294 62778 28350
rect 62598 28170 62654 28226
rect 62722 28170 62778 28226
rect 62598 28046 62654 28102
rect 62722 28046 62778 28102
rect 62598 27922 62654 27978
rect 62722 27922 62778 27978
rect 62598 10294 62654 10350
rect 62722 10294 62778 10350
rect 62598 10170 62654 10226
rect 62722 10170 62778 10226
rect 62598 10046 62654 10102
rect 62722 10046 62778 10102
rect 62598 9922 62654 9978
rect 62722 9922 62778 9978
rect 62972 6722 63028 6778
rect 61516 1502 61572 1558
rect 63644 60002 63700 60058
rect 63532 44702 63588 44758
rect 63420 18602 63476 18658
rect 63308 13742 63364 13798
rect 64428 49562 64484 49618
rect 63980 34442 64036 34498
rect 63756 7082 63812 7138
rect 64204 15542 64260 15598
rect 65100 39482 65156 39538
rect 64876 5642 64932 5698
rect 64764 5462 64820 5518
rect 65212 6542 65268 6598
rect 70674 598116 70730 598172
rect 70798 598116 70854 598172
rect 70922 598116 70978 598172
rect 71046 598116 71102 598172
rect 70674 597992 70730 598048
rect 70798 597992 70854 598048
rect 70922 597992 70978 598048
rect 71046 597992 71102 598048
rect 70674 597868 70730 597924
rect 70798 597868 70854 597924
rect 70922 597868 70978 597924
rect 71046 597868 71102 597924
rect 70674 597744 70730 597800
rect 70798 597744 70854 597800
rect 70922 597744 70978 597800
rect 71046 597744 71102 597800
rect 70674 586294 70730 586350
rect 70798 586294 70854 586350
rect 70922 586294 70978 586350
rect 71046 586294 71102 586350
rect 70674 586170 70730 586226
rect 70798 586170 70854 586226
rect 70922 586170 70978 586226
rect 71046 586170 71102 586226
rect 70674 586046 70730 586102
rect 70798 586046 70854 586102
rect 70922 586046 70978 586102
rect 71046 586046 71102 586102
rect 70674 585922 70730 585978
rect 70798 585922 70854 585978
rect 70922 585922 70978 585978
rect 71046 585922 71102 585978
rect 70674 568294 70730 568350
rect 70798 568294 70854 568350
rect 70922 568294 70978 568350
rect 71046 568294 71102 568350
rect 70674 568170 70730 568226
rect 70798 568170 70854 568226
rect 70922 568170 70978 568226
rect 71046 568170 71102 568226
rect 70674 568046 70730 568102
rect 70798 568046 70854 568102
rect 70922 568046 70978 568102
rect 71046 568046 71102 568102
rect 70674 567922 70730 567978
rect 70798 567922 70854 567978
rect 70922 567922 70978 567978
rect 71046 567922 71102 567978
rect 70674 550294 70730 550350
rect 70798 550294 70854 550350
rect 70922 550294 70978 550350
rect 71046 550294 71102 550350
rect 70674 550170 70730 550226
rect 70798 550170 70854 550226
rect 70922 550170 70978 550226
rect 71046 550170 71102 550226
rect 70674 550046 70730 550102
rect 70798 550046 70854 550102
rect 70922 550046 70978 550102
rect 71046 550046 71102 550102
rect 70674 549922 70730 549978
rect 70798 549922 70854 549978
rect 70922 549922 70978 549978
rect 71046 549922 71102 549978
rect 70674 532294 70730 532350
rect 70798 532294 70854 532350
rect 70922 532294 70978 532350
rect 71046 532294 71102 532350
rect 70674 532170 70730 532226
rect 70798 532170 70854 532226
rect 70922 532170 70978 532226
rect 71046 532170 71102 532226
rect 70674 532046 70730 532102
rect 70798 532046 70854 532102
rect 70922 532046 70978 532102
rect 71046 532046 71102 532102
rect 70674 531922 70730 531978
rect 70798 531922 70854 531978
rect 70922 531922 70978 531978
rect 71046 531922 71102 531978
rect 70674 514294 70730 514350
rect 70798 514294 70854 514350
rect 70922 514294 70978 514350
rect 71046 514294 71102 514350
rect 70674 514170 70730 514226
rect 70798 514170 70854 514226
rect 70922 514170 70978 514226
rect 71046 514170 71102 514226
rect 70674 514046 70730 514102
rect 70798 514046 70854 514102
rect 70922 514046 70978 514102
rect 71046 514046 71102 514102
rect 70674 513922 70730 513978
rect 70798 513922 70854 513978
rect 70922 513922 70978 513978
rect 71046 513922 71102 513978
rect 70674 496294 70730 496350
rect 70798 496294 70854 496350
rect 70922 496294 70978 496350
rect 71046 496294 71102 496350
rect 70674 496170 70730 496226
rect 70798 496170 70854 496226
rect 70922 496170 70978 496226
rect 71046 496170 71102 496226
rect 70674 496046 70730 496102
rect 70798 496046 70854 496102
rect 70922 496046 70978 496102
rect 71046 496046 71102 496102
rect 70674 495922 70730 495978
rect 70798 495922 70854 495978
rect 70922 495922 70978 495978
rect 71046 495922 71102 495978
rect 70674 478294 70730 478350
rect 70798 478294 70854 478350
rect 70922 478294 70978 478350
rect 71046 478294 71102 478350
rect 70674 478170 70730 478226
rect 70798 478170 70854 478226
rect 70922 478170 70978 478226
rect 71046 478170 71102 478226
rect 70674 478046 70730 478102
rect 70798 478046 70854 478102
rect 70922 478046 70978 478102
rect 71046 478046 71102 478102
rect 70674 477922 70730 477978
rect 70798 477922 70854 477978
rect 70922 477922 70978 477978
rect 71046 477922 71102 477978
rect 70674 460294 70730 460350
rect 70798 460294 70854 460350
rect 70922 460294 70978 460350
rect 71046 460294 71102 460350
rect 70674 460170 70730 460226
rect 70798 460170 70854 460226
rect 70922 460170 70978 460226
rect 71046 460170 71102 460226
rect 70674 460046 70730 460102
rect 70798 460046 70854 460102
rect 70922 460046 70978 460102
rect 71046 460046 71102 460102
rect 70674 459922 70730 459978
rect 70798 459922 70854 459978
rect 70922 459922 70978 459978
rect 71046 459922 71102 459978
rect 97674 597156 97730 597212
rect 97798 597156 97854 597212
rect 97922 597156 97978 597212
rect 98046 597156 98102 597212
rect 97674 597032 97730 597088
rect 97798 597032 97854 597088
rect 97922 597032 97978 597088
rect 98046 597032 98102 597088
rect 97674 596908 97730 596964
rect 97798 596908 97854 596964
rect 97922 596908 97978 596964
rect 98046 596908 98102 596964
rect 97674 596784 97730 596840
rect 97798 596784 97854 596840
rect 97922 596784 97978 596840
rect 98046 596784 98102 596840
rect 101394 598116 101450 598172
rect 101518 598116 101574 598172
rect 101642 598116 101698 598172
rect 101766 598116 101822 598172
rect 101394 597992 101450 598048
rect 101518 597992 101574 598048
rect 101642 597992 101698 598048
rect 101766 597992 101822 598048
rect 101394 597868 101450 597924
rect 101518 597868 101574 597924
rect 101642 597868 101698 597924
rect 101766 597868 101822 597924
rect 101394 597744 101450 597800
rect 101518 597744 101574 597800
rect 101642 597744 101698 597800
rect 101766 597744 101822 597800
rect 97674 580294 97730 580350
rect 97798 580294 97854 580350
rect 97922 580294 97978 580350
rect 98046 580294 98102 580350
rect 97674 580170 97730 580226
rect 97798 580170 97854 580226
rect 97922 580170 97978 580226
rect 98046 580170 98102 580226
rect 97674 580046 97730 580102
rect 97798 580046 97854 580102
rect 97922 580046 97978 580102
rect 98046 580046 98102 580102
rect 97674 579922 97730 579978
rect 97798 579922 97854 579978
rect 97922 579922 97978 579978
rect 98046 579922 98102 579978
rect 97674 562294 97730 562350
rect 97798 562294 97854 562350
rect 97922 562294 97978 562350
rect 98046 562294 98102 562350
rect 97674 562170 97730 562226
rect 97798 562170 97854 562226
rect 97922 562170 97978 562226
rect 98046 562170 98102 562226
rect 97674 562046 97730 562102
rect 97798 562046 97854 562102
rect 97922 562046 97978 562102
rect 98046 562046 98102 562102
rect 97674 561922 97730 561978
rect 97798 561922 97854 561978
rect 97922 561922 97978 561978
rect 98046 561922 98102 561978
rect 97674 544294 97730 544350
rect 97798 544294 97854 544350
rect 97922 544294 97978 544350
rect 98046 544294 98102 544350
rect 97674 544170 97730 544226
rect 97798 544170 97854 544226
rect 97922 544170 97978 544226
rect 98046 544170 98102 544226
rect 97674 544046 97730 544102
rect 97798 544046 97854 544102
rect 97922 544046 97978 544102
rect 98046 544046 98102 544102
rect 97674 543922 97730 543978
rect 97798 543922 97854 543978
rect 97922 543922 97978 543978
rect 98046 543922 98102 543978
rect 97674 526294 97730 526350
rect 97798 526294 97854 526350
rect 97922 526294 97978 526350
rect 98046 526294 98102 526350
rect 97674 526170 97730 526226
rect 97798 526170 97854 526226
rect 97922 526170 97978 526226
rect 98046 526170 98102 526226
rect 97674 526046 97730 526102
rect 97798 526046 97854 526102
rect 97922 526046 97978 526102
rect 98046 526046 98102 526102
rect 97674 525922 97730 525978
rect 97798 525922 97854 525978
rect 97922 525922 97978 525978
rect 98046 525922 98102 525978
rect 97674 508294 97730 508350
rect 97798 508294 97854 508350
rect 97922 508294 97978 508350
rect 98046 508294 98102 508350
rect 97674 508170 97730 508226
rect 97798 508170 97854 508226
rect 97922 508170 97978 508226
rect 98046 508170 98102 508226
rect 97674 508046 97730 508102
rect 97798 508046 97854 508102
rect 97922 508046 97978 508102
rect 98046 508046 98102 508102
rect 97674 507922 97730 507978
rect 97798 507922 97854 507978
rect 97922 507922 97978 507978
rect 98046 507922 98102 507978
rect 97674 490294 97730 490350
rect 97798 490294 97854 490350
rect 97922 490294 97978 490350
rect 98046 490294 98102 490350
rect 97674 490170 97730 490226
rect 97798 490170 97854 490226
rect 97922 490170 97978 490226
rect 98046 490170 98102 490226
rect 97674 490046 97730 490102
rect 97798 490046 97854 490102
rect 97922 490046 97978 490102
rect 98046 490046 98102 490102
rect 97674 489922 97730 489978
rect 97798 489922 97854 489978
rect 97922 489922 97978 489978
rect 98046 489922 98102 489978
rect 97674 472294 97730 472350
rect 97798 472294 97854 472350
rect 97922 472294 97978 472350
rect 98046 472294 98102 472350
rect 97674 472170 97730 472226
rect 97798 472170 97854 472226
rect 97922 472170 97978 472226
rect 98046 472170 98102 472226
rect 97674 472046 97730 472102
rect 97798 472046 97854 472102
rect 97922 472046 97978 472102
rect 98046 472046 98102 472102
rect 97674 471922 97730 471978
rect 97798 471922 97854 471978
rect 97922 471922 97978 471978
rect 98046 471922 98102 471978
rect 97674 454294 97730 454350
rect 97798 454294 97854 454350
rect 97922 454294 97978 454350
rect 98046 454294 98102 454350
rect 97674 454170 97730 454226
rect 97798 454170 97854 454226
rect 97922 454170 97978 454226
rect 98046 454170 98102 454226
rect 97674 454046 97730 454102
rect 97798 454046 97854 454102
rect 97922 454046 97978 454102
rect 98046 454046 98102 454102
rect 97674 453922 97730 453978
rect 97798 453922 97854 453978
rect 97922 453922 97978 453978
rect 98046 453922 98102 453978
rect 70674 442294 70730 442350
rect 70798 442294 70854 442350
rect 70922 442294 70978 442350
rect 71046 442294 71102 442350
rect 70674 442170 70730 442226
rect 70798 442170 70854 442226
rect 70922 442170 70978 442226
rect 71046 442170 71102 442226
rect 70674 442046 70730 442102
rect 70798 442046 70854 442102
rect 70922 442046 70978 442102
rect 71046 442046 71102 442102
rect 70674 441922 70730 441978
rect 70798 441922 70854 441978
rect 70922 441922 70978 441978
rect 71046 441922 71102 441978
rect 70674 424294 70730 424350
rect 70798 424294 70854 424350
rect 70922 424294 70978 424350
rect 71046 424294 71102 424350
rect 70674 424170 70730 424226
rect 70798 424170 70854 424226
rect 70922 424170 70978 424226
rect 71046 424170 71102 424226
rect 70674 424046 70730 424102
rect 70798 424046 70854 424102
rect 70922 424046 70978 424102
rect 71046 424046 71102 424102
rect 70674 423922 70730 423978
rect 70798 423922 70854 423978
rect 70922 423922 70978 423978
rect 71046 423922 71102 423978
rect 70674 406294 70730 406350
rect 70798 406294 70854 406350
rect 70922 406294 70978 406350
rect 71046 406294 71102 406350
rect 70674 406170 70730 406226
rect 70798 406170 70854 406226
rect 70922 406170 70978 406226
rect 71046 406170 71102 406226
rect 70674 406046 70730 406102
rect 70798 406046 70854 406102
rect 70922 406046 70978 406102
rect 71046 406046 71102 406102
rect 70674 405922 70730 405978
rect 70798 405922 70854 405978
rect 70922 405922 70978 405978
rect 71046 405922 71102 405978
rect 70674 388294 70730 388350
rect 70798 388294 70854 388350
rect 70922 388294 70978 388350
rect 71046 388294 71102 388350
rect 70674 388170 70730 388226
rect 70798 388170 70854 388226
rect 70922 388170 70978 388226
rect 71046 388170 71102 388226
rect 70674 388046 70730 388102
rect 70798 388046 70854 388102
rect 70922 388046 70978 388102
rect 71046 388046 71102 388102
rect 70674 387922 70730 387978
rect 70798 387922 70854 387978
rect 70922 387922 70978 387978
rect 71046 387922 71102 387978
rect 70674 370294 70730 370350
rect 70798 370294 70854 370350
rect 70922 370294 70978 370350
rect 71046 370294 71102 370350
rect 70674 370170 70730 370226
rect 70798 370170 70854 370226
rect 70922 370170 70978 370226
rect 71046 370170 71102 370226
rect 70674 370046 70730 370102
rect 70798 370046 70854 370102
rect 70922 370046 70978 370102
rect 71046 370046 71102 370102
rect 70674 369922 70730 369978
rect 70798 369922 70854 369978
rect 70922 369922 70978 369978
rect 71046 369922 71102 369978
rect 70674 352294 70730 352350
rect 70798 352294 70854 352350
rect 70922 352294 70978 352350
rect 71046 352294 71102 352350
rect 70674 352170 70730 352226
rect 70798 352170 70854 352226
rect 70922 352170 70978 352226
rect 71046 352170 71102 352226
rect 70674 352046 70730 352102
rect 70798 352046 70854 352102
rect 70922 352046 70978 352102
rect 71046 352046 71102 352102
rect 70674 351922 70730 351978
rect 70798 351922 70854 351978
rect 70922 351922 70978 351978
rect 71046 351922 71102 351978
rect 70674 334294 70730 334350
rect 70798 334294 70854 334350
rect 70922 334294 70978 334350
rect 71046 334294 71102 334350
rect 70674 334170 70730 334226
rect 70798 334170 70854 334226
rect 70922 334170 70978 334226
rect 71046 334170 71102 334226
rect 70674 334046 70730 334102
rect 70798 334046 70854 334102
rect 70922 334046 70978 334102
rect 71046 334046 71102 334102
rect 70674 333922 70730 333978
rect 70798 333922 70854 333978
rect 70922 333922 70978 333978
rect 71046 333922 71102 333978
rect 70674 316294 70730 316350
rect 70798 316294 70854 316350
rect 70922 316294 70978 316350
rect 71046 316294 71102 316350
rect 70674 316170 70730 316226
rect 70798 316170 70854 316226
rect 70922 316170 70978 316226
rect 71046 316170 71102 316226
rect 70674 316046 70730 316102
rect 70798 316046 70854 316102
rect 70922 316046 70978 316102
rect 71046 316046 71102 316102
rect 70674 315922 70730 315978
rect 70798 315922 70854 315978
rect 70922 315922 70978 315978
rect 71046 315922 71102 315978
rect 70674 298294 70730 298350
rect 70798 298294 70854 298350
rect 70922 298294 70978 298350
rect 71046 298294 71102 298350
rect 70674 298170 70730 298226
rect 70798 298170 70854 298226
rect 70922 298170 70978 298226
rect 71046 298170 71102 298226
rect 70674 298046 70730 298102
rect 70798 298046 70854 298102
rect 70922 298046 70978 298102
rect 71046 298046 71102 298102
rect 70674 297922 70730 297978
rect 70798 297922 70854 297978
rect 70922 297922 70978 297978
rect 71046 297922 71102 297978
rect 70674 280294 70730 280350
rect 70798 280294 70854 280350
rect 70922 280294 70978 280350
rect 71046 280294 71102 280350
rect 70674 280170 70730 280226
rect 70798 280170 70854 280226
rect 70922 280170 70978 280226
rect 71046 280170 71102 280226
rect 70674 280046 70730 280102
rect 70798 280046 70854 280102
rect 70922 280046 70978 280102
rect 71046 280046 71102 280102
rect 70674 279922 70730 279978
rect 70798 279922 70854 279978
rect 70922 279922 70978 279978
rect 71046 279922 71102 279978
rect 70674 262294 70730 262350
rect 70798 262294 70854 262350
rect 70922 262294 70978 262350
rect 71046 262294 71102 262350
rect 70674 262170 70730 262226
rect 70798 262170 70854 262226
rect 70922 262170 70978 262226
rect 71046 262170 71102 262226
rect 70674 262046 70730 262102
rect 70798 262046 70854 262102
rect 70922 262046 70978 262102
rect 71046 262046 71102 262102
rect 70674 261922 70730 261978
rect 70798 261922 70854 261978
rect 70922 261922 70978 261978
rect 71046 261922 71102 261978
rect 70674 244294 70730 244350
rect 70798 244294 70854 244350
rect 70922 244294 70978 244350
rect 71046 244294 71102 244350
rect 70674 244170 70730 244226
rect 70798 244170 70854 244226
rect 70922 244170 70978 244226
rect 71046 244170 71102 244226
rect 70674 244046 70730 244102
rect 70798 244046 70854 244102
rect 70922 244046 70978 244102
rect 71046 244046 71102 244102
rect 70674 243922 70730 243978
rect 70798 243922 70854 243978
rect 70922 243922 70978 243978
rect 71046 243922 71102 243978
rect 70674 226294 70730 226350
rect 70798 226294 70854 226350
rect 70922 226294 70978 226350
rect 71046 226294 71102 226350
rect 70674 226170 70730 226226
rect 70798 226170 70854 226226
rect 70922 226170 70978 226226
rect 71046 226170 71102 226226
rect 70674 226046 70730 226102
rect 70798 226046 70854 226102
rect 70922 226046 70978 226102
rect 71046 226046 71102 226102
rect 70674 225922 70730 225978
rect 70798 225922 70854 225978
rect 70922 225922 70978 225978
rect 71046 225922 71102 225978
rect 70674 208294 70730 208350
rect 70798 208294 70854 208350
rect 70922 208294 70978 208350
rect 71046 208294 71102 208350
rect 70674 208170 70730 208226
rect 70798 208170 70854 208226
rect 70922 208170 70978 208226
rect 71046 208170 71102 208226
rect 70674 208046 70730 208102
rect 70798 208046 70854 208102
rect 70922 208046 70978 208102
rect 71046 208046 71102 208102
rect 70674 207922 70730 207978
rect 70798 207922 70854 207978
rect 70922 207922 70978 207978
rect 71046 207922 71102 207978
rect 70674 190294 70730 190350
rect 70798 190294 70854 190350
rect 70922 190294 70978 190350
rect 71046 190294 71102 190350
rect 70674 190170 70730 190226
rect 70798 190170 70854 190226
rect 70922 190170 70978 190226
rect 71046 190170 71102 190226
rect 70674 190046 70730 190102
rect 70798 190046 70854 190102
rect 70922 190046 70978 190102
rect 71046 190046 71102 190102
rect 70674 189922 70730 189978
rect 70798 189922 70854 189978
rect 70922 189922 70978 189978
rect 71046 189922 71102 189978
rect 70674 172294 70730 172350
rect 70798 172294 70854 172350
rect 70922 172294 70978 172350
rect 71046 172294 71102 172350
rect 70674 172170 70730 172226
rect 70798 172170 70854 172226
rect 70922 172170 70978 172226
rect 71046 172170 71102 172226
rect 70674 172046 70730 172102
rect 70798 172046 70854 172102
rect 70922 172046 70978 172102
rect 71046 172046 71102 172102
rect 70674 171922 70730 171978
rect 70798 171922 70854 171978
rect 70922 171922 70978 171978
rect 71046 171922 71102 171978
rect 70674 154294 70730 154350
rect 70798 154294 70854 154350
rect 70922 154294 70978 154350
rect 71046 154294 71102 154350
rect 70674 154170 70730 154226
rect 70798 154170 70854 154226
rect 70922 154170 70978 154226
rect 71046 154170 71102 154226
rect 70674 154046 70730 154102
rect 70798 154046 70854 154102
rect 70922 154046 70978 154102
rect 71046 154046 71102 154102
rect 70674 153922 70730 153978
rect 70798 153922 70854 153978
rect 70922 153922 70978 153978
rect 71046 153922 71102 153978
rect 70674 136294 70730 136350
rect 70798 136294 70854 136350
rect 70922 136294 70978 136350
rect 71046 136294 71102 136350
rect 70674 136170 70730 136226
rect 70798 136170 70854 136226
rect 70922 136170 70978 136226
rect 71046 136170 71102 136226
rect 70674 136046 70730 136102
rect 70798 136046 70854 136102
rect 70922 136046 70978 136102
rect 71046 136046 71102 136102
rect 70674 135922 70730 135978
rect 70798 135922 70854 135978
rect 70922 135922 70978 135978
rect 71046 135922 71102 135978
rect 70674 118294 70730 118350
rect 70798 118294 70854 118350
rect 70922 118294 70978 118350
rect 71046 118294 71102 118350
rect 70674 118170 70730 118226
rect 70798 118170 70854 118226
rect 70922 118170 70978 118226
rect 71046 118170 71102 118226
rect 70674 118046 70730 118102
rect 70798 118046 70854 118102
rect 70922 118046 70978 118102
rect 71046 118046 71102 118102
rect 70674 117922 70730 117978
rect 70798 117922 70854 117978
rect 70922 117922 70978 117978
rect 71046 117922 71102 117978
rect 70674 100294 70730 100350
rect 70798 100294 70854 100350
rect 70922 100294 70978 100350
rect 71046 100294 71102 100350
rect 70674 100170 70730 100226
rect 70798 100170 70854 100226
rect 70922 100170 70978 100226
rect 71046 100170 71102 100226
rect 70674 100046 70730 100102
rect 70798 100046 70854 100102
rect 70922 100046 70978 100102
rect 71046 100046 71102 100102
rect 70674 99922 70730 99978
rect 70798 99922 70854 99978
rect 70922 99922 70978 99978
rect 71046 99922 71102 99978
rect 70674 82294 70730 82350
rect 70798 82294 70854 82350
rect 70922 82294 70978 82350
rect 71046 82294 71102 82350
rect 70674 82170 70730 82226
rect 70798 82170 70854 82226
rect 70922 82170 70978 82226
rect 71046 82170 71102 82226
rect 70674 82046 70730 82102
rect 70798 82046 70854 82102
rect 70922 82046 70978 82102
rect 71046 82046 71102 82102
rect 70674 81922 70730 81978
rect 70798 81922 70854 81978
rect 70922 81922 70978 81978
rect 71046 81922 71102 81978
rect 66954 76294 67010 76350
rect 67078 76294 67134 76350
rect 67202 76294 67258 76350
rect 67326 76294 67382 76350
rect 66954 76170 67010 76226
rect 67078 76170 67134 76226
rect 67202 76170 67258 76226
rect 67326 76170 67382 76226
rect 66954 76046 67010 76102
rect 67078 76046 67134 76102
rect 67202 76046 67258 76102
rect 67326 76046 67382 76102
rect 66954 75922 67010 75978
rect 67078 75922 67134 75978
rect 67202 75922 67258 75978
rect 67326 75922 67382 75978
rect 66556 67562 66612 67618
rect 66444 56402 66500 56458
rect 66332 32642 66388 32698
rect 66220 26162 66276 26218
rect 65996 13382 66052 13438
rect 66954 58294 67010 58350
rect 67078 58294 67134 58350
rect 67202 58294 67258 58350
rect 67326 58294 67382 58350
rect 66954 58170 67010 58226
rect 67078 58170 67134 58226
rect 67202 58170 67258 58226
rect 67326 58170 67382 58226
rect 66954 58046 67010 58102
rect 67078 58046 67134 58102
rect 67202 58046 67258 58102
rect 67326 58046 67382 58102
rect 66954 57922 67010 57978
rect 67078 57922 67134 57978
rect 67202 57922 67258 57978
rect 67326 57922 67382 57978
rect 66954 40294 67010 40350
rect 67078 40294 67134 40350
rect 67202 40294 67258 40350
rect 67326 40294 67382 40350
rect 66954 40170 67010 40226
rect 67078 40170 67134 40226
rect 67202 40170 67258 40226
rect 67326 40170 67382 40226
rect 66954 40046 67010 40102
rect 67078 40046 67134 40102
rect 67202 40046 67258 40102
rect 67326 40046 67382 40102
rect 66954 39922 67010 39978
rect 67078 39922 67134 39978
rect 67202 39922 67258 39978
rect 67326 39922 67382 39978
rect 66954 22294 67010 22350
rect 67078 22294 67134 22350
rect 67202 22294 67258 22350
rect 67326 22294 67382 22350
rect 66954 22170 67010 22226
rect 67078 22170 67134 22226
rect 67202 22170 67258 22226
rect 67326 22170 67382 22226
rect 66954 22046 67010 22102
rect 67078 22046 67134 22102
rect 67202 22046 67258 22102
rect 67326 22046 67382 22102
rect 66954 21922 67010 21978
rect 67078 21922 67134 21978
rect 67202 21922 67258 21978
rect 67326 21922 67382 21978
rect 66954 4294 67010 4350
rect 67078 4294 67134 4350
rect 67202 4294 67258 4350
rect 67326 4294 67382 4350
rect 66954 4170 67010 4226
rect 67078 4170 67134 4226
rect 67202 4170 67258 4226
rect 67326 4170 67382 4226
rect 66954 4046 67010 4102
rect 67078 4046 67134 4102
rect 67202 4046 67258 4102
rect 67326 4046 67382 4102
rect 66954 3922 67010 3978
rect 67078 3922 67134 3978
rect 67202 3922 67258 3978
rect 67326 3922 67382 3978
rect 62412 1322 62468 1378
rect 65772 1142 65828 1198
rect 58156 62 58212 118
rect 39954 -1176 40010 -1120
rect 40078 -1176 40134 -1120
rect 40202 -1176 40258 -1120
rect 40326 -1176 40382 -1120
rect 39954 -1300 40010 -1244
rect 40078 -1300 40134 -1244
rect 40202 -1300 40258 -1244
rect 40326 -1300 40382 -1244
rect 39954 -1424 40010 -1368
rect 40078 -1424 40134 -1368
rect 40202 -1424 40258 -1368
rect 40326 -1424 40382 -1368
rect 39954 -1548 40010 -1492
rect 40078 -1548 40134 -1492
rect 40202 -1548 40258 -1492
rect 40326 -1548 40382 -1492
rect 68684 70802 68740 70858
rect 68572 52622 68628 52678
rect 68460 32102 68516 32158
rect 68348 6542 68404 6598
rect 70140 69002 70196 69058
rect 69468 54782 69524 54838
rect 70028 30302 70084 30358
rect 69916 22742 69972 22798
rect 70674 64294 70730 64350
rect 70798 64294 70854 64350
rect 70922 64294 70978 64350
rect 71046 64294 71102 64350
rect 70674 64170 70730 64226
rect 70798 64170 70854 64226
rect 70922 64170 70978 64226
rect 71046 64170 71102 64226
rect 70674 64046 70730 64102
rect 70798 64046 70854 64102
rect 70922 64046 70978 64102
rect 71046 64046 71102 64102
rect 70674 63922 70730 63978
rect 70798 63922 70854 63978
rect 70922 63922 70978 63978
rect 71046 63922 71102 63978
rect 70674 46294 70730 46350
rect 70798 46294 70854 46350
rect 70922 46294 70978 46350
rect 71046 46294 71102 46350
rect 70674 46170 70730 46226
rect 70798 46170 70854 46226
rect 70922 46170 70978 46226
rect 71046 46170 71102 46226
rect 70674 46046 70730 46102
rect 70798 46046 70854 46102
rect 70922 46046 70978 46102
rect 71046 46046 71102 46102
rect 70674 45922 70730 45978
rect 70798 45922 70854 45978
rect 70922 45922 70978 45978
rect 71046 45922 71102 45978
rect 70674 28294 70730 28350
rect 70798 28294 70854 28350
rect 70922 28294 70978 28350
rect 71046 28294 71102 28350
rect 70674 28170 70730 28226
rect 70798 28170 70854 28226
rect 70922 28170 70978 28226
rect 71046 28170 71102 28226
rect 70674 28046 70730 28102
rect 70798 28046 70854 28102
rect 70922 28046 70978 28102
rect 71046 28046 71102 28102
rect 70674 27922 70730 27978
rect 70798 27922 70854 27978
rect 70922 27922 70978 27978
rect 71046 27922 71102 27978
rect 70674 10294 70730 10350
rect 70798 10294 70854 10350
rect 70922 10294 70978 10350
rect 71046 10294 71102 10350
rect 70674 10170 70730 10226
rect 70798 10170 70854 10226
rect 70922 10170 70978 10226
rect 71046 10170 71102 10226
rect 70674 10046 70730 10102
rect 70798 10046 70854 10102
rect 70922 10046 70978 10102
rect 71046 10046 71102 10102
rect 70674 9922 70730 9978
rect 70798 9922 70854 9978
rect 70922 9922 70978 9978
rect 71046 9922 71102 9978
rect 66954 -216 67010 -160
rect 67078 -216 67134 -160
rect 67202 -216 67258 -160
rect 67326 -216 67382 -160
rect 66954 -340 67010 -284
rect 67078 -340 67134 -284
rect 67202 -340 67258 -284
rect 67326 -340 67382 -284
rect 66954 -464 67010 -408
rect 67078 -464 67134 -408
rect 67202 -464 67258 -408
rect 67326 -464 67382 -408
rect 66954 -588 67010 -532
rect 67078 -588 67134 -532
rect 67202 -588 67258 -532
rect 67326 -588 67382 -532
rect 71596 13382 71652 13438
rect 72044 51542 72100 51598
rect 71932 25082 71988 25138
rect 72940 42362 72996 42418
rect 72940 34442 72996 34498
rect 73052 30302 73108 30358
rect 73164 59642 73220 59698
rect 73052 26882 73108 26938
rect 73724 40742 73780 40798
rect 73164 26162 73220 26218
rect 73612 30482 73668 30538
rect 73052 24542 73108 24598
rect 73500 25982 73556 26038
rect 73164 17162 73220 17218
rect 73948 51182 74004 51238
rect 73948 47762 74004 47818
rect 74844 59462 74900 59518
rect 75292 43802 75348 43858
rect 74956 35702 75012 35758
rect 75180 33902 75236 33958
rect 75516 45602 75572 45658
rect 75516 36242 75572 36298
rect 76412 65402 76468 65458
rect 76412 62522 76468 62578
rect 76076 42182 76132 42238
rect 76412 13382 76468 13438
rect 76636 25082 76692 25138
rect 76860 24002 76916 24058
rect 76748 19322 76804 19378
rect 76972 21662 77028 21718
rect 77958 58294 78014 58350
rect 78082 58294 78138 58350
rect 77958 58170 78014 58226
rect 78082 58170 78138 58226
rect 77958 58046 78014 58102
rect 78082 58046 78138 58102
rect 77958 57922 78014 57978
rect 78082 57922 78138 57978
rect 77958 40294 78014 40350
rect 78082 40294 78138 40350
rect 77958 40170 78014 40226
rect 78082 40170 78138 40226
rect 77958 40046 78014 40102
rect 78082 40046 78138 40102
rect 77958 39922 78014 39978
rect 78082 39922 78138 39978
rect 77644 25082 77700 25138
rect 77308 9062 77364 9118
rect 76300 1502 76356 1558
rect 77958 22294 78014 22350
rect 78082 22294 78138 22350
rect 77958 22170 78014 22226
rect 78082 22170 78138 22226
rect 77958 22046 78014 22102
rect 78082 22046 78138 22102
rect 77958 21922 78014 21978
rect 78082 21922 78138 21978
rect 78428 64682 78484 64738
rect 78428 51362 78484 51418
rect 78540 54962 78596 55018
rect 78316 21662 78372 21718
rect 78428 48662 78484 48718
rect 77980 5282 78036 5338
rect 78652 20222 78708 20278
rect 80108 72602 80164 72658
rect 79884 60362 79940 60418
rect 79772 52982 79828 53038
rect 79884 44702 79940 44758
rect 79996 55862 80052 55918
rect 79884 37142 79940 37198
rect 79996 25082 80052 25138
rect 79996 12122 80052 12178
rect 81228 65762 81284 65818
rect 80556 61262 80612 61318
rect 80556 59822 80612 59878
rect 80556 34262 80612 34318
rect 80556 32642 80612 32698
rect 80780 33722 80836 33778
rect 80556 26162 80612 26218
rect 80444 23822 80500 23878
rect 81564 48662 81620 48718
rect 81676 43982 81732 44038
rect 81564 41282 81620 41338
rect 81676 33902 81732 33958
rect 81676 23642 81732 23698
rect 81900 6722 81956 6778
rect 82796 32642 82852 32698
rect 82908 5462 82964 5518
rect 84588 72422 84644 72478
rect 83132 69182 83188 69238
rect 83356 67742 83412 67798
rect 83132 54962 83188 55018
rect 83244 60902 83300 60958
rect 83132 44342 83188 44398
rect 83356 54782 83412 54838
rect 84140 67382 84196 67438
rect 83804 35522 83860 35578
rect 83244 26162 83300 26218
rect 83692 28862 83748 28918
rect 83244 12302 83300 12358
rect 81564 1502 81620 1558
rect 81788 1502 81844 1558
rect 83580 8522 83636 8578
rect 84700 64862 84756 64918
rect 84700 60002 84756 60058
rect 85932 79262 85988 79318
rect 84924 65942 84980 65998
rect 84924 51542 84980 51598
rect 85484 51002 85540 51058
rect 84924 36962 84980 37018
rect 85036 25442 85092 25498
rect 97674 436294 97730 436350
rect 97798 436294 97854 436350
rect 97922 436294 97978 436350
rect 98046 436294 98102 436350
rect 97674 436170 97730 436226
rect 97798 436170 97854 436226
rect 97922 436170 97978 436226
rect 98046 436170 98102 436226
rect 97674 436046 97730 436102
rect 97798 436046 97854 436102
rect 97922 436046 97978 436102
rect 98046 436046 98102 436102
rect 97674 435922 97730 435978
rect 97798 435922 97854 435978
rect 97922 435922 97978 435978
rect 98046 435922 98102 435978
rect 97674 418294 97730 418350
rect 97798 418294 97854 418350
rect 97922 418294 97978 418350
rect 98046 418294 98102 418350
rect 97674 418170 97730 418226
rect 97798 418170 97854 418226
rect 97922 418170 97978 418226
rect 98046 418170 98102 418226
rect 97674 418046 97730 418102
rect 97798 418046 97854 418102
rect 97922 418046 97978 418102
rect 98046 418046 98102 418102
rect 97674 417922 97730 417978
rect 97798 417922 97854 417978
rect 97922 417922 97978 417978
rect 98046 417922 98102 417978
rect 97674 400294 97730 400350
rect 97798 400294 97854 400350
rect 97922 400294 97978 400350
rect 98046 400294 98102 400350
rect 97674 400170 97730 400226
rect 97798 400170 97854 400226
rect 97922 400170 97978 400226
rect 98046 400170 98102 400226
rect 97674 400046 97730 400102
rect 97798 400046 97854 400102
rect 97922 400046 97978 400102
rect 98046 400046 98102 400102
rect 97674 399922 97730 399978
rect 97798 399922 97854 399978
rect 97922 399922 97978 399978
rect 98046 399922 98102 399978
rect 97674 382294 97730 382350
rect 97798 382294 97854 382350
rect 97922 382294 97978 382350
rect 98046 382294 98102 382350
rect 97674 382170 97730 382226
rect 97798 382170 97854 382226
rect 97922 382170 97978 382226
rect 98046 382170 98102 382226
rect 97674 382046 97730 382102
rect 97798 382046 97854 382102
rect 97922 382046 97978 382102
rect 98046 382046 98102 382102
rect 97674 381922 97730 381978
rect 97798 381922 97854 381978
rect 97922 381922 97978 381978
rect 98046 381922 98102 381978
rect 97674 364294 97730 364350
rect 97798 364294 97854 364350
rect 97922 364294 97978 364350
rect 98046 364294 98102 364350
rect 97674 364170 97730 364226
rect 97798 364170 97854 364226
rect 97922 364170 97978 364226
rect 98046 364170 98102 364226
rect 97674 364046 97730 364102
rect 97798 364046 97854 364102
rect 97922 364046 97978 364102
rect 98046 364046 98102 364102
rect 97674 363922 97730 363978
rect 97798 363922 97854 363978
rect 97922 363922 97978 363978
rect 98046 363922 98102 363978
rect 97674 346294 97730 346350
rect 97798 346294 97854 346350
rect 97922 346294 97978 346350
rect 98046 346294 98102 346350
rect 97674 346170 97730 346226
rect 97798 346170 97854 346226
rect 97922 346170 97978 346226
rect 98046 346170 98102 346226
rect 97674 346046 97730 346102
rect 97798 346046 97854 346102
rect 97922 346046 97978 346102
rect 98046 346046 98102 346102
rect 97674 345922 97730 345978
rect 97798 345922 97854 345978
rect 97922 345922 97978 345978
rect 98046 345922 98102 345978
rect 97674 328294 97730 328350
rect 97798 328294 97854 328350
rect 97922 328294 97978 328350
rect 98046 328294 98102 328350
rect 97674 328170 97730 328226
rect 97798 328170 97854 328226
rect 97922 328170 97978 328226
rect 98046 328170 98102 328226
rect 97674 328046 97730 328102
rect 97798 328046 97854 328102
rect 97922 328046 97978 328102
rect 98046 328046 98102 328102
rect 97674 327922 97730 327978
rect 97798 327922 97854 327978
rect 97922 327922 97978 327978
rect 98046 327922 98102 327978
rect 97674 310294 97730 310350
rect 97798 310294 97854 310350
rect 97922 310294 97978 310350
rect 98046 310294 98102 310350
rect 97674 310170 97730 310226
rect 97798 310170 97854 310226
rect 97922 310170 97978 310226
rect 98046 310170 98102 310226
rect 97674 310046 97730 310102
rect 97798 310046 97854 310102
rect 97922 310046 97978 310102
rect 98046 310046 98102 310102
rect 97674 309922 97730 309978
rect 97798 309922 97854 309978
rect 97922 309922 97978 309978
rect 98046 309922 98102 309978
rect 97674 292294 97730 292350
rect 97798 292294 97854 292350
rect 97922 292294 97978 292350
rect 98046 292294 98102 292350
rect 97674 292170 97730 292226
rect 97798 292170 97854 292226
rect 97922 292170 97978 292226
rect 98046 292170 98102 292226
rect 97674 292046 97730 292102
rect 97798 292046 97854 292102
rect 97922 292046 97978 292102
rect 98046 292046 98102 292102
rect 97674 291922 97730 291978
rect 97798 291922 97854 291978
rect 97922 291922 97978 291978
rect 98046 291922 98102 291978
rect 97674 274294 97730 274350
rect 97798 274294 97854 274350
rect 97922 274294 97978 274350
rect 98046 274294 98102 274350
rect 97674 274170 97730 274226
rect 97798 274170 97854 274226
rect 97922 274170 97978 274226
rect 98046 274170 98102 274226
rect 97674 274046 97730 274102
rect 97798 274046 97854 274102
rect 97922 274046 97978 274102
rect 98046 274046 98102 274102
rect 97674 273922 97730 273978
rect 97798 273922 97854 273978
rect 97922 273922 97978 273978
rect 98046 273922 98102 273978
rect 97674 256294 97730 256350
rect 97798 256294 97854 256350
rect 97922 256294 97978 256350
rect 98046 256294 98102 256350
rect 97674 256170 97730 256226
rect 97798 256170 97854 256226
rect 97922 256170 97978 256226
rect 98046 256170 98102 256226
rect 97674 256046 97730 256102
rect 97798 256046 97854 256102
rect 97922 256046 97978 256102
rect 98046 256046 98102 256102
rect 97674 255922 97730 255978
rect 97798 255922 97854 255978
rect 97922 255922 97978 255978
rect 98046 255922 98102 255978
rect 97674 238294 97730 238350
rect 97798 238294 97854 238350
rect 97922 238294 97978 238350
rect 98046 238294 98102 238350
rect 97674 238170 97730 238226
rect 97798 238170 97854 238226
rect 97922 238170 97978 238226
rect 98046 238170 98102 238226
rect 97674 238046 97730 238102
rect 97798 238046 97854 238102
rect 97922 238046 97978 238102
rect 98046 238046 98102 238102
rect 97674 237922 97730 237978
rect 97798 237922 97854 237978
rect 97922 237922 97978 237978
rect 98046 237922 98102 237978
rect 97674 220294 97730 220350
rect 97798 220294 97854 220350
rect 97922 220294 97978 220350
rect 98046 220294 98102 220350
rect 97674 220170 97730 220226
rect 97798 220170 97854 220226
rect 97922 220170 97978 220226
rect 98046 220170 98102 220226
rect 97674 220046 97730 220102
rect 97798 220046 97854 220102
rect 97922 220046 97978 220102
rect 98046 220046 98102 220102
rect 97674 219922 97730 219978
rect 97798 219922 97854 219978
rect 97922 219922 97978 219978
rect 98046 219922 98102 219978
rect 97674 202294 97730 202350
rect 97798 202294 97854 202350
rect 97922 202294 97978 202350
rect 98046 202294 98102 202350
rect 97674 202170 97730 202226
rect 97798 202170 97854 202226
rect 97922 202170 97978 202226
rect 98046 202170 98102 202226
rect 97674 202046 97730 202102
rect 97798 202046 97854 202102
rect 97922 202046 97978 202102
rect 98046 202046 98102 202102
rect 97674 201922 97730 201978
rect 97798 201922 97854 201978
rect 97922 201922 97978 201978
rect 98046 201922 98102 201978
rect 97674 184294 97730 184350
rect 97798 184294 97854 184350
rect 97922 184294 97978 184350
rect 98046 184294 98102 184350
rect 97674 184170 97730 184226
rect 97798 184170 97854 184226
rect 97922 184170 97978 184226
rect 98046 184170 98102 184226
rect 97674 184046 97730 184102
rect 97798 184046 97854 184102
rect 97922 184046 97978 184102
rect 98046 184046 98102 184102
rect 97674 183922 97730 183978
rect 97798 183922 97854 183978
rect 97922 183922 97978 183978
rect 98046 183922 98102 183978
rect 97674 166294 97730 166350
rect 97798 166294 97854 166350
rect 97922 166294 97978 166350
rect 98046 166294 98102 166350
rect 97674 166170 97730 166226
rect 97798 166170 97854 166226
rect 97922 166170 97978 166226
rect 98046 166170 98102 166226
rect 97674 166046 97730 166102
rect 97798 166046 97854 166102
rect 97922 166046 97978 166102
rect 98046 166046 98102 166102
rect 97674 165922 97730 165978
rect 97798 165922 97854 165978
rect 97922 165922 97978 165978
rect 98046 165922 98102 165978
rect 97674 148294 97730 148350
rect 97798 148294 97854 148350
rect 97922 148294 97978 148350
rect 98046 148294 98102 148350
rect 97674 148170 97730 148226
rect 97798 148170 97854 148226
rect 97922 148170 97978 148226
rect 98046 148170 98102 148226
rect 97674 148046 97730 148102
rect 97798 148046 97854 148102
rect 97922 148046 97978 148102
rect 98046 148046 98102 148102
rect 97674 147922 97730 147978
rect 97798 147922 97854 147978
rect 97922 147922 97978 147978
rect 98046 147922 98102 147978
rect 97674 130294 97730 130350
rect 97798 130294 97854 130350
rect 97922 130294 97978 130350
rect 98046 130294 98102 130350
rect 97674 130170 97730 130226
rect 97798 130170 97854 130226
rect 97922 130170 97978 130226
rect 98046 130170 98102 130226
rect 97674 130046 97730 130102
rect 97798 130046 97854 130102
rect 97922 130046 97978 130102
rect 98046 130046 98102 130102
rect 97674 129922 97730 129978
rect 97798 129922 97854 129978
rect 97922 129922 97978 129978
rect 98046 129922 98102 129978
rect 97674 112294 97730 112350
rect 97798 112294 97854 112350
rect 97922 112294 97978 112350
rect 98046 112294 98102 112350
rect 97674 112170 97730 112226
rect 97798 112170 97854 112226
rect 97922 112170 97978 112226
rect 98046 112170 98102 112226
rect 97674 112046 97730 112102
rect 97798 112046 97854 112102
rect 97922 112046 97978 112102
rect 98046 112046 98102 112102
rect 97674 111922 97730 111978
rect 97798 111922 97854 111978
rect 97922 111922 97978 111978
rect 98046 111922 98102 111978
rect 97674 94294 97730 94350
rect 97798 94294 97854 94350
rect 97922 94294 97978 94350
rect 98046 94294 98102 94350
rect 97674 94170 97730 94226
rect 97798 94170 97854 94226
rect 97922 94170 97978 94226
rect 98046 94170 98102 94226
rect 97674 94046 97730 94102
rect 97798 94046 97854 94102
rect 97922 94046 97978 94102
rect 98046 94046 98102 94102
rect 97674 93922 97730 93978
rect 97798 93922 97854 93978
rect 97922 93922 97978 93978
rect 98046 93922 98102 93978
rect 89740 79082 89796 79138
rect 86492 63602 86548 63658
rect 86156 47402 86212 47458
rect 87276 74042 87332 74098
rect 87164 59282 87220 59338
rect 87052 54422 87108 54478
rect 86940 22562 86996 22618
rect 87388 66122 87444 66178
rect 87388 62882 87444 62938
rect 87836 28682 87892 28738
rect 87836 25442 87892 25498
rect 87500 16802 87556 16858
rect 87388 6002 87444 6058
rect 87836 11762 87892 11818
rect 88956 72242 89012 72298
rect 88284 70982 88340 71038
rect 88844 62342 88900 62398
rect 88284 49562 88340 49618
rect 88732 52442 88788 52498
rect 88172 49022 88228 49078
rect 89516 59102 89572 59158
rect 89292 50822 89348 50878
rect 89068 13562 89124 13618
rect 92316 77282 92372 77338
rect 89852 71162 89908 71218
rect 89852 60362 89908 60418
rect 90636 60722 90692 60778
rect 90412 54242 90468 54298
rect 89852 25622 89908 25678
rect 89852 19322 89908 19378
rect 89852 16982 89908 17038
rect 89404 2762 89460 2818
rect 90860 47222 90916 47278
rect 90748 45422 90804 45478
rect 90748 42722 90804 42778
rect 90748 34082 90804 34138
rect 90748 28682 90804 28738
rect 90748 8522 90804 8578
rect 91308 38762 91364 38818
rect 90972 11042 91028 11098
rect 89852 1502 89908 1558
rect 91644 67922 91700 67978
rect 91644 56222 91700 56278
rect 91756 66302 91812 66358
rect 91644 56042 91700 56098
rect 91756 52802 91812 52858
rect 91644 39482 91700 39538
rect 92204 30302 92260 30358
rect 92092 28682 92148 28738
rect 128394 597156 128450 597212
rect 128518 597156 128574 597212
rect 128642 597156 128698 597212
rect 128766 597156 128822 597212
rect 128394 597032 128450 597088
rect 128518 597032 128574 597088
rect 128642 597032 128698 597088
rect 128766 597032 128822 597088
rect 128394 596908 128450 596964
rect 128518 596908 128574 596964
rect 128642 596908 128698 596964
rect 128766 596908 128822 596964
rect 128394 596784 128450 596840
rect 128518 596784 128574 596840
rect 128642 596784 128698 596840
rect 128766 596784 128822 596840
rect 101394 586294 101450 586350
rect 101518 586294 101574 586350
rect 101642 586294 101698 586350
rect 101766 586294 101822 586350
rect 101394 586170 101450 586226
rect 101518 586170 101574 586226
rect 101642 586170 101698 586226
rect 101766 586170 101822 586226
rect 101394 586046 101450 586102
rect 101518 586046 101574 586102
rect 101642 586046 101698 586102
rect 101766 586046 101822 586102
rect 101394 585922 101450 585978
rect 101518 585922 101574 585978
rect 101642 585922 101698 585978
rect 101766 585922 101822 585978
rect 99148 79982 99204 80038
rect 101394 568294 101450 568350
rect 101518 568294 101574 568350
rect 101642 568294 101698 568350
rect 101766 568294 101822 568350
rect 101394 568170 101450 568226
rect 101518 568170 101574 568226
rect 101642 568170 101698 568226
rect 101766 568170 101822 568226
rect 101394 568046 101450 568102
rect 101518 568046 101574 568102
rect 101642 568046 101698 568102
rect 101766 568046 101822 568102
rect 101394 567922 101450 567978
rect 101518 567922 101574 567978
rect 101642 567922 101698 567978
rect 101766 567922 101822 567978
rect 101394 550294 101450 550350
rect 101518 550294 101574 550350
rect 101642 550294 101698 550350
rect 101766 550294 101822 550350
rect 101394 550170 101450 550226
rect 101518 550170 101574 550226
rect 101642 550170 101698 550226
rect 101766 550170 101822 550226
rect 101394 550046 101450 550102
rect 101518 550046 101574 550102
rect 101642 550046 101698 550102
rect 101766 550046 101822 550102
rect 101394 549922 101450 549978
rect 101518 549922 101574 549978
rect 101642 549922 101698 549978
rect 101766 549922 101822 549978
rect 101394 532294 101450 532350
rect 101518 532294 101574 532350
rect 101642 532294 101698 532350
rect 101766 532294 101822 532350
rect 101394 532170 101450 532226
rect 101518 532170 101574 532226
rect 101642 532170 101698 532226
rect 101766 532170 101822 532226
rect 101394 532046 101450 532102
rect 101518 532046 101574 532102
rect 101642 532046 101698 532102
rect 101766 532046 101822 532102
rect 101394 531922 101450 531978
rect 101518 531922 101574 531978
rect 101642 531922 101698 531978
rect 101766 531922 101822 531978
rect 101394 514294 101450 514350
rect 101518 514294 101574 514350
rect 101642 514294 101698 514350
rect 101766 514294 101822 514350
rect 101394 514170 101450 514226
rect 101518 514170 101574 514226
rect 101642 514170 101698 514226
rect 101766 514170 101822 514226
rect 101394 514046 101450 514102
rect 101518 514046 101574 514102
rect 101642 514046 101698 514102
rect 101766 514046 101822 514102
rect 101394 513922 101450 513978
rect 101518 513922 101574 513978
rect 101642 513922 101698 513978
rect 101766 513922 101822 513978
rect 101394 496294 101450 496350
rect 101518 496294 101574 496350
rect 101642 496294 101698 496350
rect 101766 496294 101822 496350
rect 101394 496170 101450 496226
rect 101518 496170 101574 496226
rect 101642 496170 101698 496226
rect 101766 496170 101822 496226
rect 101394 496046 101450 496102
rect 101518 496046 101574 496102
rect 101642 496046 101698 496102
rect 101766 496046 101822 496102
rect 101394 495922 101450 495978
rect 101518 495922 101574 495978
rect 101642 495922 101698 495978
rect 101766 495922 101822 495978
rect 101394 478294 101450 478350
rect 101518 478294 101574 478350
rect 101642 478294 101698 478350
rect 101766 478294 101822 478350
rect 101394 478170 101450 478226
rect 101518 478170 101574 478226
rect 101642 478170 101698 478226
rect 101766 478170 101822 478226
rect 101394 478046 101450 478102
rect 101518 478046 101574 478102
rect 101642 478046 101698 478102
rect 101766 478046 101822 478102
rect 101394 477922 101450 477978
rect 101518 477922 101574 477978
rect 101642 477922 101698 477978
rect 101766 477922 101822 477978
rect 101394 460294 101450 460350
rect 101518 460294 101574 460350
rect 101642 460294 101698 460350
rect 101766 460294 101822 460350
rect 101394 460170 101450 460226
rect 101518 460170 101574 460226
rect 101642 460170 101698 460226
rect 101766 460170 101822 460226
rect 101394 460046 101450 460102
rect 101518 460046 101574 460102
rect 101642 460046 101698 460102
rect 101766 460046 101822 460102
rect 101394 459922 101450 459978
rect 101518 459922 101574 459978
rect 101642 459922 101698 459978
rect 101766 459922 101822 459978
rect 101394 442294 101450 442350
rect 101518 442294 101574 442350
rect 101642 442294 101698 442350
rect 101766 442294 101822 442350
rect 101394 442170 101450 442226
rect 101518 442170 101574 442226
rect 101642 442170 101698 442226
rect 101766 442170 101822 442226
rect 101394 442046 101450 442102
rect 101518 442046 101574 442102
rect 101642 442046 101698 442102
rect 101766 442046 101822 442102
rect 101394 441922 101450 441978
rect 101518 441922 101574 441978
rect 101642 441922 101698 441978
rect 101766 441922 101822 441978
rect 101394 424294 101450 424350
rect 101518 424294 101574 424350
rect 101642 424294 101698 424350
rect 101766 424294 101822 424350
rect 101394 424170 101450 424226
rect 101518 424170 101574 424226
rect 101642 424170 101698 424226
rect 101766 424170 101822 424226
rect 101394 424046 101450 424102
rect 101518 424046 101574 424102
rect 101642 424046 101698 424102
rect 101766 424046 101822 424102
rect 101394 423922 101450 423978
rect 101518 423922 101574 423978
rect 101642 423922 101698 423978
rect 101766 423922 101822 423978
rect 101394 406294 101450 406350
rect 101518 406294 101574 406350
rect 101642 406294 101698 406350
rect 101766 406294 101822 406350
rect 101394 406170 101450 406226
rect 101518 406170 101574 406226
rect 101642 406170 101698 406226
rect 101766 406170 101822 406226
rect 101394 406046 101450 406102
rect 101518 406046 101574 406102
rect 101642 406046 101698 406102
rect 101766 406046 101822 406102
rect 101394 405922 101450 405978
rect 101518 405922 101574 405978
rect 101642 405922 101698 405978
rect 101766 405922 101822 405978
rect 101394 388294 101450 388350
rect 101518 388294 101574 388350
rect 101642 388294 101698 388350
rect 101766 388294 101822 388350
rect 101394 388170 101450 388226
rect 101518 388170 101574 388226
rect 101642 388170 101698 388226
rect 101766 388170 101822 388226
rect 101394 388046 101450 388102
rect 101518 388046 101574 388102
rect 101642 388046 101698 388102
rect 101766 388046 101822 388102
rect 101394 387922 101450 387978
rect 101518 387922 101574 387978
rect 101642 387922 101698 387978
rect 101766 387922 101822 387978
rect 101394 370294 101450 370350
rect 101518 370294 101574 370350
rect 101642 370294 101698 370350
rect 101766 370294 101822 370350
rect 101394 370170 101450 370226
rect 101518 370170 101574 370226
rect 101642 370170 101698 370226
rect 101766 370170 101822 370226
rect 101394 370046 101450 370102
rect 101518 370046 101574 370102
rect 101642 370046 101698 370102
rect 101766 370046 101822 370102
rect 101394 369922 101450 369978
rect 101518 369922 101574 369978
rect 101642 369922 101698 369978
rect 101766 369922 101822 369978
rect 101394 352294 101450 352350
rect 101518 352294 101574 352350
rect 101642 352294 101698 352350
rect 101766 352294 101822 352350
rect 101394 352170 101450 352226
rect 101518 352170 101574 352226
rect 101642 352170 101698 352226
rect 101766 352170 101822 352226
rect 101394 352046 101450 352102
rect 101518 352046 101574 352102
rect 101642 352046 101698 352102
rect 101766 352046 101822 352102
rect 101394 351922 101450 351978
rect 101518 351922 101574 351978
rect 101642 351922 101698 351978
rect 101766 351922 101822 351978
rect 101394 334294 101450 334350
rect 101518 334294 101574 334350
rect 101642 334294 101698 334350
rect 101766 334294 101822 334350
rect 101394 334170 101450 334226
rect 101518 334170 101574 334226
rect 101642 334170 101698 334226
rect 101766 334170 101822 334226
rect 101394 334046 101450 334102
rect 101518 334046 101574 334102
rect 101642 334046 101698 334102
rect 101766 334046 101822 334102
rect 101394 333922 101450 333978
rect 101518 333922 101574 333978
rect 101642 333922 101698 333978
rect 101766 333922 101822 333978
rect 101394 316294 101450 316350
rect 101518 316294 101574 316350
rect 101642 316294 101698 316350
rect 101766 316294 101822 316350
rect 101394 316170 101450 316226
rect 101518 316170 101574 316226
rect 101642 316170 101698 316226
rect 101766 316170 101822 316226
rect 101394 316046 101450 316102
rect 101518 316046 101574 316102
rect 101642 316046 101698 316102
rect 101766 316046 101822 316102
rect 101394 315922 101450 315978
rect 101518 315922 101574 315978
rect 101642 315922 101698 315978
rect 101766 315922 101822 315978
rect 101394 298294 101450 298350
rect 101518 298294 101574 298350
rect 101642 298294 101698 298350
rect 101766 298294 101822 298350
rect 101394 298170 101450 298226
rect 101518 298170 101574 298226
rect 101642 298170 101698 298226
rect 101766 298170 101822 298226
rect 101394 298046 101450 298102
rect 101518 298046 101574 298102
rect 101642 298046 101698 298102
rect 101766 298046 101822 298102
rect 101394 297922 101450 297978
rect 101518 297922 101574 297978
rect 101642 297922 101698 297978
rect 101766 297922 101822 297978
rect 101394 280294 101450 280350
rect 101518 280294 101574 280350
rect 101642 280294 101698 280350
rect 101766 280294 101822 280350
rect 101394 280170 101450 280226
rect 101518 280170 101574 280226
rect 101642 280170 101698 280226
rect 101766 280170 101822 280226
rect 101394 280046 101450 280102
rect 101518 280046 101574 280102
rect 101642 280046 101698 280102
rect 101766 280046 101822 280102
rect 101394 279922 101450 279978
rect 101518 279922 101574 279978
rect 101642 279922 101698 279978
rect 101766 279922 101822 279978
rect 101394 262294 101450 262350
rect 101518 262294 101574 262350
rect 101642 262294 101698 262350
rect 101766 262294 101822 262350
rect 101394 262170 101450 262226
rect 101518 262170 101574 262226
rect 101642 262170 101698 262226
rect 101766 262170 101822 262226
rect 101394 262046 101450 262102
rect 101518 262046 101574 262102
rect 101642 262046 101698 262102
rect 101766 262046 101822 262102
rect 101394 261922 101450 261978
rect 101518 261922 101574 261978
rect 101642 261922 101698 261978
rect 101766 261922 101822 261978
rect 101394 244294 101450 244350
rect 101518 244294 101574 244350
rect 101642 244294 101698 244350
rect 101766 244294 101822 244350
rect 101394 244170 101450 244226
rect 101518 244170 101574 244226
rect 101642 244170 101698 244226
rect 101766 244170 101822 244226
rect 101394 244046 101450 244102
rect 101518 244046 101574 244102
rect 101642 244046 101698 244102
rect 101766 244046 101822 244102
rect 101394 243922 101450 243978
rect 101518 243922 101574 243978
rect 101642 243922 101698 243978
rect 101766 243922 101822 243978
rect 101394 226294 101450 226350
rect 101518 226294 101574 226350
rect 101642 226294 101698 226350
rect 101766 226294 101822 226350
rect 101394 226170 101450 226226
rect 101518 226170 101574 226226
rect 101642 226170 101698 226226
rect 101766 226170 101822 226226
rect 101394 226046 101450 226102
rect 101518 226046 101574 226102
rect 101642 226046 101698 226102
rect 101766 226046 101822 226102
rect 101394 225922 101450 225978
rect 101518 225922 101574 225978
rect 101642 225922 101698 225978
rect 101766 225922 101822 225978
rect 101394 208294 101450 208350
rect 101518 208294 101574 208350
rect 101642 208294 101698 208350
rect 101766 208294 101822 208350
rect 101394 208170 101450 208226
rect 101518 208170 101574 208226
rect 101642 208170 101698 208226
rect 101766 208170 101822 208226
rect 101394 208046 101450 208102
rect 101518 208046 101574 208102
rect 101642 208046 101698 208102
rect 101766 208046 101822 208102
rect 101394 207922 101450 207978
rect 101518 207922 101574 207978
rect 101642 207922 101698 207978
rect 101766 207922 101822 207978
rect 101394 190294 101450 190350
rect 101518 190294 101574 190350
rect 101642 190294 101698 190350
rect 101766 190294 101822 190350
rect 101394 190170 101450 190226
rect 101518 190170 101574 190226
rect 101642 190170 101698 190226
rect 101766 190170 101822 190226
rect 101394 190046 101450 190102
rect 101518 190046 101574 190102
rect 101642 190046 101698 190102
rect 101766 190046 101822 190102
rect 101394 189922 101450 189978
rect 101518 189922 101574 189978
rect 101642 189922 101698 189978
rect 101766 189922 101822 189978
rect 101394 172294 101450 172350
rect 101518 172294 101574 172350
rect 101642 172294 101698 172350
rect 101766 172294 101822 172350
rect 101394 172170 101450 172226
rect 101518 172170 101574 172226
rect 101642 172170 101698 172226
rect 101766 172170 101822 172226
rect 101394 172046 101450 172102
rect 101518 172046 101574 172102
rect 101642 172046 101698 172102
rect 101766 172046 101822 172102
rect 101394 171922 101450 171978
rect 101518 171922 101574 171978
rect 101642 171922 101698 171978
rect 101766 171922 101822 171978
rect 101394 154294 101450 154350
rect 101518 154294 101574 154350
rect 101642 154294 101698 154350
rect 101766 154294 101822 154350
rect 101394 154170 101450 154226
rect 101518 154170 101574 154226
rect 101642 154170 101698 154226
rect 101766 154170 101822 154226
rect 101394 154046 101450 154102
rect 101518 154046 101574 154102
rect 101642 154046 101698 154102
rect 101766 154046 101822 154102
rect 101394 153922 101450 153978
rect 101518 153922 101574 153978
rect 101642 153922 101698 153978
rect 101766 153922 101822 153978
rect 101394 136294 101450 136350
rect 101518 136294 101574 136350
rect 101642 136294 101698 136350
rect 101766 136294 101822 136350
rect 101394 136170 101450 136226
rect 101518 136170 101574 136226
rect 101642 136170 101698 136226
rect 101766 136170 101822 136226
rect 101394 136046 101450 136102
rect 101518 136046 101574 136102
rect 101642 136046 101698 136102
rect 101766 136046 101822 136102
rect 101394 135922 101450 135978
rect 101518 135922 101574 135978
rect 101642 135922 101698 135978
rect 101766 135922 101822 135978
rect 101394 118294 101450 118350
rect 101518 118294 101574 118350
rect 101642 118294 101698 118350
rect 101766 118294 101822 118350
rect 101394 118170 101450 118226
rect 101518 118170 101574 118226
rect 101642 118170 101698 118226
rect 101766 118170 101822 118226
rect 101394 118046 101450 118102
rect 101518 118046 101574 118102
rect 101642 118046 101698 118102
rect 101766 118046 101822 118102
rect 101394 117922 101450 117978
rect 101518 117922 101574 117978
rect 101642 117922 101698 117978
rect 101766 117922 101822 117978
rect 101394 100294 101450 100350
rect 101518 100294 101574 100350
rect 101642 100294 101698 100350
rect 101766 100294 101822 100350
rect 101394 100170 101450 100226
rect 101518 100170 101574 100226
rect 101642 100170 101698 100226
rect 101766 100170 101822 100226
rect 101394 100046 101450 100102
rect 101518 100046 101574 100102
rect 101642 100046 101698 100102
rect 101766 100046 101822 100102
rect 101394 99922 101450 99978
rect 101518 99922 101574 99978
rect 101642 99922 101698 99978
rect 101766 99922 101822 99978
rect 101394 82294 101450 82350
rect 101518 82294 101574 82350
rect 101642 82294 101698 82350
rect 101766 82294 101822 82350
rect 101394 82170 101450 82226
rect 101518 82170 101574 82226
rect 101642 82170 101698 82226
rect 101766 82170 101822 82226
rect 101394 82046 101450 82102
rect 101518 82046 101574 82102
rect 101642 82046 101698 82102
rect 101766 82046 101822 82102
rect 101394 81922 101450 81978
rect 101518 81922 101574 81978
rect 101642 81922 101698 81978
rect 101766 81922 101822 81978
rect 97674 76294 97730 76350
rect 97798 76294 97854 76350
rect 97922 76294 97978 76350
rect 98046 76294 98102 76350
rect 97674 76170 97730 76226
rect 97798 76170 97854 76226
rect 97922 76170 97978 76226
rect 98046 76170 98102 76226
rect 97674 76046 97730 76102
rect 97798 76046 97854 76102
rect 97922 76046 97978 76102
rect 98046 76046 98102 76102
rect 97674 75922 97730 75978
rect 97798 75922 97854 75978
rect 97922 75922 97978 75978
rect 98046 75922 98102 75978
rect 93318 64294 93374 64350
rect 93442 64294 93498 64350
rect 93318 64170 93374 64226
rect 93442 64170 93498 64226
rect 93318 64046 93374 64102
rect 93442 64046 93498 64102
rect 93318 63922 93374 63978
rect 93442 63922 93498 63978
rect 92876 60542 92932 60598
rect 92764 57302 92820 57358
rect 92428 8702 92484 8758
rect 92428 5462 92484 5518
rect 94220 52262 94276 52318
rect 93318 46294 93374 46350
rect 93442 46294 93498 46350
rect 93318 46170 93374 46226
rect 93442 46170 93498 46226
rect 93318 46046 93374 46102
rect 93442 46046 93498 46102
rect 93318 45922 93374 45978
rect 93442 45922 93498 45978
rect 93318 28294 93374 28350
rect 93442 28294 93498 28350
rect 93318 28170 93374 28226
rect 93442 28170 93498 28226
rect 93318 28046 93374 28102
rect 93442 28046 93498 28102
rect 93318 27922 93374 27978
rect 93442 27922 93498 27978
rect 93884 25442 93940 25498
rect 93772 16802 93828 16858
rect 93660 15182 93716 15238
rect 93100 10682 93156 10738
rect 93318 10294 93374 10350
rect 93442 10294 93498 10350
rect 93318 10170 93374 10226
rect 93442 10170 93498 10226
rect 93318 10046 93374 10102
rect 93442 10046 93498 10102
rect 93318 9922 93374 9978
rect 93442 9922 93498 9978
rect 93212 5282 93268 5338
rect 93100 4562 93156 4618
rect 93884 11762 93940 11818
rect 93884 5102 93940 5158
rect 94892 71342 94948 71398
rect 95676 62162 95732 62218
rect 95564 58922 95620 58978
rect 94892 54602 94948 54658
rect 95452 55682 95508 55738
rect 94892 54062 94948 54118
rect 95340 44162 95396 44218
rect 95340 41282 95396 41338
rect 94892 15182 94948 15238
rect 95340 15002 95396 15058
rect 94892 7442 94948 7498
rect 85708 962 85764 1018
rect 95340 6902 95396 6958
rect 97674 58294 97730 58350
rect 97798 58294 97854 58350
rect 97922 58294 97978 58350
rect 98046 58294 98102 58350
rect 97674 58170 97730 58226
rect 97798 58170 97854 58226
rect 97922 58170 97978 58226
rect 98046 58170 98102 58226
rect 97674 58046 97730 58102
rect 97798 58046 97854 58102
rect 97922 58046 97978 58102
rect 98046 58046 98102 58102
rect 97674 57922 97730 57978
rect 97798 57922 97854 57978
rect 97922 57922 97978 57978
rect 98046 57922 98102 57978
rect 96460 57122 96516 57178
rect 96236 50642 96292 50698
rect 96012 47042 96068 47098
rect 95900 15182 95956 15238
rect 96348 5462 96404 5518
rect 96572 54602 96628 54658
rect 96572 52982 96628 53038
rect 97356 50462 97412 50518
rect 97244 40562 97300 40618
rect 97132 15182 97188 15238
rect 99932 74222 99988 74278
rect 99372 55502 99428 55558
rect 97674 40294 97730 40350
rect 97798 40294 97854 40350
rect 97922 40294 97978 40350
rect 98046 40294 98102 40350
rect 97674 40170 97730 40226
rect 97798 40170 97854 40226
rect 97922 40170 97978 40226
rect 98046 40170 98102 40226
rect 97674 40046 97730 40102
rect 97798 40046 97854 40102
rect 97922 40046 97978 40102
rect 98046 40046 98102 40102
rect 97674 39922 97730 39978
rect 97798 39922 97854 39978
rect 97922 39922 97978 39978
rect 98046 39922 98102 39978
rect 97674 22294 97730 22350
rect 97798 22294 97854 22350
rect 97922 22294 97978 22350
rect 98046 22294 98102 22350
rect 97674 22170 97730 22226
rect 97798 22170 97854 22226
rect 97922 22170 97978 22226
rect 98046 22170 98102 22226
rect 97674 22046 97730 22102
rect 97798 22046 97854 22102
rect 97922 22046 97978 22102
rect 98046 22046 98102 22102
rect 97674 21922 97730 21978
rect 97798 21922 97854 21978
rect 97922 21922 97978 21978
rect 98046 21922 98102 21978
rect 97674 4294 97730 4350
rect 97798 4294 97854 4350
rect 97922 4294 97978 4350
rect 98046 4294 98102 4350
rect 97674 4170 97730 4226
rect 97798 4170 97854 4226
rect 97922 4170 97978 4226
rect 98046 4170 98102 4226
rect 97674 4046 97730 4102
rect 97798 4046 97854 4102
rect 97922 4046 97978 4102
rect 98046 4046 98102 4102
rect 97674 3922 97730 3978
rect 97798 3922 97854 3978
rect 97922 3922 97978 3978
rect 98046 3922 98102 3978
rect 70674 -1176 70730 -1120
rect 70798 -1176 70854 -1120
rect 70922 -1176 70978 -1120
rect 71046 -1176 71102 -1120
rect 70674 -1300 70730 -1244
rect 70798 -1300 70854 -1244
rect 70922 -1300 70978 -1244
rect 71046 -1300 71102 -1244
rect 70674 -1424 70730 -1368
rect 70798 -1424 70854 -1368
rect 70922 -1424 70978 -1368
rect 71046 -1424 71102 -1368
rect 70674 -1548 70730 -1492
rect 70798 -1548 70854 -1492
rect 70922 -1548 70978 -1492
rect 71046 -1548 71102 -1492
rect 98588 52082 98644 52138
rect 98700 48842 98756 48898
rect 98812 19322 98868 19378
rect 99036 7802 99092 7858
rect 98924 3164 98980 3178
rect 98924 3122 98980 3164
rect 99820 31922 99876 31978
rect 99596 6722 99652 6778
rect 99932 19322 99988 19378
rect 100044 42002 100100 42058
rect 100044 6002 100100 6058
rect 100604 67202 100660 67258
rect 100492 53882 100548 53938
rect 101394 64294 101450 64350
rect 101518 64294 101574 64350
rect 101642 64294 101698 64350
rect 101766 64294 101822 64350
rect 101394 64170 101450 64226
rect 101518 64170 101574 64226
rect 101642 64170 101698 64226
rect 101766 64170 101822 64226
rect 101394 64046 101450 64102
rect 101518 64046 101574 64102
rect 101642 64046 101698 64102
rect 101766 64046 101822 64102
rect 101394 63922 101450 63978
rect 101518 63922 101574 63978
rect 101642 63922 101698 63978
rect 101766 63922 101822 63978
rect 101394 46294 101450 46350
rect 101518 46294 101574 46350
rect 101642 46294 101698 46350
rect 101766 46294 101822 46350
rect 101394 46170 101450 46226
rect 101518 46170 101574 46226
rect 101642 46170 101698 46226
rect 101766 46170 101822 46226
rect 101394 46046 101450 46102
rect 101518 46046 101574 46102
rect 101642 46046 101698 46102
rect 101766 46046 101822 46102
rect 101394 45922 101450 45978
rect 101518 45922 101574 45978
rect 101642 45922 101698 45978
rect 101766 45922 101822 45978
rect 101394 28294 101450 28350
rect 101518 28294 101574 28350
rect 101642 28294 101698 28350
rect 101766 28294 101822 28350
rect 101394 28170 101450 28226
rect 101518 28170 101574 28226
rect 101642 28170 101698 28226
rect 101766 28170 101822 28226
rect 101394 28046 101450 28102
rect 101518 28046 101574 28102
rect 101642 28046 101698 28102
rect 101766 28046 101822 28102
rect 101394 27922 101450 27978
rect 101518 27922 101574 27978
rect 101642 27922 101698 27978
rect 101766 27922 101822 27978
rect 101394 10294 101450 10350
rect 101518 10294 101574 10350
rect 101642 10294 101698 10350
rect 101766 10294 101822 10350
rect 101394 10170 101450 10226
rect 101518 10170 101574 10226
rect 101642 10170 101698 10226
rect 101766 10170 101822 10226
rect 101394 10046 101450 10102
rect 101518 10046 101574 10102
rect 101642 10046 101698 10102
rect 101766 10046 101822 10102
rect 101394 9922 101450 9978
rect 101518 9922 101574 9978
rect 101642 9922 101698 9978
rect 101766 9922 101822 9978
rect 100492 1502 100548 1558
rect 99148 1322 99204 1378
rect 98476 1142 98532 1198
rect 97674 -216 97730 -160
rect 97798 -216 97854 -160
rect 97922 -216 97978 -160
rect 98046 -216 98102 -160
rect 97674 -340 97730 -284
rect 97798 -340 97854 -284
rect 97922 -340 97978 -284
rect 98046 -340 98102 -284
rect 97674 -464 97730 -408
rect 97798 -464 97854 -408
rect 97922 -464 97978 -408
rect 98046 -464 98102 -408
rect 97674 -588 97730 -532
rect 97798 -588 97854 -532
rect 97922 -588 97978 -532
rect 98046 -588 98102 -532
rect 102060 65582 102116 65638
rect 108678 58294 108734 58350
rect 108802 58294 108858 58350
rect 108678 58170 108734 58226
rect 108802 58170 108858 58226
rect 108678 58046 108734 58102
rect 108802 58046 108858 58102
rect 108678 57922 108734 57978
rect 108802 57922 108858 57978
rect 110796 56402 110852 56458
rect 110796 49562 110852 49618
rect 108678 40294 108734 40350
rect 108802 40294 108858 40350
rect 108678 40170 108734 40226
rect 108802 40170 108858 40226
rect 108678 40046 108734 40102
rect 108802 40046 108858 40102
rect 108678 39922 108734 39978
rect 108802 39922 108858 39978
rect 103292 35342 103348 35398
rect 102396 20942 102452 20998
rect 109228 31202 109284 31258
rect 104076 30662 104132 30718
rect 104076 25982 104132 26038
rect 107548 25262 107604 25318
rect 104188 11942 104244 11998
rect 103404 11762 103460 11818
rect 103404 6902 103460 6958
rect 103292 4562 103348 4618
rect 108332 25262 108388 25318
rect 108678 22294 108734 22350
rect 108802 22294 108858 22350
rect 108678 22170 108734 22226
rect 108802 22170 108858 22226
rect 108678 22046 108734 22102
rect 108802 22046 108858 22102
rect 108678 21922 108734 21978
rect 108802 21922 108858 21978
rect 108332 20942 108388 20998
rect 108332 7442 108388 7498
rect 108332 6902 108388 6958
rect 111020 11942 111076 11998
rect 111020 11042 111076 11098
rect 115948 34622 116004 34678
rect 115836 33902 115892 33958
rect 115836 32642 115892 32698
rect 128394 580294 128450 580350
rect 128518 580294 128574 580350
rect 128642 580294 128698 580350
rect 128766 580294 128822 580350
rect 128394 580170 128450 580226
rect 128518 580170 128574 580226
rect 128642 580170 128698 580226
rect 128766 580170 128822 580226
rect 128394 580046 128450 580102
rect 128518 580046 128574 580102
rect 128642 580046 128698 580102
rect 128766 580046 128822 580102
rect 128394 579922 128450 579978
rect 128518 579922 128574 579978
rect 128642 579922 128698 579978
rect 128766 579922 128822 579978
rect 128394 562294 128450 562350
rect 128518 562294 128574 562350
rect 128642 562294 128698 562350
rect 128766 562294 128822 562350
rect 128394 562170 128450 562226
rect 128518 562170 128574 562226
rect 128642 562170 128698 562226
rect 128766 562170 128822 562226
rect 128394 562046 128450 562102
rect 128518 562046 128574 562102
rect 128642 562046 128698 562102
rect 128766 562046 128822 562102
rect 128394 561922 128450 561978
rect 128518 561922 128574 561978
rect 128642 561922 128698 561978
rect 128766 561922 128822 561978
rect 128394 544294 128450 544350
rect 128518 544294 128574 544350
rect 128642 544294 128698 544350
rect 128766 544294 128822 544350
rect 128394 544170 128450 544226
rect 128518 544170 128574 544226
rect 128642 544170 128698 544226
rect 128766 544170 128822 544226
rect 128394 544046 128450 544102
rect 128518 544046 128574 544102
rect 128642 544046 128698 544102
rect 128766 544046 128822 544102
rect 128394 543922 128450 543978
rect 128518 543922 128574 543978
rect 128642 543922 128698 543978
rect 128766 543922 128822 543978
rect 128394 526294 128450 526350
rect 128518 526294 128574 526350
rect 128642 526294 128698 526350
rect 128766 526294 128822 526350
rect 128394 526170 128450 526226
rect 128518 526170 128574 526226
rect 128642 526170 128698 526226
rect 128766 526170 128822 526226
rect 128394 526046 128450 526102
rect 128518 526046 128574 526102
rect 128642 526046 128698 526102
rect 128766 526046 128822 526102
rect 128394 525922 128450 525978
rect 128518 525922 128574 525978
rect 128642 525922 128698 525978
rect 128766 525922 128822 525978
rect 128394 508294 128450 508350
rect 128518 508294 128574 508350
rect 128642 508294 128698 508350
rect 128766 508294 128822 508350
rect 128394 508170 128450 508226
rect 128518 508170 128574 508226
rect 128642 508170 128698 508226
rect 128766 508170 128822 508226
rect 128394 508046 128450 508102
rect 128518 508046 128574 508102
rect 128642 508046 128698 508102
rect 128766 508046 128822 508102
rect 128394 507922 128450 507978
rect 128518 507922 128574 507978
rect 128642 507922 128698 507978
rect 128766 507922 128822 507978
rect 128394 490294 128450 490350
rect 128518 490294 128574 490350
rect 128642 490294 128698 490350
rect 128766 490294 128822 490350
rect 128394 490170 128450 490226
rect 128518 490170 128574 490226
rect 128642 490170 128698 490226
rect 128766 490170 128822 490226
rect 128394 490046 128450 490102
rect 128518 490046 128574 490102
rect 128642 490046 128698 490102
rect 128766 490046 128822 490102
rect 128394 489922 128450 489978
rect 128518 489922 128574 489978
rect 128642 489922 128698 489978
rect 128766 489922 128822 489978
rect 128394 472294 128450 472350
rect 128518 472294 128574 472350
rect 128642 472294 128698 472350
rect 128766 472294 128822 472350
rect 128394 472170 128450 472226
rect 128518 472170 128574 472226
rect 128642 472170 128698 472226
rect 128766 472170 128822 472226
rect 128394 472046 128450 472102
rect 128518 472046 128574 472102
rect 128642 472046 128698 472102
rect 128766 472046 128822 472102
rect 128394 471922 128450 471978
rect 128518 471922 128574 471978
rect 128642 471922 128698 471978
rect 128766 471922 128822 471978
rect 128394 454294 128450 454350
rect 128518 454294 128574 454350
rect 128642 454294 128698 454350
rect 128766 454294 128822 454350
rect 128394 454170 128450 454226
rect 128518 454170 128574 454226
rect 128642 454170 128698 454226
rect 128766 454170 128822 454226
rect 128394 454046 128450 454102
rect 128518 454046 128574 454102
rect 128642 454046 128698 454102
rect 128766 454046 128822 454102
rect 128394 453922 128450 453978
rect 128518 453922 128574 453978
rect 128642 453922 128698 453978
rect 128766 453922 128822 453978
rect 128394 436294 128450 436350
rect 128518 436294 128574 436350
rect 128642 436294 128698 436350
rect 128766 436294 128822 436350
rect 128394 436170 128450 436226
rect 128518 436170 128574 436226
rect 128642 436170 128698 436226
rect 128766 436170 128822 436226
rect 128394 436046 128450 436102
rect 128518 436046 128574 436102
rect 128642 436046 128698 436102
rect 128766 436046 128822 436102
rect 128394 435922 128450 435978
rect 128518 435922 128574 435978
rect 128642 435922 128698 435978
rect 128766 435922 128822 435978
rect 128394 418294 128450 418350
rect 128518 418294 128574 418350
rect 128642 418294 128698 418350
rect 128766 418294 128822 418350
rect 128394 418170 128450 418226
rect 128518 418170 128574 418226
rect 128642 418170 128698 418226
rect 128766 418170 128822 418226
rect 128394 418046 128450 418102
rect 128518 418046 128574 418102
rect 128642 418046 128698 418102
rect 128766 418046 128822 418102
rect 128394 417922 128450 417978
rect 128518 417922 128574 417978
rect 128642 417922 128698 417978
rect 128766 417922 128822 417978
rect 128394 400294 128450 400350
rect 128518 400294 128574 400350
rect 128642 400294 128698 400350
rect 128766 400294 128822 400350
rect 128394 400170 128450 400226
rect 128518 400170 128574 400226
rect 128642 400170 128698 400226
rect 128766 400170 128822 400226
rect 128394 400046 128450 400102
rect 128518 400046 128574 400102
rect 128642 400046 128698 400102
rect 128766 400046 128822 400102
rect 128394 399922 128450 399978
rect 128518 399922 128574 399978
rect 128642 399922 128698 399978
rect 128766 399922 128822 399978
rect 128394 382294 128450 382350
rect 128518 382294 128574 382350
rect 128642 382294 128698 382350
rect 128766 382294 128822 382350
rect 128394 382170 128450 382226
rect 128518 382170 128574 382226
rect 128642 382170 128698 382226
rect 128766 382170 128822 382226
rect 128394 382046 128450 382102
rect 128518 382046 128574 382102
rect 128642 382046 128698 382102
rect 128766 382046 128822 382102
rect 128394 381922 128450 381978
rect 128518 381922 128574 381978
rect 128642 381922 128698 381978
rect 128766 381922 128822 381978
rect 128394 364294 128450 364350
rect 128518 364294 128574 364350
rect 128642 364294 128698 364350
rect 128766 364294 128822 364350
rect 128394 364170 128450 364226
rect 128518 364170 128574 364226
rect 128642 364170 128698 364226
rect 128766 364170 128822 364226
rect 128394 364046 128450 364102
rect 128518 364046 128574 364102
rect 128642 364046 128698 364102
rect 128766 364046 128822 364102
rect 128394 363922 128450 363978
rect 128518 363922 128574 363978
rect 128642 363922 128698 363978
rect 128766 363922 128822 363978
rect 128394 346294 128450 346350
rect 128518 346294 128574 346350
rect 128642 346294 128698 346350
rect 128766 346294 128822 346350
rect 128394 346170 128450 346226
rect 128518 346170 128574 346226
rect 128642 346170 128698 346226
rect 128766 346170 128822 346226
rect 128394 346046 128450 346102
rect 128518 346046 128574 346102
rect 128642 346046 128698 346102
rect 128766 346046 128822 346102
rect 128394 345922 128450 345978
rect 128518 345922 128574 345978
rect 128642 345922 128698 345978
rect 128766 345922 128822 345978
rect 128394 328294 128450 328350
rect 128518 328294 128574 328350
rect 128642 328294 128698 328350
rect 128766 328294 128822 328350
rect 128394 328170 128450 328226
rect 128518 328170 128574 328226
rect 128642 328170 128698 328226
rect 128766 328170 128822 328226
rect 128394 328046 128450 328102
rect 128518 328046 128574 328102
rect 128642 328046 128698 328102
rect 128766 328046 128822 328102
rect 128394 327922 128450 327978
rect 128518 327922 128574 327978
rect 128642 327922 128698 327978
rect 128766 327922 128822 327978
rect 120988 78362 121044 78418
rect 120092 54602 120148 54658
rect 120092 42722 120148 42778
rect 120988 5282 121044 5338
rect 123788 74222 123844 74278
rect 106540 3302 106596 3358
rect 128394 310294 128450 310350
rect 128518 310294 128574 310350
rect 128642 310294 128698 310350
rect 128766 310294 128822 310350
rect 128394 310170 128450 310226
rect 128518 310170 128574 310226
rect 128642 310170 128698 310226
rect 128766 310170 128822 310226
rect 128394 310046 128450 310102
rect 128518 310046 128574 310102
rect 128642 310046 128698 310102
rect 128766 310046 128822 310102
rect 128394 309922 128450 309978
rect 128518 309922 128574 309978
rect 128642 309922 128698 309978
rect 128766 309922 128822 309978
rect 128394 292294 128450 292350
rect 128518 292294 128574 292350
rect 128642 292294 128698 292350
rect 128766 292294 128822 292350
rect 128394 292170 128450 292226
rect 128518 292170 128574 292226
rect 128642 292170 128698 292226
rect 128766 292170 128822 292226
rect 128394 292046 128450 292102
rect 128518 292046 128574 292102
rect 128642 292046 128698 292102
rect 128766 292046 128822 292102
rect 128394 291922 128450 291978
rect 128518 291922 128574 291978
rect 128642 291922 128698 291978
rect 128766 291922 128822 291978
rect 128394 274294 128450 274350
rect 128518 274294 128574 274350
rect 128642 274294 128698 274350
rect 128766 274294 128822 274350
rect 128394 274170 128450 274226
rect 128518 274170 128574 274226
rect 128642 274170 128698 274226
rect 128766 274170 128822 274226
rect 128394 274046 128450 274102
rect 128518 274046 128574 274102
rect 128642 274046 128698 274102
rect 128766 274046 128822 274102
rect 128394 273922 128450 273978
rect 128518 273922 128574 273978
rect 128642 273922 128698 273978
rect 128766 273922 128822 273978
rect 128394 256294 128450 256350
rect 128518 256294 128574 256350
rect 128642 256294 128698 256350
rect 128766 256294 128822 256350
rect 128394 256170 128450 256226
rect 128518 256170 128574 256226
rect 128642 256170 128698 256226
rect 128766 256170 128822 256226
rect 128394 256046 128450 256102
rect 128518 256046 128574 256102
rect 128642 256046 128698 256102
rect 128766 256046 128822 256102
rect 128394 255922 128450 255978
rect 128518 255922 128574 255978
rect 128642 255922 128698 255978
rect 128766 255922 128822 255978
rect 128394 238294 128450 238350
rect 128518 238294 128574 238350
rect 128642 238294 128698 238350
rect 128766 238294 128822 238350
rect 128394 238170 128450 238226
rect 128518 238170 128574 238226
rect 128642 238170 128698 238226
rect 128766 238170 128822 238226
rect 128394 238046 128450 238102
rect 128518 238046 128574 238102
rect 128642 238046 128698 238102
rect 128766 238046 128822 238102
rect 128394 237922 128450 237978
rect 128518 237922 128574 237978
rect 128642 237922 128698 237978
rect 128766 237922 128822 237978
rect 128394 220294 128450 220350
rect 128518 220294 128574 220350
rect 128642 220294 128698 220350
rect 128766 220294 128822 220350
rect 128394 220170 128450 220226
rect 128518 220170 128574 220226
rect 128642 220170 128698 220226
rect 128766 220170 128822 220226
rect 128394 220046 128450 220102
rect 128518 220046 128574 220102
rect 128642 220046 128698 220102
rect 128766 220046 128822 220102
rect 128394 219922 128450 219978
rect 128518 219922 128574 219978
rect 128642 219922 128698 219978
rect 128766 219922 128822 219978
rect 126028 45602 126084 45658
rect 128394 202294 128450 202350
rect 128518 202294 128574 202350
rect 128642 202294 128698 202350
rect 128766 202294 128822 202350
rect 128394 202170 128450 202226
rect 128518 202170 128574 202226
rect 128642 202170 128698 202226
rect 128766 202170 128822 202226
rect 128394 202046 128450 202102
rect 128518 202046 128574 202102
rect 128642 202046 128698 202102
rect 128766 202046 128822 202102
rect 128394 201922 128450 201978
rect 128518 201922 128574 201978
rect 128642 201922 128698 201978
rect 128766 201922 128822 201978
rect 128394 184294 128450 184350
rect 128518 184294 128574 184350
rect 128642 184294 128698 184350
rect 128766 184294 128822 184350
rect 128394 184170 128450 184226
rect 128518 184170 128574 184226
rect 128642 184170 128698 184226
rect 128766 184170 128822 184226
rect 128394 184046 128450 184102
rect 128518 184046 128574 184102
rect 128642 184046 128698 184102
rect 128766 184046 128822 184102
rect 128394 183922 128450 183978
rect 128518 183922 128574 183978
rect 128642 183922 128698 183978
rect 128766 183922 128822 183978
rect 128394 166294 128450 166350
rect 128518 166294 128574 166350
rect 128642 166294 128698 166350
rect 128766 166294 128822 166350
rect 128394 166170 128450 166226
rect 128518 166170 128574 166226
rect 128642 166170 128698 166226
rect 128766 166170 128822 166226
rect 128394 166046 128450 166102
rect 128518 166046 128574 166102
rect 128642 166046 128698 166102
rect 128766 166046 128822 166102
rect 128394 165922 128450 165978
rect 128518 165922 128574 165978
rect 128642 165922 128698 165978
rect 128766 165922 128822 165978
rect 128394 148294 128450 148350
rect 128518 148294 128574 148350
rect 128642 148294 128698 148350
rect 128766 148294 128822 148350
rect 128394 148170 128450 148226
rect 128518 148170 128574 148226
rect 128642 148170 128698 148226
rect 128766 148170 128822 148226
rect 128394 148046 128450 148102
rect 128518 148046 128574 148102
rect 128642 148046 128698 148102
rect 128766 148046 128822 148102
rect 128394 147922 128450 147978
rect 128518 147922 128574 147978
rect 128642 147922 128698 147978
rect 128766 147922 128822 147978
rect 128394 130294 128450 130350
rect 128518 130294 128574 130350
rect 128642 130294 128698 130350
rect 128766 130294 128822 130350
rect 128394 130170 128450 130226
rect 128518 130170 128574 130226
rect 128642 130170 128698 130226
rect 128766 130170 128822 130226
rect 128394 130046 128450 130102
rect 128518 130046 128574 130102
rect 128642 130046 128698 130102
rect 128766 130046 128822 130102
rect 128394 129922 128450 129978
rect 128518 129922 128574 129978
rect 128642 129922 128698 129978
rect 128766 129922 128822 129978
rect 132114 598116 132170 598172
rect 132238 598116 132294 598172
rect 132362 598116 132418 598172
rect 132486 598116 132542 598172
rect 132114 597992 132170 598048
rect 132238 597992 132294 598048
rect 132362 597992 132418 598048
rect 132486 597992 132542 598048
rect 132114 597868 132170 597924
rect 132238 597868 132294 597924
rect 132362 597868 132418 597924
rect 132486 597868 132542 597924
rect 132114 597744 132170 597800
rect 132238 597744 132294 597800
rect 132362 597744 132418 597800
rect 132486 597744 132542 597800
rect 132114 586294 132170 586350
rect 132238 586294 132294 586350
rect 132362 586294 132418 586350
rect 132486 586294 132542 586350
rect 132114 586170 132170 586226
rect 132238 586170 132294 586226
rect 132362 586170 132418 586226
rect 132486 586170 132542 586226
rect 132114 586046 132170 586102
rect 132238 586046 132294 586102
rect 132362 586046 132418 586102
rect 132486 586046 132542 586102
rect 132114 585922 132170 585978
rect 132238 585922 132294 585978
rect 132362 585922 132418 585978
rect 132486 585922 132542 585978
rect 132114 568294 132170 568350
rect 132238 568294 132294 568350
rect 132362 568294 132418 568350
rect 132486 568294 132542 568350
rect 132114 568170 132170 568226
rect 132238 568170 132294 568226
rect 132362 568170 132418 568226
rect 132486 568170 132542 568226
rect 132114 568046 132170 568102
rect 132238 568046 132294 568102
rect 132362 568046 132418 568102
rect 132486 568046 132542 568102
rect 132114 567922 132170 567978
rect 132238 567922 132294 567978
rect 132362 567922 132418 567978
rect 132486 567922 132542 567978
rect 132114 550294 132170 550350
rect 132238 550294 132294 550350
rect 132362 550294 132418 550350
rect 132486 550294 132542 550350
rect 132114 550170 132170 550226
rect 132238 550170 132294 550226
rect 132362 550170 132418 550226
rect 132486 550170 132542 550226
rect 132114 550046 132170 550102
rect 132238 550046 132294 550102
rect 132362 550046 132418 550102
rect 132486 550046 132542 550102
rect 132114 549922 132170 549978
rect 132238 549922 132294 549978
rect 132362 549922 132418 549978
rect 132486 549922 132542 549978
rect 132114 532294 132170 532350
rect 132238 532294 132294 532350
rect 132362 532294 132418 532350
rect 132486 532294 132542 532350
rect 132114 532170 132170 532226
rect 132238 532170 132294 532226
rect 132362 532170 132418 532226
rect 132486 532170 132542 532226
rect 132114 532046 132170 532102
rect 132238 532046 132294 532102
rect 132362 532046 132418 532102
rect 132486 532046 132542 532102
rect 132114 531922 132170 531978
rect 132238 531922 132294 531978
rect 132362 531922 132418 531978
rect 132486 531922 132542 531978
rect 132114 514294 132170 514350
rect 132238 514294 132294 514350
rect 132362 514294 132418 514350
rect 132486 514294 132542 514350
rect 132114 514170 132170 514226
rect 132238 514170 132294 514226
rect 132362 514170 132418 514226
rect 132486 514170 132542 514226
rect 132114 514046 132170 514102
rect 132238 514046 132294 514102
rect 132362 514046 132418 514102
rect 132486 514046 132542 514102
rect 132114 513922 132170 513978
rect 132238 513922 132294 513978
rect 132362 513922 132418 513978
rect 132486 513922 132542 513978
rect 132114 496294 132170 496350
rect 132238 496294 132294 496350
rect 132362 496294 132418 496350
rect 132486 496294 132542 496350
rect 132114 496170 132170 496226
rect 132238 496170 132294 496226
rect 132362 496170 132418 496226
rect 132486 496170 132542 496226
rect 132114 496046 132170 496102
rect 132238 496046 132294 496102
rect 132362 496046 132418 496102
rect 132486 496046 132542 496102
rect 132114 495922 132170 495978
rect 132238 495922 132294 495978
rect 132362 495922 132418 495978
rect 132486 495922 132542 495978
rect 132114 478294 132170 478350
rect 132238 478294 132294 478350
rect 132362 478294 132418 478350
rect 132486 478294 132542 478350
rect 132114 478170 132170 478226
rect 132238 478170 132294 478226
rect 132362 478170 132418 478226
rect 132486 478170 132542 478226
rect 132114 478046 132170 478102
rect 132238 478046 132294 478102
rect 132362 478046 132418 478102
rect 132486 478046 132542 478102
rect 132114 477922 132170 477978
rect 132238 477922 132294 477978
rect 132362 477922 132418 477978
rect 132486 477922 132542 477978
rect 132114 460294 132170 460350
rect 132238 460294 132294 460350
rect 132362 460294 132418 460350
rect 132486 460294 132542 460350
rect 132114 460170 132170 460226
rect 132238 460170 132294 460226
rect 132362 460170 132418 460226
rect 132486 460170 132542 460226
rect 132114 460046 132170 460102
rect 132238 460046 132294 460102
rect 132362 460046 132418 460102
rect 132486 460046 132542 460102
rect 132114 459922 132170 459978
rect 132238 459922 132294 459978
rect 132362 459922 132418 459978
rect 132486 459922 132542 459978
rect 132114 442294 132170 442350
rect 132238 442294 132294 442350
rect 132362 442294 132418 442350
rect 132486 442294 132542 442350
rect 132114 442170 132170 442226
rect 132238 442170 132294 442226
rect 132362 442170 132418 442226
rect 132486 442170 132542 442226
rect 132114 442046 132170 442102
rect 132238 442046 132294 442102
rect 132362 442046 132418 442102
rect 132486 442046 132542 442102
rect 132114 441922 132170 441978
rect 132238 441922 132294 441978
rect 132362 441922 132418 441978
rect 132486 441922 132542 441978
rect 132114 424294 132170 424350
rect 132238 424294 132294 424350
rect 132362 424294 132418 424350
rect 132486 424294 132542 424350
rect 132114 424170 132170 424226
rect 132238 424170 132294 424226
rect 132362 424170 132418 424226
rect 132486 424170 132542 424226
rect 132114 424046 132170 424102
rect 132238 424046 132294 424102
rect 132362 424046 132418 424102
rect 132486 424046 132542 424102
rect 132114 423922 132170 423978
rect 132238 423922 132294 423978
rect 132362 423922 132418 423978
rect 132486 423922 132542 423978
rect 132114 406294 132170 406350
rect 132238 406294 132294 406350
rect 132362 406294 132418 406350
rect 132486 406294 132542 406350
rect 132114 406170 132170 406226
rect 132238 406170 132294 406226
rect 132362 406170 132418 406226
rect 132486 406170 132542 406226
rect 132114 406046 132170 406102
rect 132238 406046 132294 406102
rect 132362 406046 132418 406102
rect 132486 406046 132542 406102
rect 132114 405922 132170 405978
rect 132238 405922 132294 405978
rect 132362 405922 132418 405978
rect 132486 405922 132542 405978
rect 132114 388294 132170 388350
rect 132238 388294 132294 388350
rect 132362 388294 132418 388350
rect 132486 388294 132542 388350
rect 132114 388170 132170 388226
rect 132238 388170 132294 388226
rect 132362 388170 132418 388226
rect 132486 388170 132542 388226
rect 132114 388046 132170 388102
rect 132238 388046 132294 388102
rect 132362 388046 132418 388102
rect 132486 388046 132542 388102
rect 132114 387922 132170 387978
rect 132238 387922 132294 387978
rect 132362 387922 132418 387978
rect 132486 387922 132542 387978
rect 132114 370294 132170 370350
rect 132238 370294 132294 370350
rect 132362 370294 132418 370350
rect 132486 370294 132542 370350
rect 132114 370170 132170 370226
rect 132238 370170 132294 370226
rect 132362 370170 132418 370226
rect 132486 370170 132542 370226
rect 132114 370046 132170 370102
rect 132238 370046 132294 370102
rect 132362 370046 132418 370102
rect 132486 370046 132542 370102
rect 132114 369922 132170 369978
rect 132238 369922 132294 369978
rect 132362 369922 132418 369978
rect 132486 369922 132542 369978
rect 132114 352294 132170 352350
rect 132238 352294 132294 352350
rect 132362 352294 132418 352350
rect 132486 352294 132542 352350
rect 132114 352170 132170 352226
rect 132238 352170 132294 352226
rect 132362 352170 132418 352226
rect 132486 352170 132542 352226
rect 132114 352046 132170 352102
rect 132238 352046 132294 352102
rect 132362 352046 132418 352102
rect 132486 352046 132542 352102
rect 132114 351922 132170 351978
rect 132238 351922 132294 351978
rect 132362 351922 132418 351978
rect 132486 351922 132542 351978
rect 132114 334294 132170 334350
rect 132238 334294 132294 334350
rect 132362 334294 132418 334350
rect 132486 334294 132542 334350
rect 132114 334170 132170 334226
rect 132238 334170 132294 334226
rect 132362 334170 132418 334226
rect 132486 334170 132542 334226
rect 132114 334046 132170 334102
rect 132238 334046 132294 334102
rect 132362 334046 132418 334102
rect 132486 334046 132542 334102
rect 132114 333922 132170 333978
rect 132238 333922 132294 333978
rect 132362 333922 132418 333978
rect 132486 333922 132542 333978
rect 132114 316294 132170 316350
rect 132238 316294 132294 316350
rect 132362 316294 132418 316350
rect 132486 316294 132542 316350
rect 132114 316170 132170 316226
rect 132238 316170 132294 316226
rect 132362 316170 132418 316226
rect 132486 316170 132542 316226
rect 132114 316046 132170 316102
rect 132238 316046 132294 316102
rect 132362 316046 132418 316102
rect 132486 316046 132542 316102
rect 132114 315922 132170 315978
rect 132238 315922 132294 315978
rect 132362 315922 132418 315978
rect 132486 315922 132542 315978
rect 132114 298294 132170 298350
rect 132238 298294 132294 298350
rect 132362 298294 132418 298350
rect 132486 298294 132542 298350
rect 132114 298170 132170 298226
rect 132238 298170 132294 298226
rect 132362 298170 132418 298226
rect 132486 298170 132542 298226
rect 132114 298046 132170 298102
rect 132238 298046 132294 298102
rect 132362 298046 132418 298102
rect 132486 298046 132542 298102
rect 132114 297922 132170 297978
rect 132238 297922 132294 297978
rect 132362 297922 132418 297978
rect 132486 297922 132542 297978
rect 159114 597156 159170 597212
rect 159238 597156 159294 597212
rect 159362 597156 159418 597212
rect 159486 597156 159542 597212
rect 159114 597032 159170 597088
rect 159238 597032 159294 597088
rect 159362 597032 159418 597088
rect 159486 597032 159542 597088
rect 159114 596908 159170 596964
rect 159238 596908 159294 596964
rect 159362 596908 159418 596964
rect 159486 596908 159542 596964
rect 159114 596784 159170 596840
rect 159238 596784 159294 596840
rect 159362 596784 159418 596840
rect 159486 596784 159542 596840
rect 159114 580294 159170 580350
rect 159238 580294 159294 580350
rect 159362 580294 159418 580350
rect 159486 580294 159542 580350
rect 159114 580170 159170 580226
rect 159238 580170 159294 580226
rect 159362 580170 159418 580226
rect 159486 580170 159542 580226
rect 159114 580046 159170 580102
rect 159238 580046 159294 580102
rect 159362 580046 159418 580102
rect 159486 580046 159542 580102
rect 159114 579922 159170 579978
rect 159238 579922 159294 579978
rect 159362 579922 159418 579978
rect 159486 579922 159542 579978
rect 159114 562294 159170 562350
rect 159238 562294 159294 562350
rect 159362 562294 159418 562350
rect 159486 562294 159542 562350
rect 159114 562170 159170 562226
rect 159238 562170 159294 562226
rect 159362 562170 159418 562226
rect 159486 562170 159542 562226
rect 159114 562046 159170 562102
rect 159238 562046 159294 562102
rect 159362 562046 159418 562102
rect 159486 562046 159542 562102
rect 159114 561922 159170 561978
rect 159238 561922 159294 561978
rect 159362 561922 159418 561978
rect 159486 561922 159542 561978
rect 159114 544294 159170 544350
rect 159238 544294 159294 544350
rect 159362 544294 159418 544350
rect 159486 544294 159542 544350
rect 159114 544170 159170 544226
rect 159238 544170 159294 544226
rect 159362 544170 159418 544226
rect 159486 544170 159542 544226
rect 159114 544046 159170 544102
rect 159238 544046 159294 544102
rect 159362 544046 159418 544102
rect 159486 544046 159542 544102
rect 159114 543922 159170 543978
rect 159238 543922 159294 543978
rect 159362 543922 159418 543978
rect 159486 543922 159542 543978
rect 159114 526294 159170 526350
rect 159238 526294 159294 526350
rect 159362 526294 159418 526350
rect 159486 526294 159542 526350
rect 159114 526170 159170 526226
rect 159238 526170 159294 526226
rect 159362 526170 159418 526226
rect 159486 526170 159542 526226
rect 159114 526046 159170 526102
rect 159238 526046 159294 526102
rect 159362 526046 159418 526102
rect 159486 526046 159542 526102
rect 159114 525922 159170 525978
rect 159238 525922 159294 525978
rect 159362 525922 159418 525978
rect 159486 525922 159542 525978
rect 159114 508294 159170 508350
rect 159238 508294 159294 508350
rect 159362 508294 159418 508350
rect 159486 508294 159542 508350
rect 159114 508170 159170 508226
rect 159238 508170 159294 508226
rect 159362 508170 159418 508226
rect 159486 508170 159542 508226
rect 159114 508046 159170 508102
rect 159238 508046 159294 508102
rect 159362 508046 159418 508102
rect 159486 508046 159542 508102
rect 159114 507922 159170 507978
rect 159238 507922 159294 507978
rect 159362 507922 159418 507978
rect 159486 507922 159542 507978
rect 159114 490294 159170 490350
rect 159238 490294 159294 490350
rect 159362 490294 159418 490350
rect 159486 490294 159542 490350
rect 159114 490170 159170 490226
rect 159238 490170 159294 490226
rect 159362 490170 159418 490226
rect 159486 490170 159542 490226
rect 159114 490046 159170 490102
rect 159238 490046 159294 490102
rect 159362 490046 159418 490102
rect 159486 490046 159542 490102
rect 159114 489922 159170 489978
rect 159238 489922 159294 489978
rect 159362 489922 159418 489978
rect 159486 489922 159542 489978
rect 159114 472294 159170 472350
rect 159238 472294 159294 472350
rect 159362 472294 159418 472350
rect 159486 472294 159542 472350
rect 159114 472170 159170 472226
rect 159238 472170 159294 472226
rect 159362 472170 159418 472226
rect 159486 472170 159542 472226
rect 159114 472046 159170 472102
rect 159238 472046 159294 472102
rect 159362 472046 159418 472102
rect 159486 472046 159542 472102
rect 159114 471922 159170 471978
rect 159238 471922 159294 471978
rect 159362 471922 159418 471978
rect 159486 471922 159542 471978
rect 159114 454294 159170 454350
rect 159238 454294 159294 454350
rect 159362 454294 159418 454350
rect 159486 454294 159542 454350
rect 159114 454170 159170 454226
rect 159238 454170 159294 454226
rect 159362 454170 159418 454226
rect 159486 454170 159542 454226
rect 159114 454046 159170 454102
rect 159238 454046 159294 454102
rect 159362 454046 159418 454102
rect 159486 454046 159542 454102
rect 159114 453922 159170 453978
rect 159238 453922 159294 453978
rect 159362 453922 159418 453978
rect 159486 453922 159542 453978
rect 159114 436294 159170 436350
rect 159238 436294 159294 436350
rect 159362 436294 159418 436350
rect 159486 436294 159542 436350
rect 159114 436170 159170 436226
rect 159238 436170 159294 436226
rect 159362 436170 159418 436226
rect 159486 436170 159542 436226
rect 159114 436046 159170 436102
rect 159238 436046 159294 436102
rect 159362 436046 159418 436102
rect 159486 436046 159542 436102
rect 159114 435922 159170 435978
rect 159238 435922 159294 435978
rect 159362 435922 159418 435978
rect 159486 435922 159542 435978
rect 159114 418294 159170 418350
rect 159238 418294 159294 418350
rect 159362 418294 159418 418350
rect 159486 418294 159542 418350
rect 159114 418170 159170 418226
rect 159238 418170 159294 418226
rect 159362 418170 159418 418226
rect 159486 418170 159542 418226
rect 159114 418046 159170 418102
rect 159238 418046 159294 418102
rect 159362 418046 159418 418102
rect 159486 418046 159542 418102
rect 159114 417922 159170 417978
rect 159238 417922 159294 417978
rect 159362 417922 159418 417978
rect 159486 417922 159542 417978
rect 159114 400294 159170 400350
rect 159238 400294 159294 400350
rect 159362 400294 159418 400350
rect 159486 400294 159542 400350
rect 159114 400170 159170 400226
rect 159238 400170 159294 400226
rect 159362 400170 159418 400226
rect 159486 400170 159542 400226
rect 159114 400046 159170 400102
rect 159238 400046 159294 400102
rect 159362 400046 159418 400102
rect 159486 400046 159542 400102
rect 159114 399922 159170 399978
rect 159238 399922 159294 399978
rect 159362 399922 159418 399978
rect 159486 399922 159542 399978
rect 159114 382294 159170 382350
rect 159238 382294 159294 382350
rect 159362 382294 159418 382350
rect 159486 382294 159542 382350
rect 159114 382170 159170 382226
rect 159238 382170 159294 382226
rect 159362 382170 159418 382226
rect 159486 382170 159542 382226
rect 159114 382046 159170 382102
rect 159238 382046 159294 382102
rect 159362 382046 159418 382102
rect 159486 382046 159542 382102
rect 159114 381922 159170 381978
rect 159238 381922 159294 381978
rect 159362 381922 159418 381978
rect 159486 381922 159542 381978
rect 159114 364294 159170 364350
rect 159238 364294 159294 364350
rect 159362 364294 159418 364350
rect 159486 364294 159542 364350
rect 159114 364170 159170 364226
rect 159238 364170 159294 364226
rect 159362 364170 159418 364226
rect 159486 364170 159542 364226
rect 159114 364046 159170 364102
rect 159238 364046 159294 364102
rect 159362 364046 159418 364102
rect 159486 364046 159542 364102
rect 159114 363922 159170 363978
rect 159238 363922 159294 363978
rect 159362 363922 159418 363978
rect 159486 363922 159542 363978
rect 159114 346294 159170 346350
rect 159238 346294 159294 346350
rect 159362 346294 159418 346350
rect 159486 346294 159542 346350
rect 159114 346170 159170 346226
rect 159238 346170 159294 346226
rect 159362 346170 159418 346226
rect 159486 346170 159542 346226
rect 159114 346046 159170 346102
rect 159238 346046 159294 346102
rect 159362 346046 159418 346102
rect 159486 346046 159542 346102
rect 159114 345922 159170 345978
rect 159238 345922 159294 345978
rect 159362 345922 159418 345978
rect 159486 345922 159542 345978
rect 159114 328294 159170 328350
rect 159238 328294 159294 328350
rect 159362 328294 159418 328350
rect 159486 328294 159542 328350
rect 159114 328170 159170 328226
rect 159238 328170 159294 328226
rect 159362 328170 159418 328226
rect 159486 328170 159542 328226
rect 159114 328046 159170 328102
rect 159238 328046 159294 328102
rect 159362 328046 159418 328102
rect 159486 328046 159542 328102
rect 159114 327922 159170 327978
rect 159238 327922 159294 327978
rect 159362 327922 159418 327978
rect 159486 327922 159542 327978
rect 159114 310294 159170 310350
rect 159238 310294 159294 310350
rect 159362 310294 159418 310350
rect 159486 310294 159542 310350
rect 159114 310170 159170 310226
rect 159238 310170 159294 310226
rect 159362 310170 159418 310226
rect 159486 310170 159542 310226
rect 159114 310046 159170 310102
rect 159238 310046 159294 310102
rect 159362 310046 159418 310102
rect 159486 310046 159542 310102
rect 159114 309922 159170 309978
rect 159238 309922 159294 309978
rect 159362 309922 159418 309978
rect 159486 309922 159542 309978
rect 132114 280294 132170 280350
rect 132238 280294 132294 280350
rect 132362 280294 132418 280350
rect 132486 280294 132542 280350
rect 132114 280170 132170 280226
rect 132238 280170 132294 280226
rect 132362 280170 132418 280226
rect 132486 280170 132542 280226
rect 132114 280046 132170 280102
rect 132238 280046 132294 280102
rect 132362 280046 132418 280102
rect 132486 280046 132542 280102
rect 132114 279922 132170 279978
rect 132238 279922 132294 279978
rect 132362 279922 132418 279978
rect 132486 279922 132542 279978
rect 132114 262294 132170 262350
rect 132238 262294 132294 262350
rect 132362 262294 132418 262350
rect 132486 262294 132542 262350
rect 132114 262170 132170 262226
rect 132238 262170 132294 262226
rect 132362 262170 132418 262226
rect 132486 262170 132542 262226
rect 132114 262046 132170 262102
rect 132238 262046 132294 262102
rect 132362 262046 132418 262102
rect 132486 262046 132542 262102
rect 132114 261922 132170 261978
rect 132238 261922 132294 261978
rect 132362 261922 132418 261978
rect 132486 261922 132542 261978
rect 132114 244294 132170 244350
rect 132238 244294 132294 244350
rect 132362 244294 132418 244350
rect 132486 244294 132542 244350
rect 132114 244170 132170 244226
rect 132238 244170 132294 244226
rect 132362 244170 132418 244226
rect 132486 244170 132542 244226
rect 132114 244046 132170 244102
rect 132238 244046 132294 244102
rect 132362 244046 132418 244102
rect 132486 244046 132542 244102
rect 132114 243922 132170 243978
rect 132238 243922 132294 243978
rect 132362 243922 132418 243978
rect 132486 243922 132542 243978
rect 132114 226294 132170 226350
rect 132238 226294 132294 226350
rect 132362 226294 132418 226350
rect 132486 226294 132542 226350
rect 132114 226170 132170 226226
rect 132238 226170 132294 226226
rect 132362 226170 132418 226226
rect 132486 226170 132542 226226
rect 132114 226046 132170 226102
rect 132238 226046 132294 226102
rect 132362 226046 132418 226102
rect 132486 226046 132542 226102
rect 132114 225922 132170 225978
rect 132238 225922 132294 225978
rect 132362 225922 132418 225978
rect 132486 225922 132542 225978
rect 132114 208294 132170 208350
rect 132238 208294 132294 208350
rect 132362 208294 132418 208350
rect 132486 208294 132542 208350
rect 132114 208170 132170 208226
rect 132238 208170 132294 208226
rect 132362 208170 132418 208226
rect 132486 208170 132542 208226
rect 132114 208046 132170 208102
rect 132238 208046 132294 208102
rect 132362 208046 132418 208102
rect 132486 208046 132542 208102
rect 132114 207922 132170 207978
rect 132238 207922 132294 207978
rect 132362 207922 132418 207978
rect 132486 207922 132542 207978
rect 132114 190294 132170 190350
rect 132238 190294 132294 190350
rect 132362 190294 132418 190350
rect 132486 190294 132542 190350
rect 132114 190170 132170 190226
rect 132238 190170 132294 190226
rect 132362 190170 132418 190226
rect 132486 190170 132542 190226
rect 132114 190046 132170 190102
rect 132238 190046 132294 190102
rect 132362 190046 132418 190102
rect 132486 190046 132542 190102
rect 132114 189922 132170 189978
rect 132238 189922 132294 189978
rect 132362 189922 132418 189978
rect 132486 189922 132542 189978
rect 132114 172294 132170 172350
rect 132238 172294 132294 172350
rect 132362 172294 132418 172350
rect 132486 172294 132542 172350
rect 132114 172170 132170 172226
rect 132238 172170 132294 172226
rect 132362 172170 132418 172226
rect 132486 172170 132542 172226
rect 132114 172046 132170 172102
rect 132238 172046 132294 172102
rect 132362 172046 132418 172102
rect 132486 172046 132542 172102
rect 132114 171922 132170 171978
rect 132238 171922 132294 171978
rect 132362 171922 132418 171978
rect 132486 171922 132542 171978
rect 132114 154294 132170 154350
rect 132238 154294 132294 154350
rect 132362 154294 132418 154350
rect 132486 154294 132542 154350
rect 132114 154170 132170 154226
rect 132238 154170 132294 154226
rect 132362 154170 132418 154226
rect 132486 154170 132542 154226
rect 132114 154046 132170 154102
rect 132238 154046 132294 154102
rect 132362 154046 132418 154102
rect 132486 154046 132542 154102
rect 132114 153922 132170 153978
rect 132238 153922 132294 153978
rect 132362 153922 132418 153978
rect 132486 153922 132542 153978
rect 132114 136294 132170 136350
rect 132238 136294 132294 136350
rect 132362 136294 132418 136350
rect 132486 136294 132542 136350
rect 132114 136170 132170 136226
rect 132238 136170 132294 136226
rect 132362 136170 132418 136226
rect 132486 136170 132542 136226
rect 132114 136046 132170 136102
rect 132238 136046 132294 136102
rect 132362 136046 132418 136102
rect 132486 136046 132542 136102
rect 132114 135922 132170 135978
rect 132238 135922 132294 135978
rect 132362 135922 132418 135978
rect 132486 135922 132542 135978
rect 128394 112294 128450 112350
rect 128518 112294 128574 112350
rect 128642 112294 128698 112350
rect 128766 112294 128822 112350
rect 128394 112170 128450 112226
rect 128518 112170 128574 112226
rect 128642 112170 128698 112226
rect 128766 112170 128822 112226
rect 128394 112046 128450 112102
rect 128518 112046 128574 112102
rect 128642 112046 128698 112102
rect 128766 112046 128822 112102
rect 128394 111922 128450 111978
rect 128518 111922 128574 111978
rect 128642 111922 128698 111978
rect 128766 111922 128822 111978
rect 128394 94294 128450 94350
rect 128518 94294 128574 94350
rect 128642 94294 128698 94350
rect 128766 94294 128822 94350
rect 128394 94170 128450 94226
rect 128518 94170 128574 94226
rect 128642 94170 128698 94226
rect 128766 94170 128822 94226
rect 128394 94046 128450 94102
rect 128518 94046 128574 94102
rect 128642 94046 128698 94102
rect 128766 94046 128822 94102
rect 128394 93922 128450 93978
rect 128518 93922 128574 93978
rect 128642 93922 128698 93978
rect 128766 93922 128822 93978
rect 128394 76294 128450 76350
rect 128518 76294 128574 76350
rect 128642 76294 128698 76350
rect 128766 76294 128822 76350
rect 128394 76170 128450 76226
rect 128518 76170 128574 76226
rect 128642 76170 128698 76226
rect 128766 76170 128822 76226
rect 128394 76046 128450 76102
rect 128518 76046 128574 76102
rect 128642 76046 128698 76102
rect 128766 76046 128822 76102
rect 128394 75922 128450 75978
rect 128518 75922 128574 75978
rect 128642 75922 128698 75978
rect 128766 75922 128822 75978
rect 128394 58294 128450 58350
rect 128518 58294 128574 58350
rect 128642 58294 128698 58350
rect 128766 58294 128822 58350
rect 128394 58170 128450 58226
rect 128518 58170 128574 58226
rect 128642 58170 128698 58226
rect 128766 58170 128822 58226
rect 128394 58046 128450 58102
rect 128518 58046 128574 58102
rect 128642 58046 128698 58102
rect 128766 58046 128822 58102
rect 128394 57922 128450 57978
rect 128518 57922 128574 57978
rect 128642 57922 128698 57978
rect 128766 57922 128822 57978
rect 128394 40294 128450 40350
rect 128518 40294 128574 40350
rect 128642 40294 128698 40350
rect 128766 40294 128822 40350
rect 128394 40170 128450 40226
rect 128518 40170 128574 40226
rect 128642 40170 128698 40226
rect 128766 40170 128822 40226
rect 128394 40046 128450 40102
rect 128518 40046 128574 40102
rect 128642 40046 128698 40102
rect 128766 40046 128822 40102
rect 128394 39922 128450 39978
rect 128518 39922 128574 39978
rect 128642 39922 128698 39978
rect 128766 39922 128822 39978
rect 132114 118294 132170 118350
rect 132238 118294 132294 118350
rect 132362 118294 132418 118350
rect 132486 118294 132542 118350
rect 132114 118170 132170 118226
rect 132238 118170 132294 118226
rect 132362 118170 132418 118226
rect 132486 118170 132542 118226
rect 132114 118046 132170 118102
rect 132238 118046 132294 118102
rect 132362 118046 132418 118102
rect 132486 118046 132542 118102
rect 132114 117922 132170 117978
rect 132238 117922 132294 117978
rect 132362 117922 132418 117978
rect 132486 117922 132542 117978
rect 132114 100294 132170 100350
rect 132238 100294 132294 100350
rect 132362 100294 132418 100350
rect 132486 100294 132542 100350
rect 132114 100170 132170 100226
rect 132238 100170 132294 100226
rect 132362 100170 132418 100226
rect 132486 100170 132542 100226
rect 132114 100046 132170 100102
rect 132238 100046 132294 100102
rect 132362 100046 132418 100102
rect 132486 100046 132542 100102
rect 132114 99922 132170 99978
rect 132238 99922 132294 99978
rect 132362 99922 132418 99978
rect 132486 99922 132542 99978
rect 132114 82294 132170 82350
rect 132238 82294 132294 82350
rect 132362 82294 132418 82350
rect 132486 82294 132542 82350
rect 132114 82170 132170 82226
rect 132238 82170 132294 82226
rect 132362 82170 132418 82226
rect 132486 82170 132542 82226
rect 132114 82046 132170 82102
rect 132238 82046 132294 82102
rect 132362 82046 132418 82102
rect 132486 82046 132542 82102
rect 132114 81922 132170 81978
rect 132238 81922 132294 81978
rect 132362 81922 132418 81978
rect 132486 81922 132542 81978
rect 132114 64294 132170 64350
rect 132238 64294 132294 64350
rect 132362 64294 132418 64350
rect 132486 64294 132542 64350
rect 132114 64170 132170 64226
rect 132238 64170 132294 64226
rect 132362 64170 132418 64226
rect 132486 64170 132542 64226
rect 132114 64046 132170 64102
rect 132238 64046 132294 64102
rect 132362 64046 132418 64102
rect 132486 64046 132542 64102
rect 132114 63922 132170 63978
rect 132238 63922 132294 63978
rect 132362 63922 132418 63978
rect 132486 63922 132542 63978
rect 132114 46294 132170 46350
rect 132238 46294 132294 46350
rect 132362 46294 132418 46350
rect 132486 46294 132542 46350
rect 132114 46170 132170 46226
rect 132238 46170 132294 46226
rect 132362 46170 132418 46226
rect 132486 46170 132542 46226
rect 132114 46046 132170 46102
rect 132238 46046 132294 46102
rect 132362 46046 132418 46102
rect 132486 46046 132542 46102
rect 132114 45922 132170 45978
rect 132238 45922 132294 45978
rect 132362 45922 132418 45978
rect 132486 45922 132542 45978
rect 132114 28294 132170 28350
rect 132238 28294 132294 28350
rect 132362 28294 132418 28350
rect 132486 28294 132542 28350
rect 132114 28170 132170 28226
rect 132238 28170 132294 28226
rect 132362 28170 132418 28226
rect 132486 28170 132542 28226
rect 132114 28046 132170 28102
rect 132238 28046 132294 28102
rect 132362 28046 132418 28102
rect 132486 28046 132542 28102
rect 132114 27922 132170 27978
rect 132238 27922 132294 27978
rect 132362 27922 132418 27978
rect 132486 27922 132542 27978
rect 128394 22294 128450 22350
rect 128518 22294 128574 22350
rect 128642 22294 128698 22350
rect 128766 22294 128822 22350
rect 128394 22170 128450 22226
rect 128518 22170 128574 22226
rect 128642 22170 128698 22226
rect 128766 22170 128822 22226
rect 128394 22046 128450 22102
rect 128518 22046 128574 22102
rect 128642 22046 128698 22102
rect 128766 22046 128822 22102
rect 128394 21922 128450 21978
rect 128518 21922 128574 21978
rect 128642 21922 128698 21978
rect 128766 21922 128822 21978
rect 128394 4294 128450 4350
rect 128518 4294 128574 4350
rect 128642 4294 128698 4350
rect 128766 4294 128822 4350
rect 128394 4170 128450 4226
rect 128518 4170 128574 4226
rect 128642 4170 128698 4226
rect 128766 4170 128822 4226
rect 128394 4046 128450 4102
rect 128518 4046 128574 4102
rect 128642 4046 128698 4102
rect 128766 4046 128822 4102
rect 128394 3922 128450 3978
rect 128518 3922 128574 3978
rect 128642 3922 128698 3978
rect 128766 3922 128822 3978
rect 117964 2402 118020 2458
rect 101394 -1176 101450 -1120
rect 101518 -1176 101574 -1120
rect 101642 -1176 101698 -1120
rect 101766 -1176 101822 -1120
rect 101394 -1300 101450 -1244
rect 101518 -1300 101574 -1244
rect 101642 -1300 101698 -1244
rect 101766 -1300 101822 -1244
rect 101394 -1424 101450 -1368
rect 101518 -1424 101574 -1368
rect 101642 -1424 101698 -1368
rect 101766 -1424 101822 -1368
rect 101394 -1548 101450 -1492
rect 101518 -1548 101574 -1492
rect 101642 -1548 101698 -1492
rect 101766 -1548 101822 -1492
rect 131292 14282 131348 14338
rect 132114 10294 132170 10350
rect 132238 10294 132294 10350
rect 132362 10294 132418 10350
rect 132486 10294 132542 10350
rect 132114 10170 132170 10226
rect 132238 10170 132294 10226
rect 132362 10170 132418 10226
rect 132486 10170 132542 10226
rect 132114 10046 132170 10102
rect 132238 10046 132294 10102
rect 132362 10046 132418 10102
rect 132486 10046 132542 10102
rect 132114 9922 132170 9978
rect 132238 9922 132294 9978
rect 132362 9922 132418 9978
rect 132486 9922 132542 9978
rect 130172 1142 130228 1198
rect 128394 -216 128450 -160
rect 128518 -216 128574 -160
rect 128642 -216 128698 -160
rect 128766 -216 128822 -160
rect 128394 -340 128450 -284
rect 128518 -340 128574 -284
rect 128642 -340 128698 -284
rect 128766 -340 128822 -284
rect 128394 -464 128450 -408
rect 128518 -464 128574 -408
rect 128642 -464 128698 -408
rect 128766 -464 128822 -408
rect 128394 -588 128450 -532
rect 128518 -588 128574 -532
rect 128642 -588 128698 -532
rect 128766 -588 128822 -532
rect 132748 44522 132804 44578
rect 134428 51182 134484 51238
rect 159114 292294 159170 292350
rect 159238 292294 159294 292350
rect 159362 292294 159418 292350
rect 159486 292294 159542 292350
rect 159114 292170 159170 292226
rect 159238 292170 159294 292226
rect 159362 292170 159418 292226
rect 159486 292170 159542 292226
rect 159114 292046 159170 292102
rect 159238 292046 159294 292102
rect 159362 292046 159418 292102
rect 159486 292046 159542 292102
rect 159114 291922 159170 291978
rect 159238 291922 159294 291978
rect 159362 291922 159418 291978
rect 159486 291922 159542 291978
rect 159114 274294 159170 274350
rect 159238 274294 159294 274350
rect 159362 274294 159418 274350
rect 159486 274294 159542 274350
rect 159114 274170 159170 274226
rect 159238 274170 159294 274226
rect 159362 274170 159418 274226
rect 159486 274170 159542 274226
rect 159114 274046 159170 274102
rect 159238 274046 159294 274102
rect 159362 274046 159418 274102
rect 159486 274046 159542 274102
rect 159114 273922 159170 273978
rect 159238 273922 159294 273978
rect 159362 273922 159418 273978
rect 159486 273922 159542 273978
rect 159114 256294 159170 256350
rect 159238 256294 159294 256350
rect 159362 256294 159418 256350
rect 159486 256294 159542 256350
rect 159114 256170 159170 256226
rect 159238 256170 159294 256226
rect 159362 256170 159418 256226
rect 159486 256170 159542 256226
rect 159114 256046 159170 256102
rect 159238 256046 159294 256102
rect 159362 256046 159418 256102
rect 159486 256046 159542 256102
rect 159114 255922 159170 255978
rect 159238 255922 159294 255978
rect 159362 255922 159418 255978
rect 159486 255922 159542 255978
rect 159114 238294 159170 238350
rect 159238 238294 159294 238350
rect 159362 238294 159418 238350
rect 159486 238294 159542 238350
rect 159114 238170 159170 238226
rect 159238 238170 159294 238226
rect 159362 238170 159418 238226
rect 159486 238170 159542 238226
rect 159114 238046 159170 238102
rect 159238 238046 159294 238102
rect 159362 238046 159418 238102
rect 159486 238046 159542 238102
rect 159114 237922 159170 237978
rect 159238 237922 159294 237978
rect 159362 237922 159418 237978
rect 159486 237922 159542 237978
rect 159114 220294 159170 220350
rect 159238 220294 159294 220350
rect 159362 220294 159418 220350
rect 159486 220294 159542 220350
rect 159114 220170 159170 220226
rect 159238 220170 159294 220226
rect 159362 220170 159418 220226
rect 159486 220170 159542 220226
rect 159114 220046 159170 220102
rect 159238 220046 159294 220102
rect 159362 220046 159418 220102
rect 159486 220046 159542 220102
rect 159114 219922 159170 219978
rect 159238 219922 159294 219978
rect 159362 219922 159418 219978
rect 159486 219922 159542 219978
rect 159114 202294 159170 202350
rect 159238 202294 159294 202350
rect 159362 202294 159418 202350
rect 159486 202294 159542 202350
rect 159114 202170 159170 202226
rect 159238 202170 159294 202226
rect 159362 202170 159418 202226
rect 159486 202170 159542 202226
rect 159114 202046 159170 202102
rect 159238 202046 159294 202102
rect 159362 202046 159418 202102
rect 159486 202046 159542 202102
rect 159114 201922 159170 201978
rect 159238 201922 159294 201978
rect 159362 201922 159418 201978
rect 159486 201922 159542 201978
rect 159114 184294 159170 184350
rect 159238 184294 159294 184350
rect 159362 184294 159418 184350
rect 159486 184294 159542 184350
rect 159114 184170 159170 184226
rect 159238 184170 159294 184226
rect 159362 184170 159418 184226
rect 159486 184170 159542 184226
rect 159114 184046 159170 184102
rect 159238 184046 159294 184102
rect 159362 184046 159418 184102
rect 159486 184046 159542 184102
rect 159114 183922 159170 183978
rect 159238 183922 159294 183978
rect 159362 183922 159418 183978
rect 159486 183922 159542 183978
rect 159114 166294 159170 166350
rect 159238 166294 159294 166350
rect 159362 166294 159418 166350
rect 159486 166294 159542 166350
rect 159114 166170 159170 166226
rect 159238 166170 159294 166226
rect 159362 166170 159418 166226
rect 159486 166170 159542 166226
rect 159114 166046 159170 166102
rect 159238 166046 159294 166102
rect 159362 166046 159418 166102
rect 159486 166046 159542 166102
rect 159114 165922 159170 165978
rect 159238 165922 159294 165978
rect 159362 165922 159418 165978
rect 159486 165922 159542 165978
rect 159114 148294 159170 148350
rect 159238 148294 159294 148350
rect 159362 148294 159418 148350
rect 159486 148294 159542 148350
rect 159114 148170 159170 148226
rect 159238 148170 159294 148226
rect 159362 148170 159418 148226
rect 159486 148170 159542 148226
rect 159114 148046 159170 148102
rect 159238 148046 159294 148102
rect 159362 148046 159418 148102
rect 159486 148046 159542 148102
rect 159114 147922 159170 147978
rect 159238 147922 159294 147978
rect 159362 147922 159418 147978
rect 159486 147922 159542 147978
rect 159114 130294 159170 130350
rect 159238 130294 159294 130350
rect 159362 130294 159418 130350
rect 159486 130294 159542 130350
rect 159114 130170 159170 130226
rect 159238 130170 159294 130226
rect 159362 130170 159418 130226
rect 159486 130170 159542 130226
rect 159114 130046 159170 130102
rect 159238 130046 159294 130102
rect 159362 130046 159418 130102
rect 159486 130046 159542 130102
rect 159114 129922 159170 129978
rect 159238 129922 159294 129978
rect 159362 129922 159418 129978
rect 159486 129922 159542 129978
rect 159114 112294 159170 112350
rect 159238 112294 159294 112350
rect 159362 112294 159418 112350
rect 159486 112294 159542 112350
rect 159114 112170 159170 112226
rect 159238 112170 159294 112226
rect 159362 112170 159418 112226
rect 159486 112170 159542 112226
rect 159114 112046 159170 112102
rect 159238 112046 159294 112102
rect 159362 112046 159418 112102
rect 159486 112046 159542 112102
rect 159114 111922 159170 111978
rect 159238 111922 159294 111978
rect 159362 111922 159418 111978
rect 159486 111922 159542 111978
rect 159114 94294 159170 94350
rect 159238 94294 159294 94350
rect 159362 94294 159418 94350
rect 159486 94294 159542 94350
rect 159114 94170 159170 94226
rect 159238 94170 159294 94226
rect 159362 94170 159418 94226
rect 159486 94170 159542 94226
rect 159114 94046 159170 94102
rect 159238 94046 159294 94102
rect 159362 94046 159418 94102
rect 159486 94046 159542 94102
rect 159114 93922 159170 93978
rect 159238 93922 159294 93978
rect 159362 93922 159418 93978
rect 159486 93922 159542 93978
rect 159114 76294 159170 76350
rect 159238 76294 159294 76350
rect 159362 76294 159418 76350
rect 159486 76294 159542 76350
rect 159114 76170 159170 76226
rect 159238 76170 159294 76226
rect 159362 76170 159418 76226
rect 159486 76170 159542 76226
rect 159114 76046 159170 76102
rect 159238 76046 159294 76102
rect 159362 76046 159418 76102
rect 159486 76046 159542 76102
rect 159114 75922 159170 75978
rect 159238 75922 159294 75978
rect 159362 75922 159418 75978
rect 159486 75922 159542 75978
rect 159114 58294 159170 58350
rect 159238 58294 159294 58350
rect 159362 58294 159418 58350
rect 159486 58294 159542 58350
rect 159114 58170 159170 58226
rect 159238 58170 159294 58226
rect 159362 58170 159418 58226
rect 159486 58170 159542 58226
rect 159114 58046 159170 58102
rect 159238 58046 159294 58102
rect 159362 58046 159418 58102
rect 159486 58046 159542 58102
rect 159114 57922 159170 57978
rect 159238 57922 159294 57978
rect 159362 57922 159418 57978
rect 159486 57922 159542 57978
rect 147868 41102 147924 41158
rect 142828 29222 142884 29278
rect 137788 19142 137844 19198
rect 139468 12482 139524 12538
rect 144508 24362 144564 24418
rect 146188 15902 146244 15958
rect 159114 40294 159170 40350
rect 159238 40294 159294 40350
rect 159362 40294 159418 40350
rect 159486 40294 159542 40350
rect 159114 40170 159170 40226
rect 159238 40170 159294 40226
rect 159362 40170 159418 40226
rect 159486 40170 159542 40226
rect 159114 40046 159170 40102
rect 159238 40046 159294 40102
rect 159362 40046 159418 40102
rect 159486 40046 159542 40102
rect 159114 39922 159170 39978
rect 159238 39922 159294 39978
rect 159362 39922 159418 39978
rect 159486 39922 159542 39978
rect 151228 37682 151284 37738
rect 149548 17522 149604 17578
rect 154588 30842 154644 30898
rect 152908 24182 152964 24238
rect 159114 22294 159170 22350
rect 159238 22294 159294 22350
rect 159362 22294 159418 22350
rect 159486 22294 159542 22350
rect 159114 22170 159170 22226
rect 159238 22170 159294 22226
rect 159362 22170 159418 22226
rect 159486 22170 159542 22226
rect 159114 22046 159170 22102
rect 159238 22046 159294 22102
rect 159362 22046 159418 22102
rect 159486 22046 159542 22102
rect 159114 21922 159170 21978
rect 159238 21922 159294 21978
rect 159362 21922 159418 21978
rect 159486 21922 159542 21978
rect 157948 18962 158004 19018
rect 162834 598116 162890 598172
rect 162958 598116 163014 598172
rect 163082 598116 163138 598172
rect 163206 598116 163262 598172
rect 162834 597992 162890 598048
rect 162958 597992 163014 598048
rect 163082 597992 163138 598048
rect 163206 597992 163262 598048
rect 162834 597868 162890 597924
rect 162958 597868 163014 597924
rect 163082 597868 163138 597924
rect 163206 597868 163262 597924
rect 162834 597744 162890 597800
rect 162958 597744 163014 597800
rect 163082 597744 163138 597800
rect 163206 597744 163262 597800
rect 189834 597156 189890 597212
rect 189958 597156 190014 597212
rect 190082 597156 190138 597212
rect 190206 597156 190262 597212
rect 189834 597032 189890 597088
rect 189958 597032 190014 597088
rect 190082 597032 190138 597088
rect 190206 597032 190262 597088
rect 189834 596908 189890 596964
rect 189958 596908 190014 596964
rect 190082 596908 190138 596964
rect 190206 596908 190262 596964
rect 189834 596784 189890 596840
rect 189958 596784 190014 596840
rect 190082 596784 190138 596840
rect 190206 596784 190262 596840
rect 162834 586294 162890 586350
rect 162958 586294 163014 586350
rect 163082 586294 163138 586350
rect 163206 586294 163262 586350
rect 162834 586170 162890 586226
rect 162958 586170 163014 586226
rect 163082 586170 163138 586226
rect 163206 586170 163262 586226
rect 162834 586046 162890 586102
rect 162958 586046 163014 586102
rect 163082 586046 163138 586102
rect 163206 586046 163262 586102
rect 162834 585922 162890 585978
rect 162958 585922 163014 585978
rect 163082 585922 163138 585978
rect 163206 585922 163262 585978
rect 162834 568294 162890 568350
rect 162958 568294 163014 568350
rect 163082 568294 163138 568350
rect 163206 568294 163262 568350
rect 162834 568170 162890 568226
rect 162958 568170 163014 568226
rect 163082 568170 163138 568226
rect 163206 568170 163262 568226
rect 162834 568046 162890 568102
rect 162958 568046 163014 568102
rect 163082 568046 163138 568102
rect 163206 568046 163262 568102
rect 162834 567922 162890 567978
rect 162958 567922 163014 567978
rect 163082 567922 163138 567978
rect 163206 567922 163262 567978
rect 162834 550294 162890 550350
rect 162958 550294 163014 550350
rect 163082 550294 163138 550350
rect 163206 550294 163262 550350
rect 162834 550170 162890 550226
rect 162958 550170 163014 550226
rect 163082 550170 163138 550226
rect 163206 550170 163262 550226
rect 162834 550046 162890 550102
rect 162958 550046 163014 550102
rect 163082 550046 163138 550102
rect 163206 550046 163262 550102
rect 162834 549922 162890 549978
rect 162958 549922 163014 549978
rect 163082 549922 163138 549978
rect 163206 549922 163262 549978
rect 162834 532294 162890 532350
rect 162958 532294 163014 532350
rect 163082 532294 163138 532350
rect 163206 532294 163262 532350
rect 162834 532170 162890 532226
rect 162958 532170 163014 532226
rect 163082 532170 163138 532226
rect 163206 532170 163262 532226
rect 162834 532046 162890 532102
rect 162958 532046 163014 532102
rect 163082 532046 163138 532102
rect 163206 532046 163262 532102
rect 162834 531922 162890 531978
rect 162958 531922 163014 531978
rect 163082 531922 163138 531978
rect 163206 531922 163262 531978
rect 162834 514294 162890 514350
rect 162958 514294 163014 514350
rect 163082 514294 163138 514350
rect 163206 514294 163262 514350
rect 162834 514170 162890 514226
rect 162958 514170 163014 514226
rect 163082 514170 163138 514226
rect 163206 514170 163262 514226
rect 162834 514046 162890 514102
rect 162958 514046 163014 514102
rect 163082 514046 163138 514102
rect 163206 514046 163262 514102
rect 162834 513922 162890 513978
rect 162958 513922 163014 513978
rect 163082 513922 163138 513978
rect 163206 513922 163262 513978
rect 162834 496294 162890 496350
rect 162958 496294 163014 496350
rect 163082 496294 163138 496350
rect 163206 496294 163262 496350
rect 162834 496170 162890 496226
rect 162958 496170 163014 496226
rect 163082 496170 163138 496226
rect 163206 496170 163262 496226
rect 162834 496046 162890 496102
rect 162958 496046 163014 496102
rect 163082 496046 163138 496102
rect 163206 496046 163262 496102
rect 162834 495922 162890 495978
rect 162958 495922 163014 495978
rect 163082 495922 163138 495978
rect 163206 495922 163262 495978
rect 162834 478294 162890 478350
rect 162958 478294 163014 478350
rect 163082 478294 163138 478350
rect 163206 478294 163262 478350
rect 162834 478170 162890 478226
rect 162958 478170 163014 478226
rect 163082 478170 163138 478226
rect 163206 478170 163262 478226
rect 162834 478046 162890 478102
rect 162958 478046 163014 478102
rect 163082 478046 163138 478102
rect 163206 478046 163262 478102
rect 162834 477922 162890 477978
rect 162958 477922 163014 477978
rect 163082 477922 163138 477978
rect 163206 477922 163262 477978
rect 162834 460294 162890 460350
rect 162958 460294 163014 460350
rect 163082 460294 163138 460350
rect 163206 460294 163262 460350
rect 162834 460170 162890 460226
rect 162958 460170 163014 460226
rect 163082 460170 163138 460226
rect 163206 460170 163262 460226
rect 162834 460046 162890 460102
rect 162958 460046 163014 460102
rect 163082 460046 163138 460102
rect 163206 460046 163262 460102
rect 162834 459922 162890 459978
rect 162958 459922 163014 459978
rect 163082 459922 163138 459978
rect 163206 459922 163262 459978
rect 162834 442294 162890 442350
rect 162958 442294 163014 442350
rect 163082 442294 163138 442350
rect 163206 442294 163262 442350
rect 162834 442170 162890 442226
rect 162958 442170 163014 442226
rect 163082 442170 163138 442226
rect 163206 442170 163262 442226
rect 162834 442046 162890 442102
rect 162958 442046 163014 442102
rect 163082 442046 163138 442102
rect 163206 442046 163262 442102
rect 162834 441922 162890 441978
rect 162958 441922 163014 441978
rect 163082 441922 163138 441978
rect 163206 441922 163262 441978
rect 162834 424294 162890 424350
rect 162958 424294 163014 424350
rect 163082 424294 163138 424350
rect 163206 424294 163262 424350
rect 162834 424170 162890 424226
rect 162958 424170 163014 424226
rect 163082 424170 163138 424226
rect 163206 424170 163262 424226
rect 162834 424046 162890 424102
rect 162958 424046 163014 424102
rect 163082 424046 163138 424102
rect 163206 424046 163262 424102
rect 162834 423922 162890 423978
rect 162958 423922 163014 423978
rect 163082 423922 163138 423978
rect 163206 423922 163262 423978
rect 162834 406294 162890 406350
rect 162958 406294 163014 406350
rect 163082 406294 163138 406350
rect 163206 406294 163262 406350
rect 162834 406170 162890 406226
rect 162958 406170 163014 406226
rect 163082 406170 163138 406226
rect 163206 406170 163262 406226
rect 162834 406046 162890 406102
rect 162958 406046 163014 406102
rect 163082 406046 163138 406102
rect 163206 406046 163262 406102
rect 162834 405922 162890 405978
rect 162958 405922 163014 405978
rect 163082 405922 163138 405978
rect 163206 405922 163262 405978
rect 162834 388294 162890 388350
rect 162958 388294 163014 388350
rect 163082 388294 163138 388350
rect 163206 388294 163262 388350
rect 162834 388170 162890 388226
rect 162958 388170 163014 388226
rect 163082 388170 163138 388226
rect 163206 388170 163262 388226
rect 162834 388046 162890 388102
rect 162958 388046 163014 388102
rect 163082 388046 163138 388102
rect 163206 388046 163262 388102
rect 162834 387922 162890 387978
rect 162958 387922 163014 387978
rect 163082 387922 163138 387978
rect 163206 387922 163262 387978
rect 162834 370294 162890 370350
rect 162958 370294 163014 370350
rect 163082 370294 163138 370350
rect 163206 370294 163262 370350
rect 162834 370170 162890 370226
rect 162958 370170 163014 370226
rect 163082 370170 163138 370226
rect 163206 370170 163262 370226
rect 162834 370046 162890 370102
rect 162958 370046 163014 370102
rect 163082 370046 163138 370102
rect 163206 370046 163262 370102
rect 162834 369922 162890 369978
rect 162958 369922 163014 369978
rect 163082 369922 163138 369978
rect 163206 369922 163262 369978
rect 162834 352294 162890 352350
rect 162958 352294 163014 352350
rect 163082 352294 163138 352350
rect 163206 352294 163262 352350
rect 162834 352170 162890 352226
rect 162958 352170 163014 352226
rect 163082 352170 163138 352226
rect 163206 352170 163262 352226
rect 162834 352046 162890 352102
rect 162958 352046 163014 352102
rect 163082 352046 163138 352102
rect 163206 352046 163262 352102
rect 162834 351922 162890 351978
rect 162958 351922 163014 351978
rect 163082 351922 163138 351978
rect 163206 351922 163262 351978
rect 162834 334294 162890 334350
rect 162958 334294 163014 334350
rect 163082 334294 163138 334350
rect 163206 334294 163262 334350
rect 162834 334170 162890 334226
rect 162958 334170 163014 334226
rect 163082 334170 163138 334226
rect 163206 334170 163262 334226
rect 162834 334046 162890 334102
rect 162958 334046 163014 334102
rect 163082 334046 163138 334102
rect 163206 334046 163262 334102
rect 162834 333922 162890 333978
rect 162958 333922 163014 333978
rect 163082 333922 163138 333978
rect 163206 333922 163262 333978
rect 162834 316294 162890 316350
rect 162958 316294 163014 316350
rect 163082 316294 163138 316350
rect 163206 316294 163262 316350
rect 162834 316170 162890 316226
rect 162958 316170 163014 316226
rect 163082 316170 163138 316226
rect 163206 316170 163262 316226
rect 162834 316046 162890 316102
rect 162958 316046 163014 316102
rect 163082 316046 163138 316102
rect 163206 316046 163262 316102
rect 162834 315922 162890 315978
rect 162958 315922 163014 315978
rect 163082 315922 163138 315978
rect 163206 315922 163262 315978
rect 162834 298294 162890 298350
rect 162958 298294 163014 298350
rect 163082 298294 163138 298350
rect 163206 298294 163262 298350
rect 162834 298170 162890 298226
rect 162958 298170 163014 298226
rect 163082 298170 163138 298226
rect 163206 298170 163262 298226
rect 162834 298046 162890 298102
rect 162958 298046 163014 298102
rect 163082 298046 163138 298102
rect 163206 298046 163262 298102
rect 162834 297922 162890 297978
rect 162958 297922 163014 297978
rect 163082 297922 163138 297978
rect 163206 297922 163262 297978
rect 162834 280294 162890 280350
rect 162958 280294 163014 280350
rect 163082 280294 163138 280350
rect 163206 280294 163262 280350
rect 162834 280170 162890 280226
rect 162958 280170 163014 280226
rect 163082 280170 163138 280226
rect 163206 280170 163262 280226
rect 162834 280046 162890 280102
rect 162958 280046 163014 280102
rect 163082 280046 163138 280102
rect 163206 280046 163262 280102
rect 162834 279922 162890 279978
rect 162958 279922 163014 279978
rect 163082 279922 163138 279978
rect 163206 279922 163262 279978
rect 162834 262294 162890 262350
rect 162958 262294 163014 262350
rect 163082 262294 163138 262350
rect 163206 262294 163262 262350
rect 162834 262170 162890 262226
rect 162958 262170 163014 262226
rect 163082 262170 163138 262226
rect 163206 262170 163262 262226
rect 162834 262046 162890 262102
rect 162958 262046 163014 262102
rect 163082 262046 163138 262102
rect 163206 262046 163262 262102
rect 162834 261922 162890 261978
rect 162958 261922 163014 261978
rect 163082 261922 163138 261978
rect 163206 261922 163262 261978
rect 162834 244294 162890 244350
rect 162958 244294 163014 244350
rect 163082 244294 163138 244350
rect 163206 244294 163262 244350
rect 162834 244170 162890 244226
rect 162958 244170 163014 244226
rect 163082 244170 163138 244226
rect 163206 244170 163262 244226
rect 162834 244046 162890 244102
rect 162958 244046 163014 244102
rect 163082 244046 163138 244102
rect 163206 244046 163262 244102
rect 162834 243922 162890 243978
rect 162958 243922 163014 243978
rect 163082 243922 163138 243978
rect 163206 243922 163262 243978
rect 162834 226294 162890 226350
rect 162958 226294 163014 226350
rect 163082 226294 163138 226350
rect 163206 226294 163262 226350
rect 162834 226170 162890 226226
rect 162958 226170 163014 226226
rect 163082 226170 163138 226226
rect 163206 226170 163262 226226
rect 162834 226046 162890 226102
rect 162958 226046 163014 226102
rect 163082 226046 163138 226102
rect 163206 226046 163262 226102
rect 162834 225922 162890 225978
rect 162958 225922 163014 225978
rect 163082 225922 163138 225978
rect 163206 225922 163262 225978
rect 162834 208294 162890 208350
rect 162958 208294 163014 208350
rect 163082 208294 163138 208350
rect 163206 208294 163262 208350
rect 162834 208170 162890 208226
rect 162958 208170 163014 208226
rect 163082 208170 163138 208226
rect 163206 208170 163262 208226
rect 162834 208046 162890 208102
rect 162958 208046 163014 208102
rect 163082 208046 163138 208102
rect 163206 208046 163262 208102
rect 162834 207922 162890 207978
rect 162958 207922 163014 207978
rect 163082 207922 163138 207978
rect 163206 207922 163262 207978
rect 162834 190294 162890 190350
rect 162958 190294 163014 190350
rect 163082 190294 163138 190350
rect 163206 190294 163262 190350
rect 162834 190170 162890 190226
rect 162958 190170 163014 190226
rect 163082 190170 163138 190226
rect 163206 190170 163262 190226
rect 162834 190046 162890 190102
rect 162958 190046 163014 190102
rect 163082 190046 163138 190102
rect 163206 190046 163262 190102
rect 162834 189922 162890 189978
rect 162958 189922 163014 189978
rect 163082 189922 163138 189978
rect 163206 189922 163262 189978
rect 162834 172294 162890 172350
rect 162958 172294 163014 172350
rect 163082 172294 163138 172350
rect 163206 172294 163262 172350
rect 162834 172170 162890 172226
rect 162958 172170 163014 172226
rect 163082 172170 163138 172226
rect 163206 172170 163262 172226
rect 162834 172046 162890 172102
rect 162958 172046 163014 172102
rect 163082 172046 163138 172102
rect 163206 172046 163262 172102
rect 162834 171922 162890 171978
rect 162958 171922 163014 171978
rect 163082 171922 163138 171978
rect 163206 171922 163262 171978
rect 162834 154294 162890 154350
rect 162958 154294 163014 154350
rect 163082 154294 163138 154350
rect 163206 154294 163262 154350
rect 162834 154170 162890 154226
rect 162958 154170 163014 154226
rect 163082 154170 163138 154226
rect 163206 154170 163262 154226
rect 162834 154046 162890 154102
rect 162958 154046 163014 154102
rect 163082 154046 163138 154102
rect 163206 154046 163262 154102
rect 162834 153922 162890 153978
rect 162958 153922 163014 153978
rect 163082 153922 163138 153978
rect 163206 153922 163262 153978
rect 162834 136294 162890 136350
rect 162958 136294 163014 136350
rect 163082 136294 163138 136350
rect 163206 136294 163262 136350
rect 162834 136170 162890 136226
rect 162958 136170 163014 136226
rect 163082 136170 163138 136226
rect 163206 136170 163262 136226
rect 162834 136046 162890 136102
rect 162958 136046 163014 136102
rect 163082 136046 163138 136102
rect 163206 136046 163262 136102
rect 162834 135922 162890 135978
rect 162958 135922 163014 135978
rect 163082 135922 163138 135978
rect 163206 135922 163262 135978
rect 162834 118294 162890 118350
rect 162958 118294 163014 118350
rect 163082 118294 163138 118350
rect 163206 118294 163262 118350
rect 162834 118170 162890 118226
rect 162958 118170 163014 118226
rect 163082 118170 163138 118226
rect 163206 118170 163262 118226
rect 162834 118046 162890 118102
rect 162958 118046 163014 118102
rect 163082 118046 163138 118102
rect 163206 118046 163262 118102
rect 162834 117922 162890 117978
rect 162958 117922 163014 117978
rect 163082 117922 163138 117978
rect 163206 117922 163262 117978
rect 162834 100294 162890 100350
rect 162958 100294 163014 100350
rect 163082 100294 163138 100350
rect 163206 100294 163262 100350
rect 162834 100170 162890 100226
rect 162958 100170 163014 100226
rect 163082 100170 163138 100226
rect 163206 100170 163262 100226
rect 162834 100046 162890 100102
rect 162958 100046 163014 100102
rect 163082 100046 163138 100102
rect 163206 100046 163262 100102
rect 162834 99922 162890 99978
rect 162958 99922 163014 99978
rect 163082 99922 163138 99978
rect 163206 99922 163262 99978
rect 162834 82294 162890 82350
rect 162958 82294 163014 82350
rect 163082 82294 163138 82350
rect 163206 82294 163262 82350
rect 162834 82170 162890 82226
rect 162958 82170 163014 82226
rect 163082 82170 163138 82226
rect 163206 82170 163262 82226
rect 162834 82046 162890 82102
rect 162958 82046 163014 82102
rect 163082 82046 163138 82102
rect 163206 82046 163262 82102
rect 162834 81922 162890 81978
rect 162958 81922 163014 81978
rect 163082 81922 163138 81978
rect 163206 81922 163262 81978
rect 164668 74942 164724 74998
rect 186508 74762 186564 74818
rect 189834 580294 189890 580350
rect 189958 580294 190014 580350
rect 190082 580294 190138 580350
rect 190206 580294 190262 580350
rect 189834 580170 189890 580226
rect 189958 580170 190014 580226
rect 190082 580170 190138 580226
rect 190206 580170 190262 580226
rect 189834 580046 189890 580102
rect 189958 580046 190014 580102
rect 190082 580046 190138 580102
rect 190206 580046 190262 580102
rect 189834 579922 189890 579978
rect 189958 579922 190014 579978
rect 190082 579922 190138 579978
rect 190206 579922 190262 579978
rect 189834 562294 189890 562350
rect 189958 562294 190014 562350
rect 190082 562294 190138 562350
rect 190206 562294 190262 562350
rect 189834 562170 189890 562226
rect 189958 562170 190014 562226
rect 190082 562170 190138 562226
rect 190206 562170 190262 562226
rect 189834 562046 189890 562102
rect 189958 562046 190014 562102
rect 190082 562046 190138 562102
rect 190206 562046 190262 562102
rect 189834 561922 189890 561978
rect 189958 561922 190014 561978
rect 190082 561922 190138 561978
rect 190206 561922 190262 561978
rect 189834 544294 189890 544350
rect 189958 544294 190014 544350
rect 190082 544294 190138 544350
rect 190206 544294 190262 544350
rect 189834 544170 189890 544226
rect 189958 544170 190014 544226
rect 190082 544170 190138 544226
rect 190206 544170 190262 544226
rect 189834 544046 189890 544102
rect 189958 544046 190014 544102
rect 190082 544046 190138 544102
rect 190206 544046 190262 544102
rect 189834 543922 189890 543978
rect 189958 543922 190014 543978
rect 190082 543922 190138 543978
rect 190206 543922 190262 543978
rect 189834 526294 189890 526350
rect 189958 526294 190014 526350
rect 190082 526294 190138 526350
rect 190206 526294 190262 526350
rect 189834 526170 189890 526226
rect 189958 526170 190014 526226
rect 190082 526170 190138 526226
rect 190206 526170 190262 526226
rect 189834 526046 189890 526102
rect 189958 526046 190014 526102
rect 190082 526046 190138 526102
rect 190206 526046 190262 526102
rect 189834 525922 189890 525978
rect 189958 525922 190014 525978
rect 190082 525922 190138 525978
rect 190206 525922 190262 525978
rect 189834 508294 189890 508350
rect 189958 508294 190014 508350
rect 190082 508294 190138 508350
rect 190206 508294 190262 508350
rect 189834 508170 189890 508226
rect 189958 508170 190014 508226
rect 190082 508170 190138 508226
rect 190206 508170 190262 508226
rect 189834 508046 189890 508102
rect 189958 508046 190014 508102
rect 190082 508046 190138 508102
rect 190206 508046 190262 508102
rect 189834 507922 189890 507978
rect 189958 507922 190014 507978
rect 190082 507922 190138 507978
rect 190206 507922 190262 507978
rect 189834 490294 189890 490350
rect 189958 490294 190014 490350
rect 190082 490294 190138 490350
rect 190206 490294 190262 490350
rect 189834 490170 189890 490226
rect 189958 490170 190014 490226
rect 190082 490170 190138 490226
rect 190206 490170 190262 490226
rect 189834 490046 189890 490102
rect 189958 490046 190014 490102
rect 190082 490046 190138 490102
rect 190206 490046 190262 490102
rect 189834 489922 189890 489978
rect 189958 489922 190014 489978
rect 190082 489922 190138 489978
rect 190206 489922 190262 489978
rect 189834 472294 189890 472350
rect 189958 472294 190014 472350
rect 190082 472294 190138 472350
rect 190206 472294 190262 472350
rect 189834 472170 189890 472226
rect 189958 472170 190014 472226
rect 190082 472170 190138 472226
rect 190206 472170 190262 472226
rect 189834 472046 189890 472102
rect 189958 472046 190014 472102
rect 190082 472046 190138 472102
rect 190206 472046 190262 472102
rect 189834 471922 189890 471978
rect 189958 471922 190014 471978
rect 190082 471922 190138 471978
rect 190206 471922 190262 471978
rect 189834 454294 189890 454350
rect 189958 454294 190014 454350
rect 190082 454294 190138 454350
rect 190206 454294 190262 454350
rect 189834 454170 189890 454226
rect 189958 454170 190014 454226
rect 190082 454170 190138 454226
rect 190206 454170 190262 454226
rect 189834 454046 189890 454102
rect 189958 454046 190014 454102
rect 190082 454046 190138 454102
rect 190206 454046 190262 454102
rect 189834 453922 189890 453978
rect 189958 453922 190014 453978
rect 190082 453922 190138 453978
rect 190206 453922 190262 453978
rect 189834 436294 189890 436350
rect 189958 436294 190014 436350
rect 190082 436294 190138 436350
rect 190206 436294 190262 436350
rect 189834 436170 189890 436226
rect 189958 436170 190014 436226
rect 190082 436170 190138 436226
rect 190206 436170 190262 436226
rect 189834 436046 189890 436102
rect 189958 436046 190014 436102
rect 190082 436046 190138 436102
rect 190206 436046 190262 436102
rect 189834 435922 189890 435978
rect 189958 435922 190014 435978
rect 190082 435922 190138 435978
rect 190206 435922 190262 435978
rect 189834 418294 189890 418350
rect 189958 418294 190014 418350
rect 190082 418294 190138 418350
rect 190206 418294 190262 418350
rect 189834 418170 189890 418226
rect 189958 418170 190014 418226
rect 190082 418170 190138 418226
rect 190206 418170 190262 418226
rect 189834 418046 189890 418102
rect 189958 418046 190014 418102
rect 190082 418046 190138 418102
rect 190206 418046 190262 418102
rect 189834 417922 189890 417978
rect 189958 417922 190014 417978
rect 190082 417922 190138 417978
rect 190206 417922 190262 417978
rect 189834 400294 189890 400350
rect 189958 400294 190014 400350
rect 190082 400294 190138 400350
rect 190206 400294 190262 400350
rect 189834 400170 189890 400226
rect 189958 400170 190014 400226
rect 190082 400170 190138 400226
rect 190206 400170 190262 400226
rect 189834 400046 189890 400102
rect 189958 400046 190014 400102
rect 190082 400046 190138 400102
rect 190206 400046 190262 400102
rect 189834 399922 189890 399978
rect 189958 399922 190014 399978
rect 190082 399922 190138 399978
rect 190206 399922 190262 399978
rect 189834 382294 189890 382350
rect 189958 382294 190014 382350
rect 190082 382294 190138 382350
rect 190206 382294 190262 382350
rect 189834 382170 189890 382226
rect 189958 382170 190014 382226
rect 190082 382170 190138 382226
rect 190206 382170 190262 382226
rect 189834 382046 189890 382102
rect 189958 382046 190014 382102
rect 190082 382046 190138 382102
rect 190206 382046 190262 382102
rect 189834 381922 189890 381978
rect 189958 381922 190014 381978
rect 190082 381922 190138 381978
rect 190206 381922 190262 381978
rect 189834 364294 189890 364350
rect 189958 364294 190014 364350
rect 190082 364294 190138 364350
rect 190206 364294 190262 364350
rect 189834 364170 189890 364226
rect 189958 364170 190014 364226
rect 190082 364170 190138 364226
rect 190206 364170 190262 364226
rect 189834 364046 189890 364102
rect 189958 364046 190014 364102
rect 190082 364046 190138 364102
rect 190206 364046 190262 364102
rect 189834 363922 189890 363978
rect 189958 363922 190014 363978
rect 190082 363922 190138 363978
rect 190206 363922 190262 363978
rect 189834 346294 189890 346350
rect 189958 346294 190014 346350
rect 190082 346294 190138 346350
rect 190206 346294 190262 346350
rect 189834 346170 189890 346226
rect 189958 346170 190014 346226
rect 190082 346170 190138 346226
rect 190206 346170 190262 346226
rect 189834 346046 189890 346102
rect 189958 346046 190014 346102
rect 190082 346046 190138 346102
rect 190206 346046 190262 346102
rect 189834 345922 189890 345978
rect 189958 345922 190014 345978
rect 190082 345922 190138 345978
rect 190206 345922 190262 345978
rect 189834 328294 189890 328350
rect 189958 328294 190014 328350
rect 190082 328294 190138 328350
rect 190206 328294 190262 328350
rect 189834 328170 189890 328226
rect 189958 328170 190014 328226
rect 190082 328170 190138 328226
rect 190206 328170 190262 328226
rect 189834 328046 189890 328102
rect 189958 328046 190014 328102
rect 190082 328046 190138 328102
rect 190206 328046 190262 328102
rect 189834 327922 189890 327978
rect 189958 327922 190014 327978
rect 190082 327922 190138 327978
rect 190206 327922 190262 327978
rect 189834 310294 189890 310350
rect 189958 310294 190014 310350
rect 190082 310294 190138 310350
rect 190206 310294 190262 310350
rect 189834 310170 189890 310226
rect 189958 310170 190014 310226
rect 190082 310170 190138 310226
rect 190206 310170 190262 310226
rect 189834 310046 189890 310102
rect 189958 310046 190014 310102
rect 190082 310046 190138 310102
rect 190206 310046 190262 310102
rect 189834 309922 189890 309978
rect 189958 309922 190014 309978
rect 190082 309922 190138 309978
rect 190206 309922 190262 309978
rect 189834 292294 189890 292350
rect 189958 292294 190014 292350
rect 190082 292294 190138 292350
rect 190206 292294 190262 292350
rect 189834 292170 189890 292226
rect 189958 292170 190014 292226
rect 190082 292170 190138 292226
rect 190206 292170 190262 292226
rect 189834 292046 189890 292102
rect 189958 292046 190014 292102
rect 190082 292046 190138 292102
rect 190206 292046 190262 292102
rect 189834 291922 189890 291978
rect 189958 291922 190014 291978
rect 190082 291922 190138 291978
rect 190206 291922 190262 291978
rect 189834 274294 189890 274350
rect 189958 274294 190014 274350
rect 190082 274294 190138 274350
rect 190206 274294 190262 274350
rect 189834 274170 189890 274226
rect 189958 274170 190014 274226
rect 190082 274170 190138 274226
rect 190206 274170 190262 274226
rect 189834 274046 189890 274102
rect 189958 274046 190014 274102
rect 190082 274046 190138 274102
rect 190206 274046 190262 274102
rect 189834 273922 189890 273978
rect 189958 273922 190014 273978
rect 190082 273922 190138 273978
rect 190206 273922 190262 273978
rect 189834 256294 189890 256350
rect 189958 256294 190014 256350
rect 190082 256294 190138 256350
rect 190206 256294 190262 256350
rect 189834 256170 189890 256226
rect 189958 256170 190014 256226
rect 190082 256170 190138 256226
rect 190206 256170 190262 256226
rect 189834 256046 189890 256102
rect 189958 256046 190014 256102
rect 190082 256046 190138 256102
rect 190206 256046 190262 256102
rect 189834 255922 189890 255978
rect 189958 255922 190014 255978
rect 190082 255922 190138 255978
rect 190206 255922 190262 255978
rect 189834 238294 189890 238350
rect 189958 238294 190014 238350
rect 190082 238294 190138 238350
rect 190206 238294 190262 238350
rect 189834 238170 189890 238226
rect 189958 238170 190014 238226
rect 190082 238170 190138 238226
rect 190206 238170 190262 238226
rect 189834 238046 189890 238102
rect 189958 238046 190014 238102
rect 190082 238046 190138 238102
rect 190206 238046 190262 238102
rect 189834 237922 189890 237978
rect 189958 237922 190014 237978
rect 190082 237922 190138 237978
rect 190206 237922 190262 237978
rect 189834 220294 189890 220350
rect 189958 220294 190014 220350
rect 190082 220294 190138 220350
rect 190206 220294 190262 220350
rect 189834 220170 189890 220226
rect 189958 220170 190014 220226
rect 190082 220170 190138 220226
rect 190206 220170 190262 220226
rect 189834 220046 189890 220102
rect 189958 220046 190014 220102
rect 190082 220046 190138 220102
rect 190206 220046 190262 220102
rect 189834 219922 189890 219978
rect 189958 219922 190014 219978
rect 190082 219922 190138 219978
rect 190206 219922 190262 219978
rect 189834 202294 189890 202350
rect 189958 202294 190014 202350
rect 190082 202294 190138 202350
rect 190206 202294 190262 202350
rect 189834 202170 189890 202226
rect 189958 202170 190014 202226
rect 190082 202170 190138 202226
rect 190206 202170 190262 202226
rect 189834 202046 189890 202102
rect 189958 202046 190014 202102
rect 190082 202046 190138 202102
rect 190206 202046 190262 202102
rect 189834 201922 189890 201978
rect 189958 201922 190014 201978
rect 190082 201922 190138 201978
rect 190206 201922 190262 201978
rect 189834 184294 189890 184350
rect 189958 184294 190014 184350
rect 190082 184294 190138 184350
rect 190206 184294 190262 184350
rect 189834 184170 189890 184226
rect 189958 184170 190014 184226
rect 190082 184170 190138 184226
rect 190206 184170 190262 184226
rect 189834 184046 189890 184102
rect 189958 184046 190014 184102
rect 190082 184046 190138 184102
rect 190206 184046 190262 184102
rect 189834 183922 189890 183978
rect 189958 183922 190014 183978
rect 190082 183922 190138 183978
rect 190206 183922 190262 183978
rect 189834 166294 189890 166350
rect 189958 166294 190014 166350
rect 190082 166294 190138 166350
rect 190206 166294 190262 166350
rect 189834 166170 189890 166226
rect 189958 166170 190014 166226
rect 190082 166170 190138 166226
rect 190206 166170 190262 166226
rect 189834 166046 189890 166102
rect 189958 166046 190014 166102
rect 190082 166046 190138 166102
rect 190206 166046 190262 166102
rect 189834 165922 189890 165978
rect 189958 165922 190014 165978
rect 190082 165922 190138 165978
rect 190206 165922 190262 165978
rect 189834 148294 189890 148350
rect 189958 148294 190014 148350
rect 190082 148294 190138 148350
rect 190206 148294 190262 148350
rect 189834 148170 189890 148226
rect 189958 148170 190014 148226
rect 190082 148170 190138 148226
rect 190206 148170 190262 148226
rect 189834 148046 189890 148102
rect 189958 148046 190014 148102
rect 190082 148046 190138 148102
rect 190206 148046 190262 148102
rect 189834 147922 189890 147978
rect 189958 147922 190014 147978
rect 190082 147922 190138 147978
rect 190206 147922 190262 147978
rect 189834 130294 189890 130350
rect 189958 130294 190014 130350
rect 190082 130294 190138 130350
rect 190206 130294 190262 130350
rect 189834 130170 189890 130226
rect 189958 130170 190014 130226
rect 190082 130170 190138 130226
rect 190206 130170 190262 130226
rect 189834 130046 189890 130102
rect 189958 130046 190014 130102
rect 190082 130046 190138 130102
rect 190206 130046 190262 130102
rect 189834 129922 189890 129978
rect 189958 129922 190014 129978
rect 190082 129922 190138 129978
rect 190206 129922 190262 129978
rect 189834 112294 189890 112350
rect 189958 112294 190014 112350
rect 190082 112294 190138 112350
rect 190206 112294 190262 112350
rect 189834 112170 189890 112226
rect 189958 112170 190014 112226
rect 190082 112170 190138 112226
rect 190206 112170 190262 112226
rect 189834 112046 189890 112102
rect 189958 112046 190014 112102
rect 190082 112046 190138 112102
rect 190206 112046 190262 112102
rect 189834 111922 189890 111978
rect 189958 111922 190014 111978
rect 190082 111922 190138 111978
rect 190206 111922 190262 111978
rect 189834 94294 189890 94350
rect 189958 94294 190014 94350
rect 190082 94294 190138 94350
rect 190206 94294 190262 94350
rect 189834 94170 189890 94226
rect 189958 94170 190014 94226
rect 190082 94170 190138 94226
rect 190206 94170 190262 94226
rect 189834 94046 189890 94102
rect 189958 94046 190014 94102
rect 190082 94046 190138 94102
rect 190206 94046 190262 94102
rect 189834 93922 189890 93978
rect 189958 93922 190014 93978
rect 190082 93922 190138 93978
rect 190206 93922 190262 93978
rect 189834 76294 189890 76350
rect 189958 76294 190014 76350
rect 190082 76294 190138 76350
rect 190206 76294 190262 76350
rect 189834 76170 189890 76226
rect 189958 76170 190014 76226
rect 190082 76170 190138 76226
rect 190206 76170 190262 76226
rect 189834 76046 189890 76102
rect 189958 76046 190014 76102
rect 190082 76046 190138 76102
rect 190206 76046 190262 76102
rect 189834 75922 189890 75978
rect 189958 75922 190014 75978
rect 190082 75922 190138 75978
rect 190206 75922 190262 75978
rect 162834 64294 162890 64350
rect 162958 64294 163014 64350
rect 163082 64294 163138 64350
rect 163206 64294 163262 64350
rect 162834 64170 162890 64226
rect 162958 64170 163014 64226
rect 163082 64170 163138 64226
rect 163206 64170 163262 64226
rect 162834 64046 162890 64102
rect 162958 64046 163014 64102
rect 163082 64046 163138 64102
rect 163206 64046 163262 64102
rect 162834 63922 162890 63978
rect 162958 63922 163014 63978
rect 163082 63922 163138 63978
rect 163206 63922 163262 63978
rect 162834 46294 162890 46350
rect 162958 46294 163014 46350
rect 163082 46294 163138 46350
rect 163206 46294 163262 46350
rect 162834 46170 162890 46226
rect 162958 46170 163014 46226
rect 163082 46170 163138 46226
rect 163206 46170 163262 46226
rect 162834 46046 162890 46102
rect 162958 46046 163014 46102
rect 163082 46046 163138 46102
rect 163206 46046 163262 46102
rect 162834 45922 162890 45978
rect 162958 45922 163014 45978
rect 163082 45922 163138 45978
rect 163206 45922 163262 45978
rect 166348 61262 166404 61318
rect 162834 28294 162890 28350
rect 162958 28294 163014 28350
rect 163082 28294 163138 28350
rect 163206 28294 163262 28350
rect 162834 28170 162890 28226
rect 162958 28170 163014 28226
rect 163082 28170 163138 28226
rect 163206 28170 163262 28226
rect 162834 28046 162890 28102
rect 162958 28046 163014 28102
rect 163082 28046 163138 28102
rect 163206 28046 163262 28102
rect 162834 27922 162890 27978
rect 162958 27922 163014 27978
rect 163082 27922 163138 27978
rect 163206 27922 163262 27978
rect 159114 4294 159170 4350
rect 159238 4294 159294 4350
rect 159362 4294 159418 4350
rect 159486 4294 159542 4350
rect 159114 4170 159170 4226
rect 159238 4170 159294 4226
rect 159362 4170 159418 4226
rect 159486 4170 159542 4226
rect 132114 -1176 132170 -1120
rect 132238 -1176 132294 -1120
rect 132362 -1176 132418 -1120
rect 132486 -1176 132542 -1120
rect 132114 -1300 132170 -1244
rect 132238 -1300 132294 -1244
rect 132362 -1300 132418 -1244
rect 132486 -1300 132542 -1244
rect 132114 -1424 132170 -1368
rect 132238 -1424 132294 -1368
rect 132362 -1424 132418 -1368
rect 132486 -1424 132542 -1368
rect 132114 -1548 132170 -1492
rect 132238 -1548 132294 -1492
rect 132362 -1548 132418 -1492
rect 132486 -1548 132542 -1492
rect 161308 14102 161364 14158
rect 162834 10294 162890 10350
rect 162958 10294 163014 10350
rect 163082 10294 163138 10350
rect 163206 10294 163262 10350
rect 162834 10170 162890 10226
rect 162958 10170 163014 10226
rect 163082 10170 163138 10226
rect 163206 10170 163262 10226
rect 162834 10046 162890 10102
rect 162958 10046 163014 10102
rect 163082 10046 163138 10102
rect 163206 10046 163262 10102
rect 162834 9922 162890 9978
rect 162958 9922 163014 9978
rect 163082 9922 163138 9978
rect 163206 9922 163262 9978
rect 159114 4046 159170 4102
rect 159238 4046 159294 4102
rect 159362 4046 159418 4102
rect 159486 4046 159542 4102
rect 159114 3922 159170 3978
rect 159238 3922 159294 3978
rect 159362 3922 159418 3978
rect 159486 3922 159542 3978
rect 159114 -216 159170 -160
rect 159238 -216 159294 -160
rect 159362 -216 159418 -160
rect 159486 -216 159542 -160
rect 159114 -340 159170 -284
rect 159238 -340 159294 -284
rect 159362 -340 159418 -284
rect 159486 -340 159542 -284
rect 159114 -464 159170 -408
rect 159238 -464 159294 -408
rect 159362 -464 159418 -408
rect 159486 -464 159542 -408
rect 159114 -588 159170 -532
rect 159238 -588 159294 -532
rect 159362 -588 159418 -532
rect 159486 -588 159542 -532
rect 164668 29042 164724 29098
rect 163660 9062 163716 9118
rect 189834 58294 189890 58350
rect 189958 58294 190014 58350
rect 190082 58294 190138 58350
rect 190206 58294 190262 58350
rect 189834 58170 189890 58226
rect 189958 58170 190014 58226
rect 190082 58170 190138 58226
rect 190206 58170 190262 58226
rect 189834 58046 189890 58102
rect 189958 58046 190014 58102
rect 190082 58046 190138 58102
rect 190206 58046 190262 58102
rect 189834 57922 189890 57978
rect 189958 57922 190014 57978
rect 190082 57922 190138 57978
rect 190206 57922 190262 57978
rect 193554 598116 193610 598172
rect 193678 598116 193734 598172
rect 193802 598116 193858 598172
rect 193926 598116 193982 598172
rect 193554 597992 193610 598048
rect 193678 597992 193734 598048
rect 193802 597992 193858 598048
rect 193926 597992 193982 598048
rect 193554 597868 193610 597924
rect 193678 597868 193734 597924
rect 193802 597868 193858 597924
rect 193926 597868 193982 597924
rect 193554 597744 193610 597800
rect 193678 597744 193734 597800
rect 193802 597744 193858 597800
rect 193926 597744 193982 597800
rect 193554 586294 193610 586350
rect 193678 586294 193734 586350
rect 193802 586294 193858 586350
rect 193926 586294 193982 586350
rect 193554 586170 193610 586226
rect 193678 586170 193734 586226
rect 193802 586170 193858 586226
rect 193926 586170 193982 586226
rect 193554 586046 193610 586102
rect 193678 586046 193734 586102
rect 193802 586046 193858 586102
rect 193926 586046 193982 586102
rect 193554 585922 193610 585978
rect 193678 585922 193734 585978
rect 193802 585922 193858 585978
rect 193926 585922 193982 585978
rect 193554 568294 193610 568350
rect 193678 568294 193734 568350
rect 193802 568294 193858 568350
rect 193926 568294 193982 568350
rect 193554 568170 193610 568226
rect 193678 568170 193734 568226
rect 193802 568170 193858 568226
rect 193926 568170 193982 568226
rect 193554 568046 193610 568102
rect 193678 568046 193734 568102
rect 193802 568046 193858 568102
rect 193926 568046 193982 568102
rect 193554 567922 193610 567978
rect 193678 567922 193734 567978
rect 193802 567922 193858 567978
rect 193926 567922 193982 567978
rect 193554 550294 193610 550350
rect 193678 550294 193734 550350
rect 193802 550294 193858 550350
rect 193926 550294 193982 550350
rect 193554 550170 193610 550226
rect 193678 550170 193734 550226
rect 193802 550170 193858 550226
rect 193926 550170 193982 550226
rect 193554 550046 193610 550102
rect 193678 550046 193734 550102
rect 193802 550046 193858 550102
rect 193926 550046 193982 550102
rect 193554 549922 193610 549978
rect 193678 549922 193734 549978
rect 193802 549922 193858 549978
rect 193926 549922 193982 549978
rect 193554 532294 193610 532350
rect 193678 532294 193734 532350
rect 193802 532294 193858 532350
rect 193926 532294 193982 532350
rect 193554 532170 193610 532226
rect 193678 532170 193734 532226
rect 193802 532170 193858 532226
rect 193926 532170 193982 532226
rect 193554 532046 193610 532102
rect 193678 532046 193734 532102
rect 193802 532046 193858 532102
rect 193926 532046 193982 532102
rect 193554 531922 193610 531978
rect 193678 531922 193734 531978
rect 193802 531922 193858 531978
rect 193926 531922 193982 531978
rect 193554 514294 193610 514350
rect 193678 514294 193734 514350
rect 193802 514294 193858 514350
rect 193926 514294 193982 514350
rect 193554 514170 193610 514226
rect 193678 514170 193734 514226
rect 193802 514170 193858 514226
rect 193926 514170 193982 514226
rect 193554 514046 193610 514102
rect 193678 514046 193734 514102
rect 193802 514046 193858 514102
rect 193926 514046 193982 514102
rect 193554 513922 193610 513978
rect 193678 513922 193734 513978
rect 193802 513922 193858 513978
rect 193926 513922 193982 513978
rect 193554 496294 193610 496350
rect 193678 496294 193734 496350
rect 193802 496294 193858 496350
rect 193926 496294 193982 496350
rect 193554 496170 193610 496226
rect 193678 496170 193734 496226
rect 193802 496170 193858 496226
rect 193926 496170 193982 496226
rect 193554 496046 193610 496102
rect 193678 496046 193734 496102
rect 193802 496046 193858 496102
rect 193926 496046 193982 496102
rect 193554 495922 193610 495978
rect 193678 495922 193734 495978
rect 193802 495922 193858 495978
rect 193926 495922 193982 495978
rect 193554 478294 193610 478350
rect 193678 478294 193734 478350
rect 193802 478294 193858 478350
rect 193926 478294 193982 478350
rect 193554 478170 193610 478226
rect 193678 478170 193734 478226
rect 193802 478170 193858 478226
rect 193926 478170 193982 478226
rect 193554 478046 193610 478102
rect 193678 478046 193734 478102
rect 193802 478046 193858 478102
rect 193926 478046 193982 478102
rect 193554 477922 193610 477978
rect 193678 477922 193734 477978
rect 193802 477922 193858 477978
rect 193926 477922 193982 477978
rect 193554 460294 193610 460350
rect 193678 460294 193734 460350
rect 193802 460294 193858 460350
rect 193926 460294 193982 460350
rect 193554 460170 193610 460226
rect 193678 460170 193734 460226
rect 193802 460170 193858 460226
rect 193926 460170 193982 460226
rect 193554 460046 193610 460102
rect 193678 460046 193734 460102
rect 193802 460046 193858 460102
rect 193926 460046 193982 460102
rect 193554 459922 193610 459978
rect 193678 459922 193734 459978
rect 193802 459922 193858 459978
rect 193926 459922 193982 459978
rect 193554 442294 193610 442350
rect 193678 442294 193734 442350
rect 193802 442294 193858 442350
rect 193926 442294 193982 442350
rect 193554 442170 193610 442226
rect 193678 442170 193734 442226
rect 193802 442170 193858 442226
rect 193926 442170 193982 442226
rect 193554 442046 193610 442102
rect 193678 442046 193734 442102
rect 193802 442046 193858 442102
rect 193926 442046 193982 442102
rect 193554 441922 193610 441978
rect 193678 441922 193734 441978
rect 193802 441922 193858 441978
rect 193926 441922 193982 441978
rect 193554 424294 193610 424350
rect 193678 424294 193734 424350
rect 193802 424294 193858 424350
rect 193926 424294 193982 424350
rect 193554 424170 193610 424226
rect 193678 424170 193734 424226
rect 193802 424170 193858 424226
rect 193926 424170 193982 424226
rect 193554 424046 193610 424102
rect 193678 424046 193734 424102
rect 193802 424046 193858 424102
rect 193926 424046 193982 424102
rect 193554 423922 193610 423978
rect 193678 423922 193734 423978
rect 193802 423922 193858 423978
rect 193926 423922 193982 423978
rect 193554 406294 193610 406350
rect 193678 406294 193734 406350
rect 193802 406294 193858 406350
rect 193926 406294 193982 406350
rect 193554 406170 193610 406226
rect 193678 406170 193734 406226
rect 193802 406170 193858 406226
rect 193926 406170 193982 406226
rect 193554 406046 193610 406102
rect 193678 406046 193734 406102
rect 193802 406046 193858 406102
rect 193926 406046 193982 406102
rect 193554 405922 193610 405978
rect 193678 405922 193734 405978
rect 193802 405922 193858 405978
rect 193926 405922 193982 405978
rect 193554 388294 193610 388350
rect 193678 388294 193734 388350
rect 193802 388294 193858 388350
rect 193926 388294 193982 388350
rect 193554 388170 193610 388226
rect 193678 388170 193734 388226
rect 193802 388170 193858 388226
rect 193926 388170 193982 388226
rect 193554 388046 193610 388102
rect 193678 388046 193734 388102
rect 193802 388046 193858 388102
rect 193926 388046 193982 388102
rect 193554 387922 193610 387978
rect 193678 387922 193734 387978
rect 193802 387922 193858 387978
rect 193926 387922 193982 387978
rect 193554 370294 193610 370350
rect 193678 370294 193734 370350
rect 193802 370294 193858 370350
rect 193926 370294 193982 370350
rect 193554 370170 193610 370226
rect 193678 370170 193734 370226
rect 193802 370170 193858 370226
rect 193926 370170 193982 370226
rect 193554 370046 193610 370102
rect 193678 370046 193734 370102
rect 193802 370046 193858 370102
rect 193926 370046 193982 370102
rect 193554 369922 193610 369978
rect 193678 369922 193734 369978
rect 193802 369922 193858 369978
rect 193926 369922 193982 369978
rect 193554 352294 193610 352350
rect 193678 352294 193734 352350
rect 193802 352294 193858 352350
rect 193926 352294 193982 352350
rect 193554 352170 193610 352226
rect 193678 352170 193734 352226
rect 193802 352170 193858 352226
rect 193926 352170 193982 352226
rect 193554 352046 193610 352102
rect 193678 352046 193734 352102
rect 193802 352046 193858 352102
rect 193926 352046 193982 352102
rect 193554 351922 193610 351978
rect 193678 351922 193734 351978
rect 193802 351922 193858 351978
rect 193926 351922 193982 351978
rect 193554 334294 193610 334350
rect 193678 334294 193734 334350
rect 193802 334294 193858 334350
rect 193926 334294 193982 334350
rect 193554 334170 193610 334226
rect 193678 334170 193734 334226
rect 193802 334170 193858 334226
rect 193926 334170 193982 334226
rect 193554 334046 193610 334102
rect 193678 334046 193734 334102
rect 193802 334046 193858 334102
rect 193926 334046 193982 334102
rect 193554 333922 193610 333978
rect 193678 333922 193734 333978
rect 193802 333922 193858 333978
rect 193926 333922 193982 333978
rect 193554 316294 193610 316350
rect 193678 316294 193734 316350
rect 193802 316294 193858 316350
rect 193926 316294 193982 316350
rect 193554 316170 193610 316226
rect 193678 316170 193734 316226
rect 193802 316170 193858 316226
rect 193926 316170 193982 316226
rect 193554 316046 193610 316102
rect 193678 316046 193734 316102
rect 193802 316046 193858 316102
rect 193926 316046 193982 316102
rect 193554 315922 193610 315978
rect 193678 315922 193734 315978
rect 193802 315922 193858 315978
rect 193926 315922 193982 315978
rect 193554 298294 193610 298350
rect 193678 298294 193734 298350
rect 193802 298294 193858 298350
rect 193926 298294 193982 298350
rect 193554 298170 193610 298226
rect 193678 298170 193734 298226
rect 193802 298170 193858 298226
rect 193926 298170 193982 298226
rect 193554 298046 193610 298102
rect 193678 298046 193734 298102
rect 193802 298046 193858 298102
rect 193926 298046 193982 298102
rect 193554 297922 193610 297978
rect 193678 297922 193734 297978
rect 193802 297922 193858 297978
rect 193926 297922 193982 297978
rect 193554 280294 193610 280350
rect 193678 280294 193734 280350
rect 193802 280294 193858 280350
rect 193926 280294 193982 280350
rect 193554 280170 193610 280226
rect 193678 280170 193734 280226
rect 193802 280170 193858 280226
rect 193926 280170 193982 280226
rect 193554 280046 193610 280102
rect 193678 280046 193734 280102
rect 193802 280046 193858 280102
rect 193926 280046 193982 280102
rect 193554 279922 193610 279978
rect 193678 279922 193734 279978
rect 193802 279922 193858 279978
rect 193926 279922 193982 279978
rect 193554 262294 193610 262350
rect 193678 262294 193734 262350
rect 193802 262294 193858 262350
rect 193926 262294 193982 262350
rect 193554 262170 193610 262226
rect 193678 262170 193734 262226
rect 193802 262170 193858 262226
rect 193926 262170 193982 262226
rect 193554 262046 193610 262102
rect 193678 262046 193734 262102
rect 193802 262046 193858 262102
rect 193926 262046 193982 262102
rect 193554 261922 193610 261978
rect 193678 261922 193734 261978
rect 193802 261922 193858 261978
rect 193926 261922 193982 261978
rect 193554 244294 193610 244350
rect 193678 244294 193734 244350
rect 193802 244294 193858 244350
rect 193926 244294 193982 244350
rect 193554 244170 193610 244226
rect 193678 244170 193734 244226
rect 193802 244170 193858 244226
rect 193926 244170 193982 244226
rect 193554 244046 193610 244102
rect 193678 244046 193734 244102
rect 193802 244046 193858 244102
rect 193926 244046 193982 244102
rect 193554 243922 193610 243978
rect 193678 243922 193734 243978
rect 193802 243922 193858 243978
rect 193926 243922 193982 243978
rect 193554 226294 193610 226350
rect 193678 226294 193734 226350
rect 193802 226294 193858 226350
rect 193926 226294 193982 226350
rect 193554 226170 193610 226226
rect 193678 226170 193734 226226
rect 193802 226170 193858 226226
rect 193926 226170 193982 226226
rect 193554 226046 193610 226102
rect 193678 226046 193734 226102
rect 193802 226046 193858 226102
rect 193926 226046 193982 226102
rect 193554 225922 193610 225978
rect 193678 225922 193734 225978
rect 193802 225922 193858 225978
rect 193926 225922 193982 225978
rect 193554 208294 193610 208350
rect 193678 208294 193734 208350
rect 193802 208294 193858 208350
rect 193926 208294 193982 208350
rect 193554 208170 193610 208226
rect 193678 208170 193734 208226
rect 193802 208170 193858 208226
rect 193926 208170 193982 208226
rect 193554 208046 193610 208102
rect 193678 208046 193734 208102
rect 193802 208046 193858 208102
rect 193926 208046 193982 208102
rect 193554 207922 193610 207978
rect 193678 207922 193734 207978
rect 193802 207922 193858 207978
rect 193926 207922 193982 207978
rect 193554 190294 193610 190350
rect 193678 190294 193734 190350
rect 193802 190294 193858 190350
rect 193926 190294 193982 190350
rect 193554 190170 193610 190226
rect 193678 190170 193734 190226
rect 193802 190170 193858 190226
rect 193926 190170 193982 190226
rect 193554 190046 193610 190102
rect 193678 190046 193734 190102
rect 193802 190046 193858 190102
rect 193926 190046 193982 190102
rect 193554 189922 193610 189978
rect 193678 189922 193734 189978
rect 193802 189922 193858 189978
rect 193926 189922 193982 189978
rect 193554 172294 193610 172350
rect 193678 172294 193734 172350
rect 193802 172294 193858 172350
rect 193926 172294 193982 172350
rect 193554 172170 193610 172226
rect 193678 172170 193734 172226
rect 193802 172170 193858 172226
rect 193926 172170 193982 172226
rect 193554 172046 193610 172102
rect 193678 172046 193734 172102
rect 193802 172046 193858 172102
rect 193926 172046 193982 172102
rect 193554 171922 193610 171978
rect 193678 171922 193734 171978
rect 193802 171922 193858 171978
rect 193926 171922 193982 171978
rect 193554 154294 193610 154350
rect 193678 154294 193734 154350
rect 193802 154294 193858 154350
rect 193926 154294 193982 154350
rect 193554 154170 193610 154226
rect 193678 154170 193734 154226
rect 193802 154170 193858 154226
rect 193926 154170 193982 154226
rect 193554 154046 193610 154102
rect 193678 154046 193734 154102
rect 193802 154046 193858 154102
rect 193926 154046 193982 154102
rect 193554 153922 193610 153978
rect 193678 153922 193734 153978
rect 193802 153922 193858 153978
rect 193926 153922 193982 153978
rect 193554 136294 193610 136350
rect 193678 136294 193734 136350
rect 193802 136294 193858 136350
rect 193926 136294 193982 136350
rect 193554 136170 193610 136226
rect 193678 136170 193734 136226
rect 193802 136170 193858 136226
rect 193926 136170 193982 136226
rect 193554 136046 193610 136102
rect 193678 136046 193734 136102
rect 193802 136046 193858 136102
rect 193926 136046 193982 136102
rect 193554 135922 193610 135978
rect 193678 135922 193734 135978
rect 193802 135922 193858 135978
rect 193926 135922 193982 135978
rect 193554 118294 193610 118350
rect 193678 118294 193734 118350
rect 193802 118294 193858 118350
rect 193926 118294 193982 118350
rect 193554 118170 193610 118226
rect 193678 118170 193734 118226
rect 193802 118170 193858 118226
rect 193926 118170 193982 118226
rect 193554 118046 193610 118102
rect 193678 118046 193734 118102
rect 193802 118046 193858 118102
rect 193926 118046 193982 118102
rect 193554 117922 193610 117978
rect 193678 117922 193734 117978
rect 193802 117922 193858 117978
rect 193926 117922 193982 117978
rect 193554 100294 193610 100350
rect 193678 100294 193734 100350
rect 193802 100294 193858 100350
rect 193926 100294 193982 100350
rect 193554 100170 193610 100226
rect 193678 100170 193734 100226
rect 193802 100170 193858 100226
rect 193926 100170 193982 100226
rect 193554 100046 193610 100102
rect 193678 100046 193734 100102
rect 193802 100046 193858 100102
rect 193926 100046 193982 100102
rect 193554 99922 193610 99978
rect 193678 99922 193734 99978
rect 193802 99922 193858 99978
rect 193926 99922 193982 99978
rect 193554 82294 193610 82350
rect 193678 82294 193734 82350
rect 193802 82294 193858 82350
rect 193926 82294 193982 82350
rect 193554 82170 193610 82226
rect 193678 82170 193734 82226
rect 193802 82170 193858 82226
rect 193926 82170 193982 82226
rect 193554 82046 193610 82102
rect 193678 82046 193734 82102
rect 193802 82046 193858 82102
rect 193926 82046 193982 82102
rect 193554 81922 193610 81978
rect 193678 81922 193734 81978
rect 193802 81922 193858 81978
rect 193926 81922 193982 81978
rect 220554 597156 220610 597212
rect 220678 597156 220734 597212
rect 220802 597156 220858 597212
rect 220926 597156 220982 597212
rect 220554 597032 220610 597088
rect 220678 597032 220734 597088
rect 220802 597032 220858 597088
rect 220926 597032 220982 597088
rect 220554 596908 220610 596964
rect 220678 596908 220734 596964
rect 220802 596908 220858 596964
rect 220926 596908 220982 596964
rect 220554 596784 220610 596840
rect 220678 596784 220734 596840
rect 220802 596784 220858 596840
rect 220926 596784 220982 596840
rect 220554 580294 220610 580350
rect 220678 580294 220734 580350
rect 220802 580294 220858 580350
rect 220926 580294 220982 580350
rect 220554 580170 220610 580226
rect 220678 580170 220734 580226
rect 220802 580170 220858 580226
rect 220926 580170 220982 580226
rect 220554 580046 220610 580102
rect 220678 580046 220734 580102
rect 220802 580046 220858 580102
rect 220926 580046 220982 580102
rect 220554 579922 220610 579978
rect 220678 579922 220734 579978
rect 220802 579922 220858 579978
rect 220926 579922 220982 579978
rect 220554 562294 220610 562350
rect 220678 562294 220734 562350
rect 220802 562294 220858 562350
rect 220926 562294 220982 562350
rect 220554 562170 220610 562226
rect 220678 562170 220734 562226
rect 220802 562170 220858 562226
rect 220926 562170 220982 562226
rect 220554 562046 220610 562102
rect 220678 562046 220734 562102
rect 220802 562046 220858 562102
rect 220926 562046 220982 562102
rect 220554 561922 220610 561978
rect 220678 561922 220734 561978
rect 220802 561922 220858 561978
rect 220926 561922 220982 561978
rect 220554 544294 220610 544350
rect 220678 544294 220734 544350
rect 220802 544294 220858 544350
rect 220926 544294 220982 544350
rect 220554 544170 220610 544226
rect 220678 544170 220734 544226
rect 220802 544170 220858 544226
rect 220926 544170 220982 544226
rect 220554 544046 220610 544102
rect 220678 544046 220734 544102
rect 220802 544046 220858 544102
rect 220926 544046 220982 544102
rect 220554 543922 220610 543978
rect 220678 543922 220734 543978
rect 220802 543922 220858 543978
rect 220926 543922 220982 543978
rect 220554 526294 220610 526350
rect 220678 526294 220734 526350
rect 220802 526294 220858 526350
rect 220926 526294 220982 526350
rect 220554 526170 220610 526226
rect 220678 526170 220734 526226
rect 220802 526170 220858 526226
rect 220926 526170 220982 526226
rect 220554 526046 220610 526102
rect 220678 526046 220734 526102
rect 220802 526046 220858 526102
rect 220926 526046 220982 526102
rect 220554 525922 220610 525978
rect 220678 525922 220734 525978
rect 220802 525922 220858 525978
rect 220926 525922 220982 525978
rect 220554 508294 220610 508350
rect 220678 508294 220734 508350
rect 220802 508294 220858 508350
rect 220926 508294 220982 508350
rect 220554 508170 220610 508226
rect 220678 508170 220734 508226
rect 220802 508170 220858 508226
rect 220926 508170 220982 508226
rect 220554 508046 220610 508102
rect 220678 508046 220734 508102
rect 220802 508046 220858 508102
rect 220926 508046 220982 508102
rect 220554 507922 220610 507978
rect 220678 507922 220734 507978
rect 220802 507922 220858 507978
rect 220926 507922 220982 507978
rect 220554 490294 220610 490350
rect 220678 490294 220734 490350
rect 220802 490294 220858 490350
rect 220926 490294 220982 490350
rect 220554 490170 220610 490226
rect 220678 490170 220734 490226
rect 220802 490170 220858 490226
rect 220926 490170 220982 490226
rect 220554 490046 220610 490102
rect 220678 490046 220734 490102
rect 220802 490046 220858 490102
rect 220926 490046 220982 490102
rect 220554 489922 220610 489978
rect 220678 489922 220734 489978
rect 220802 489922 220858 489978
rect 220926 489922 220982 489978
rect 220554 472294 220610 472350
rect 220678 472294 220734 472350
rect 220802 472294 220858 472350
rect 220926 472294 220982 472350
rect 220554 472170 220610 472226
rect 220678 472170 220734 472226
rect 220802 472170 220858 472226
rect 220926 472170 220982 472226
rect 220554 472046 220610 472102
rect 220678 472046 220734 472102
rect 220802 472046 220858 472102
rect 220926 472046 220982 472102
rect 220554 471922 220610 471978
rect 220678 471922 220734 471978
rect 220802 471922 220858 471978
rect 220926 471922 220982 471978
rect 220554 454294 220610 454350
rect 220678 454294 220734 454350
rect 220802 454294 220858 454350
rect 220926 454294 220982 454350
rect 220554 454170 220610 454226
rect 220678 454170 220734 454226
rect 220802 454170 220858 454226
rect 220926 454170 220982 454226
rect 220554 454046 220610 454102
rect 220678 454046 220734 454102
rect 220802 454046 220858 454102
rect 220926 454046 220982 454102
rect 220554 453922 220610 453978
rect 220678 453922 220734 453978
rect 220802 453922 220858 453978
rect 220926 453922 220982 453978
rect 220554 436294 220610 436350
rect 220678 436294 220734 436350
rect 220802 436294 220858 436350
rect 220926 436294 220982 436350
rect 220554 436170 220610 436226
rect 220678 436170 220734 436226
rect 220802 436170 220858 436226
rect 220926 436170 220982 436226
rect 220554 436046 220610 436102
rect 220678 436046 220734 436102
rect 220802 436046 220858 436102
rect 220926 436046 220982 436102
rect 220554 435922 220610 435978
rect 220678 435922 220734 435978
rect 220802 435922 220858 435978
rect 220926 435922 220982 435978
rect 220554 418294 220610 418350
rect 220678 418294 220734 418350
rect 220802 418294 220858 418350
rect 220926 418294 220982 418350
rect 220554 418170 220610 418226
rect 220678 418170 220734 418226
rect 220802 418170 220858 418226
rect 220926 418170 220982 418226
rect 220554 418046 220610 418102
rect 220678 418046 220734 418102
rect 220802 418046 220858 418102
rect 220926 418046 220982 418102
rect 220554 417922 220610 417978
rect 220678 417922 220734 417978
rect 220802 417922 220858 417978
rect 220926 417922 220982 417978
rect 220554 400294 220610 400350
rect 220678 400294 220734 400350
rect 220802 400294 220858 400350
rect 220926 400294 220982 400350
rect 220554 400170 220610 400226
rect 220678 400170 220734 400226
rect 220802 400170 220858 400226
rect 220926 400170 220982 400226
rect 220554 400046 220610 400102
rect 220678 400046 220734 400102
rect 220802 400046 220858 400102
rect 220926 400046 220982 400102
rect 220554 399922 220610 399978
rect 220678 399922 220734 399978
rect 220802 399922 220858 399978
rect 220926 399922 220982 399978
rect 220554 382294 220610 382350
rect 220678 382294 220734 382350
rect 220802 382294 220858 382350
rect 220926 382294 220982 382350
rect 220554 382170 220610 382226
rect 220678 382170 220734 382226
rect 220802 382170 220858 382226
rect 220926 382170 220982 382226
rect 220554 382046 220610 382102
rect 220678 382046 220734 382102
rect 220802 382046 220858 382102
rect 220926 382046 220982 382102
rect 220554 381922 220610 381978
rect 220678 381922 220734 381978
rect 220802 381922 220858 381978
rect 220926 381922 220982 381978
rect 220554 364294 220610 364350
rect 220678 364294 220734 364350
rect 220802 364294 220858 364350
rect 220926 364294 220982 364350
rect 220554 364170 220610 364226
rect 220678 364170 220734 364226
rect 220802 364170 220858 364226
rect 220926 364170 220982 364226
rect 220554 364046 220610 364102
rect 220678 364046 220734 364102
rect 220802 364046 220858 364102
rect 220926 364046 220982 364102
rect 220554 363922 220610 363978
rect 220678 363922 220734 363978
rect 220802 363922 220858 363978
rect 220926 363922 220982 363978
rect 220554 346294 220610 346350
rect 220678 346294 220734 346350
rect 220802 346294 220858 346350
rect 220926 346294 220982 346350
rect 220554 346170 220610 346226
rect 220678 346170 220734 346226
rect 220802 346170 220858 346226
rect 220926 346170 220982 346226
rect 220554 346046 220610 346102
rect 220678 346046 220734 346102
rect 220802 346046 220858 346102
rect 220926 346046 220982 346102
rect 220554 345922 220610 345978
rect 220678 345922 220734 345978
rect 220802 345922 220858 345978
rect 220926 345922 220982 345978
rect 220554 328294 220610 328350
rect 220678 328294 220734 328350
rect 220802 328294 220858 328350
rect 220926 328294 220982 328350
rect 220554 328170 220610 328226
rect 220678 328170 220734 328226
rect 220802 328170 220858 328226
rect 220926 328170 220982 328226
rect 220554 328046 220610 328102
rect 220678 328046 220734 328102
rect 220802 328046 220858 328102
rect 220926 328046 220982 328102
rect 220554 327922 220610 327978
rect 220678 327922 220734 327978
rect 220802 327922 220858 327978
rect 220926 327922 220982 327978
rect 220554 310294 220610 310350
rect 220678 310294 220734 310350
rect 220802 310294 220858 310350
rect 220926 310294 220982 310350
rect 220554 310170 220610 310226
rect 220678 310170 220734 310226
rect 220802 310170 220858 310226
rect 220926 310170 220982 310226
rect 220554 310046 220610 310102
rect 220678 310046 220734 310102
rect 220802 310046 220858 310102
rect 220926 310046 220982 310102
rect 220554 309922 220610 309978
rect 220678 309922 220734 309978
rect 220802 309922 220858 309978
rect 220926 309922 220982 309978
rect 220554 292294 220610 292350
rect 220678 292294 220734 292350
rect 220802 292294 220858 292350
rect 220926 292294 220982 292350
rect 220554 292170 220610 292226
rect 220678 292170 220734 292226
rect 220802 292170 220858 292226
rect 220926 292170 220982 292226
rect 220554 292046 220610 292102
rect 220678 292046 220734 292102
rect 220802 292046 220858 292102
rect 220926 292046 220982 292102
rect 220554 291922 220610 291978
rect 220678 291922 220734 291978
rect 220802 291922 220858 291978
rect 220926 291922 220982 291978
rect 220554 274294 220610 274350
rect 220678 274294 220734 274350
rect 220802 274294 220858 274350
rect 220926 274294 220982 274350
rect 220554 274170 220610 274226
rect 220678 274170 220734 274226
rect 220802 274170 220858 274226
rect 220926 274170 220982 274226
rect 220554 274046 220610 274102
rect 220678 274046 220734 274102
rect 220802 274046 220858 274102
rect 220926 274046 220982 274102
rect 220554 273922 220610 273978
rect 220678 273922 220734 273978
rect 220802 273922 220858 273978
rect 220926 273922 220982 273978
rect 220554 256294 220610 256350
rect 220678 256294 220734 256350
rect 220802 256294 220858 256350
rect 220926 256294 220982 256350
rect 220554 256170 220610 256226
rect 220678 256170 220734 256226
rect 220802 256170 220858 256226
rect 220926 256170 220982 256226
rect 220554 256046 220610 256102
rect 220678 256046 220734 256102
rect 220802 256046 220858 256102
rect 220926 256046 220982 256102
rect 220554 255922 220610 255978
rect 220678 255922 220734 255978
rect 220802 255922 220858 255978
rect 220926 255922 220982 255978
rect 220554 238294 220610 238350
rect 220678 238294 220734 238350
rect 220802 238294 220858 238350
rect 220926 238294 220982 238350
rect 220554 238170 220610 238226
rect 220678 238170 220734 238226
rect 220802 238170 220858 238226
rect 220926 238170 220982 238226
rect 220554 238046 220610 238102
rect 220678 238046 220734 238102
rect 220802 238046 220858 238102
rect 220926 238046 220982 238102
rect 220554 237922 220610 237978
rect 220678 237922 220734 237978
rect 220802 237922 220858 237978
rect 220926 237922 220982 237978
rect 220554 220294 220610 220350
rect 220678 220294 220734 220350
rect 220802 220294 220858 220350
rect 220926 220294 220982 220350
rect 220554 220170 220610 220226
rect 220678 220170 220734 220226
rect 220802 220170 220858 220226
rect 220926 220170 220982 220226
rect 220554 220046 220610 220102
rect 220678 220046 220734 220102
rect 220802 220046 220858 220102
rect 220926 220046 220982 220102
rect 220554 219922 220610 219978
rect 220678 219922 220734 219978
rect 220802 219922 220858 219978
rect 220926 219922 220982 219978
rect 220554 202294 220610 202350
rect 220678 202294 220734 202350
rect 220802 202294 220858 202350
rect 220926 202294 220982 202350
rect 220554 202170 220610 202226
rect 220678 202170 220734 202226
rect 220802 202170 220858 202226
rect 220926 202170 220982 202226
rect 220554 202046 220610 202102
rect 220678 202046 220734 202102
rect 220802 202046 220858 202102
rect 220926 202046 220982 202102
rect 220554 201922 220610 201978
rect 220678 201922 220734 201978
rect 220802 201922 220858 201978
rect 220926 201922 220982 201978
rect 220554 184294 220610 184350
rect 220678 184294 220734 184350
rect 220802 184294 220858 184350
rect 220926 184294 220982 184350
rect 220554 184170 220610 184226
rect 220678 184170 220734 184226
rect 220802 184170 220858 184226
rect 220926 184170 220982 184226
rect 220554 184046 220610 184102
rect 220678 184046 220734 184102
rect 220802 184046 220858 184102
rect 220926 184046 220982 184102
rect 220554 183922 220610 183978
rect 220678 183922 220734 183978
rect 220802 183922 220858 183978
rect 220926 183922 220982 183978
rect 220554 166294 220610 166350
rect 220678 166294 220734 166350
rect 220802 166294 220858 166350
rect 220926 166294 220982 166350
rect 220554 166170 220610 166226
rect 220678 166170 220734 166226
rect 220802 166170 220858 166226
rect 220926 166170 220982 166226
rect 220554 166046 220610 166102
rect 220678 166046 220734 166102
rect 220802 166046 220858 166102
rect 220926 166046 220982 166102
rect 220554 165922 220610 165978
rect 220678 165922 220734 165978
rect 220802 165922 220858 165978
rect 220926 165922 220982 165978
rect 220554 148294 220610 148350
rect 220678 148294 220734 148350
rect 220802 148294 220858 148350
rect 220926 148294 220982 148350
rect 220554 148170 220610 148226
rect 220678 148170 220734 148226
rect 220802 148170 220858 148226
rect 220926 148170 220982 148226
rect 220554 148046 220610 148102
rect 220678 148046 220734 148102
rect 220802 148046 220858 148102
rect 220926 148046 220982 148102
rect 220554 147922 220610 147978
rect 220678 147922 220734 147978
rect 220802 147922 220858 147978
rect 220926 147922 220982 147978
rect 220554 130294 220610 130350
rect 220678 130294 220734 130350
rect 220802 130294 220858 130350
rect 220926 130294 220982 130350
rect 220554 130170 220610 130226
rect 220678 130170 220734 130226
rect 220802 130170 220858 130226
rect 220926 130170 220982 130226
rect 220554 130046 220610 130102
rect 220678 130046 220734 130102
rect 220802 130046 220858 130102
rect 220926 130046 220982 130102
rect 220554 129922 220610 129978
rect 220678 129922 220734 129978
rect 220802 129922 220858 129978
rect 220926 129922 220982 129978
rect 220554 112294 220610 112350
rect 220678 112294 220734 112350
rect 220802 112294 220858 112350
rect 220926 112294 220982 112350
rect 220554 112170 220610 112226
rect 220678 112170 220734 112226
rect 220802 112170 220858 112226
rect 220926 112170 220982 112226
rect 220554 112046 220610 112102
rect 220678 112046 220734 112102
rect 220802 112046 220858 112102
rect 220926 112046 220982 112102
rect 220554 111922 220610 111978
rect 220678 111922 220734 111978
rect 220802 111922 220858 111978
rect 220926 111922 220982 111978
rect 220554 94294 220610 94350
rect 220678 94294 220734 94350
rect 220802 94294 220858 94350
rect 220926 94294 220982 94350
rect 220554 94170 220610 94226
rect 220678 94170 220734 94226
rect 220802 94170 220858 94226
rect 220926 94170 220982 94226
rect 220554 94046 220610 94102
rect 220678 94046 220734 94102
rect 220802 94046 220858 94102
rect 220926 94046 220982 94102
rect 220554 93922 220610 93978
rect 220678 93922 220734 93978
rect 220802 93922 220858 93978
rect 220926 93922 220982 93978
rect 220554 76294 220610 76350
rect 220678 76294 220734 76350
rect 220802 76294 220858 76350
rect 220926 76294 220982 76350
rect 220554 76170 220610 76226
rect 220678 76170 220734 76226
rect 220802 76170 220858 76226
rect 220926 76170 220982 76226
rect 220554 76046 220610 76102
rect 220678 76046 220734 76102
rect 220802 76046 220858 76102
rect 220926 76046 220982 76102
rect 220554 75922 220610 75978
rect 220678 75922 220734 75978
rect 220802 75922 220858 75978
rect 220926 75922 220982 75978
rect 193554 64294 193610 64350
rect 193678 64294 193734 64350
rect 193802 64294 193858 64350
rect 193926 64294 193982 64350
rect 193554 64170 193610 64226
rect 193678 64170 193734 64226
rect 193802 64170 193858 64226
rect 193926 64170 193982 64226
rect 193554 64046 193610 64102
rect 193678 64046 193734 64102
rect 193802 64046 193858 64102
rect 193926 64046 193982 64102
rect 193554 63922 193610 63978
rect 193678 63922 193734 63978
rect 193802 63922 193858 63978
rect 193926 63922 193982 63978
rect 193554 46294 193610 46350
rect 193678 46294 193734 46350
rect 193802 46294 193858 46350
rect 193926 46294 193982 46350
rect 193554 46170 193610 46226
rect 193678 46170 193734 46226
rect 193802 46170 193858 46226
rect 193926 46170 193982 46226
rect 193554 46046 193610 46102
rect 193678 46046 193734 46102
rect 193802 46046 193858 46102
rect 193926 46046 193982 46102
rect 193554 45922 193610 45978
rect 193678 45922 193734 45978
rect 193802 45922 193858 45978
rect 193926 45922 193982 45978
rect 189834 40294 189890 40350
rect 189958 40294 190014 40350
rect 190082 40294 190138 40350
rect 190206 40294 190262 40350
rect 189834 40170 189890 40226
rect 189958 40170 190014 40226
rect 190082 40170 190138 40226
rect 190206 40170 190262 40226
rect 189834 40046 189890 40102
rect 189958 40046 190014 40102
rect 190082 40046 190138 40102
rect 190206 40046 190262 40102
rect 189834 39922 189890 39978
rect 189958 39922 190014 39978
rect 190082 39922 190138 39978
rect 190206 39922 190262 39978
rect 178108 32462 178164 32518
rect 173068 26882 173124 26938
rect 174748 20582 174804 20638
rect 169372 8882 169428 8938
rect 189834 22294 189890 22350
rect 189958 22294 190014 22350
rect 190082 22294 190138 22350
rect 190206 22294 190262 22350
rect 189834 22170 189890 22226
rect 189958 22170 190014 22226
rect 190082 22170 190138 22226
rect 190206 22170 190262 22226
rect 189834 22046 189890 22102
rect 189958 22046 190014 22102
rect 190082 22046 190138 22102
rect 190206 22046 190262 22102
rect 189834 21922 189890 21978
rect 189958 21922 190014 21978
rect 190082 21922 190138 21978
rect 190206 21922 190262 21978
rect 183148 17342 183204 17398
rect 179788 13922 179844 13978
rect 189834 4294 189890 4350
rect 189958 4294 190014 4350
rect 190082 4294 190138 4350
rect 190206 4294 190262 4350
rect 189834 4170 189890 4226
rect 189958 4170 190014 4226
rect 190082 4170 190138 4226
rect 190206 4170 190262 4226
rect 162834 -1176 162890 -1120
rect 162958 -1176 163014 -1120
rect 163082 -1176 163138 -1120
rect 163206 -1176 163262 -1120
rect 162834 -1300 162890 -1244
rect 162958 -1300 163014 -1244
rect 163082 -1300 163138 -1244
rect 163206 -1300 163262 -1244
rect 162834 -1424 162890 -1368
rect 162958 -1424 163014 -1368
rect 163082 -1424 163138 -1368
rect 163206 -1424 163262 -1368
rect 162834 -1548 162890 -1492
rect 162958 -1548 163014 -1492
rect 163082 -1548 163138 -1492
rect 163206 -1548 163262 -1492
rect 190428 45422 190484 45478
rect 193554 28294 193610 28350
rect 193678 28294 193734 28350
rect 193802 28294 193858 28350
rect 193926 28294 193982 28350
rect 193554 28170 193610 28226
rect 193678 28170 193734 28226
rect 193802 28170 193858 28226
rect 193926 28170 193982 28226
rect 193554 28046 193610 28102
rect 193678 28046 193734 28102
rect 193802 28046 193858 28102
rect 193926 28046 193982 28102
rect 193554 27922 193610 27978
rect 193678 27922 193734 27978
rect 193802 27922 193858 27978
rect 193926 27922 193982 27978
rect 191548 18782 191604 18838
rect 206668 71342 206724 71398
rect 193554 10294 193610 10350
rect 193678 10294 193734 10350
rect 193802 10294 193858 10350
rect 193926 10294 193982 10350
rect 193554 10170 193610 10226
rect 193678 10170 193734 10226
rect 193802 10170 193858 10226
rect 193926 10170 193982 10226
rect 193554 10046 193610 10102
rect 193678 10046 193734 10102
rect 193802 10046 193858 10102
rect 193926 10046 193982 10102
rect 193554 9922 193610 9978
rect 193678 9922 193734 9978
rect 193802 9922 193858 9978
rect 193926 9922 193982 9978
rect 189834 4046 189890 4102
rect 189958 4046 190014 4102
rect 190082 4046 190138 4102
rect 190206 4046 190262 4102
rect 189834 3922 189890 3978
rect 189958 3922 190014 3978
rect 190082 3922 190138 3978
rect 190206 3922 190262 3978
rect 193228 3482 193284 3538
rect 189834 -216 189890 -160
rect 189958 -216 190014 -160
rect 190082 -216 190138 -160
rect 190206 -216 190262 -160
rect 189834 -340 189890 -284
rect 189958 -340 190014 -284
rect 190082 -340 190138 -284
rect 190206 -340 190262 -284
rect 189834 -464 189890 -408
rect 189958 -464 190014 -408
rect 190082 -464 190138 -408
rect 190206 -464 190262 -408
rect 189834 -588 189890 -532
rect 189958 -588 190014 -532
rect 190082 -588 190138 -532
rect 190206 -588 190262 -532
rect 194908 20402 194964 20458
rect 201740 15722 201796 15778
rect 203644 10862 203700 10918
rect 216748 61082 216804 61138
rect 215068 37502 215124 37558
rect 209356 7262 209412 7318
rect 224274 598116 224330 598172
rect 224398 598116 224454 598172
rect 224522 598116 224578 598172
rect 224646 598116 224702 598172
rect 224274 597992 224330 598048
rect 224398 597992 224454 598048
rect 224522 597992 224578 598048
rect 224646 597992 224702 598048
rect 224274 597868 224330 597924
rect 224398 597868 224454 597924
rect 224522 597868 224578 597924
rect 224646 597868 224702 597924
rect 224274 597744 224330 597800
rect 224398 597744 224454 597800
rect 224522 597744 224578 597800
rect 224646 597744 224702 597800
rect 224274 586294 224330 586350
rect 224398 586294 224454 586350
rect 224522 586294 224578 586350
rect 224646 586294 224702 586350
rect 224274 586170 224330 586226
rect 224398 586170 224454 586226
rect 224522 586170 224578 586226
rect 224646 586170 224702 586226
rect 224274 586046 224330 586102
rect 224398 586046 224454 586102
rect 224522 586046 224578 586102
rect 224646 586046 224702 586102
rect 224274 585922 224330 585978
rect 224398 585922 224454 585978
rect 224522 585922 224578 585978
rect 224646 585922 224702 585978
rect 224274 568294 224330 568350
rect 224398 568294 224454 568350
rect 224522 568294 224578 568350
rect 224646 568294 224702 568350
rect 224274 568170 224330 568226
rect 224398 568170 224454 568226
rect 224522 568170 224578 568226
rect 224646 568170 224702 568226
rect 224274 568046 224330 568102
rect 224398 568046 224454 568102
rect 224522 568046 224578 568102
rect 224646 568046 224702 568102
rect 224274 567922 224330 567978
rect 224398 567922 224454 567978
rect 224522 567922 224578 567978
rect 224646 567922 224702 567978
rect 224274 550294 224330 550350
rect 224398 550294 224454 550350
rect 224522 550294 224578 550350
rect 224646 550294 224702 550350
rect 224274 550170 224330 550226
rect 224398 550170 224454 550226
rect 224522 550170 224578 550226
rect 224646 550170 224702 550226
rect 224274 550046 224330 550102
rect 224398 550046 224454 550102
rect 224522 550046 224578 550102
rect 224646 550046 224702 550102
rect 224274 549922 224330 549978
rect 224398 549922 224454 549978
rect 224522 549922 224578 549978
rect 224646 549922 224702 549978
rect 224274 532294 224330 532350
rect 224398 532294 224454 532350
rect 224522 532294 224578 532350
rect 224646 532294 224702 532350
rect 224274 532170 224330 532226
rect 224398 532170 224454 532226
rect 224522 532170 224578 532226
rect 224646 532170 224702 532226
rect 224274 532046 224330 532102
rect 224398 532046 224454 532102
rect 224522 532046 224578 532102
rect 224646 532046 224702 532102
rect 224274 531922 224330 531978
rect 224398 531922 224454 531978
rect 224522 531922 224578 531978
rect 224646 531922 224702 531978
rect 224274 514294 224330 514350
rect 224398 514294 224454 514350
rect 224522 514294 224578 514350
rect 224646 514294 224702 514350
rect 224274 514170 224330 514226
rect 224398 514170 224454 514226
rect 224522 514170 224578 514226
rect 224646 514170 224702 514226
rect 224274 514046 224330 514102
rect 224398 514046 224454 514102
rect 224522 514046 224578 514102
rect 224646 514046 224702 514102
rect 224274 513922 224330 513978
rect 224398 513922 224454 513978
rect 224522 513922 224578 513978
rect 224646 513922 224702 513978
rect 224274 496294 224330 496350
rect 224398 496294 224454 496350
rect 224522 496294 224578 496350
rect 224646 496294 224702 496350
rect 224274 496170 224330 496226
rect 224398 496170 224454 496226
rect 224522 496170 224578 496226
rect 224646 496170 224702 496226
rect 224274 496046 224330 496102
rect 224398 496046 224454 496102
rect 224522 496046 224578 496102
rect 224646 496046 224702 496102
rect 224274 495922 224330 495978
rect 224398 495922 224454 495978
rect 224522 495922 224578 495978
rect 224646 495922 224702 495978
rect 224274 478294 224330 478350
rect 224398 478294 224454 478350
rect 224522 478294 224578 478350
rect 224646 478294 224702 478350
rect 224274 478170 224330 478226
rect 224398 478170 224454 478226
rect 224522 478170 224578 478226
rect 224646 478170 224702 478226
rect 224274 478046 224330 478102
rect 224398 478046 224454 478102
rect 224522 478046 224578 478102
rect 224646 478046 224702 478102
rect 224274 477922 224330 477978
rect 224398 477922 224454 477978
rect 224522 477922 224578 477978
rect 224646 477922 224702 477978
rect 224274 460294 224330 460350
rect 224398 460294 224454 460350
rect 224522 460294 224578 460350
rect 224646 460294 224702 460350
rect 224274 460170 224330 460226
rect 224398 460170 224454 460226
rect 224522 460170 224578 460226
rect 224646 460170 224702 460226
rect 224274 460046 224330 460102
rect 224398 460046 224454 460102
rect 224522 460046 224578 460102
rect 224646 460046 224702 460102
rect 224274 459922 224330 459978
rect 224398 459922 224454 459978
rect 224522 459922 224578 459978
rect 224646 459922 224702 459978
rect 224274 442294 224330 442350
rect 224398 442294 224454 442350
rect 224522 442294 224578 442350
rect 224646 442294 224702 442350
rect 224274 442170 224330 442226
rect 224398 442170 224454 442226
rect 224522 442170 224578 442226
rect 224646 442170 224702 442226
rect 224274 442046 224330 442102
rect 224398 442046 224454 442102
rect 224522 442046 224578 442102
rect 224646 442046 224702 442102
rect 224274 441922 224330 441978
rect 224398 441922 224454 441978
rect 224522 441922 224578 441978
rect 224646 441922 224702 441978
rect 224274 424294 224330 424350
rect 224398 424294 224454 424350
rect 224522 424294 224578 424350
rect 224646 424294 224702 424350
rect 224274 424170 224330 424226
rect 224398 424170 224454 424226
rect 224522 424170 224578 424226
rect 224646 424170 224702 424226
rect 224274 424046 224330 424102
rect 224398 424046 224454 424102
rect 224522 424046 224578 424102
rect 224646 424046 224702 424102
rect 224274 423922 224330 423978
rect 224398 423922 224454 423978
rect 224522 423922 224578 423978
rect 224646 423922 224702 423978
rect 224274 406294 224330 406350
rect 224398 406294 224454 406350
rect 224522 406294 224578 406350
rect 224646 406294 224702 406350
rect 224274 406170 224330 406226
rect 224398 406170 224454 406226
rect 224522 406170 224578 406226
rect 224646 406170 224702 406226
rect 224274 406046 224330 406102
rect 224398 406046 224454 406102
rect 224522 406046 224578 406102
rect 224646 406046 224702 406102
rect 224274 405922 224330 405978
rect 224398 405922 224454 405978
rect 224522 405922 224578 405978
rect 224646 405922 224702 405978
rect 224274 388294 224330 388350
rect 224398 388294 224454 388350
rect 224522 388294 224578 388350
rect 224646 388294 224702 388350
rect 224274 388170 224330 388226
rect 224398 388170 224454 388226
rect 224522 388170 224578 388226
rect 224646 388170 224702 388226
rect 224274 388046 224330 388102
rect 224398 388046 224454 388102
rect 224522 388046 224578 388102
rect 224646 388046 224702 388102
rect 224274 387922 224330 387978
rect 224398 387922 224454 387978
rect 224522 387922 224578 387978
rect 224646 387922 224702 387978
rect 224274 370294 224330 370350
rect 224398 370294 224454 370350
rect 224522 370294 224578 370350
rect 224646 370294 224702 370350
rect 224274 370170 224330 370226
rect 224398 370170 224454 370226
rect 224522 370170 224578 370226
rect 224646 370170 224702 370226
rect 224274 370046 224330 370102
rect 224398 370046 224454 370102
rect 224522 370046 224578 370102
rect 224646 370046 224702 370102
rect 224274 369922 224330 369978
rect 224398 369922 224454 369978
rect 224522 369922 224578 369978
rect 224646 369922 224702 369978
rect 224274 352294 224330 352350
rect 224398 352294 224454 352350
rect 224522 352294 224578 352350
rect 224646 352294 224702 352350
rect 224274 352170 224330 352226
rect 224398 352170 224454 352226
rect 224522 352170 224578 352226
rect 224646 352170 224702 352226
rect 224274 352046 224330 352102
rect 224398 352046 224454 352102
rect 224522 352046 224578 352102
rect 224646 352046 224702 352102
rect 224274 351922 224330 351978
rect 224398 351922 224454 351978
rect 224522 351922 224578 351978
rect 224646 351922 224702 351978
rect 224274 334294 224330 334350
rect 224398 334294 224454 334350
rect 224522 334294 224578 334350
rect 224646 334294 224702 334350
rect 224274 334170 224330 334226
rect 224398 334170 224454 334226
rect 224522 334170 224578 334226
rect 224646 334170 224702 334226
rect 224274 334046 224330 334102
rect 224398 334046 224454 334102
rect 224522 334046 224578 334102
rect 224646 334046 224702 334102
rect 224274 333922 224330 333978
rect 224398 333922 224454 333978
rect 224522 333922 224578 333978
rect 224646 333922 224702 333978
rect 224274 316294 224330 316350
rect 224398 316294 224454 316350
rect 224522 316294 224578 316350
rect 224646 316294 224702 316350
rect 224274 316170 224330 316226
rect 224398 316170 224454 316226
rect 224522 316170 224578 316226
rect 224646 316170 224702 316226
rect 224274 316046 224330 316102
rect 224398 316046 224454 316102
rect 224522 316046 224578 316102
rect 224646 316046 224702 316102
rect 224274 315922 224330 315978
rect 224398 315922 224454 315978
rect 224522 315922 224578 315978
rect 224646 315922 224702 315978
rect 224274 298294 224330 298350
rect 224398 298294 224454 298350
rect 224522 298294 224578 298350
rect 224646 298294 224702 298350
rect 224274 298170 224330 298226
rect 224398 298170 224454 298226
rect 224522 298170 224578 298226
rect 224646 298170 224702 298226
rect 224274 298046 224330 298102
rect 224398 298046 224454 298102
rect 224522 298046 224578 298102
rect 224646 298046 224702 298102
rect 224274 297922 224330 297978
rect 224398 297922 224454 297978
rect 224522 297922 224578 297978
rect 224646 297922 224702 297978
rect 224274 280294 224330 280350
rect 224398 280294 224454 280350
rect 224522 280294 224578 280350
rect 224646 280294 224702 280350
rect 224274 280170 224330 280226
rect 224398 280170 224454 280226
rect 224522 280170 224578 280226
rect 224646 280170 224702 280226
rect 224274 280046 224330 280102
rect 224398 280046 224454 280102
rect 224522 280046 224578 280102
rect 224646 280046 224702 280102
rect 224274 279922 224330 279978
rect 224398 279922 224454 279978
rect 224522 279922 224578 279978
rect 224646 279922 224702 279978
rect 224274 262294 224330 262350
rect 224398 262294 224454 262350
rect 224522 262294 224578 262350
rect 224646 262294 224702 262350
rect 224274 262170 224330 262226
rect 224398 262170 224454 262226
rect 224522 262170 224578 262226
rect 224646 262170 224702 262226
rect 224274 262046 224330 262102
rect 224398 262046 224454 262102
rect 224522 262046 224578 262102
rect 224646 262046 224702 262102
rect 224274 261922 224330 261978
rect 224398 261922 224454 261978
rect 224522 261922 224578 261978
rect 224646 261922 224702 261978
rect 224274 244294 224330 244350
rect 224398 244294 224454 244350
rect 224522 244294 224578 244350
rect 224646 244294 224702 244350
rect 224274 244170 224330 244226
rect 224398 244170 224454 244226
rect 224522 244170 224578 244226
rect 224646 244170 224702 244226
rect 224274 244046 224330 244102
rect 224398 244046 224454 244102
rect 224522 244046 224578 244102
rect 224646 244046 224702 244102
rect 224274 243922 224330 243978
rect 224398 243922 224454 243978
rect 224522 243922 224578 243978
rect 224646 243922 224702 243978
rect 224274 226294 224330 226350
rect 224398 226294 224454 226350
rect 224522 226294 224578 226350
rect 224646 226294 224702 226350
rect 224274 226170 224330 226226
rect 224398 226170 224454 226226
rect 224522 226170 224578 226226
rect 224646 226170 224702 226226
rect 224274 226046 224330 226102
rect 224398 226046 224454 226102
rect 224522 226046 224578 226102
rect 224646 226046 224702 226102
rect 224274 225922 224330 225978
rect 224398 225922 224454 225978
rect 224522 225922 224578 225978
rect 224646 225922 224702 225978
rect 224274 208294 224330 208350
rect 224398 208294 224454 208350
rect 224522 208294 224578 208350
rect 224646 208294 224702 208350
rect 224274 208170 224330 208226
rect 224398 208170 224454 208226
rect 224522 208170 224578 208226
rect 224646 208170 224702 208226
rect 224274 208046 224330 208102
rect 224398 208046 224454 208102
rect 224522 208046 224578 208102
rect 224646 208046 224702 208102
rect 224274 207922 224330 207978
rect 224398 207922 224454 207978
rect 224522 207922 224578 207978
rect 224646 207922 224702 207978
rect 224274 190294 224330 190350
rect 224398 190294 224454 190350
rect 224522 190294 224578 190350
rect 224646 190294 224702 190350
rect 224274 190170 224330 190226
rect 224398 190170 224454 190226
rect 224522 190170 224578 190226
rect 224646 190170 224702 190226
rect 224274 190046 224330 190102
rect 224398 190046 224454 190102
rect 224522 190046 224578 190102
rect 224646 190046 224702 190102
rect 224274 189922 224330 189978
rect 224398 189922 224454 189978
rect 224522 189922 224578 189978
rect 224646 189922 224702 189978
rect 224274 172294 224330 172350
rect 224398 172294 224454 172350
rect 224522 172294 224578 172350
rect 224646 172294 224702 172350
rect 224274 172170 224330 172226
rect 224398 172170 224454 172226
rect 224522 172170 224578 172226
rect 224646 172170 224702 172226
rect 224274 172046 224330 172102
rect 224398 172046 224454 172102
rect 224522 172046 224578 172102
rect 224646 172046 224702 172102
rect 224274 171922 224330 171978
rect 224398 171922 224454 171978
rect 224522 171922 224578 171978
rect 224646 171922 224702 171978
rect 224274 154294 224330 154350
rect 224398 154294 224454 154350
rect 224522 154294 224578 154350
rect 224646 154294 224702 154350
rect 224274 154170 224330 154226
rect 224398 154170 224454 154226
rect 224522 154170 224578 154226
rect 224646 154170 224702 154226
rect 224274 154046 224330 154102
rect 224398 154046 224454 154102
rect 224522 154046 224578 154102
rect 224646 154046 224702 154102
rect 224274 153922 224330 153978
rect 224398 153922 224454 153978
rect 224522 153922 224578 153978
rect 224646 153922 224702 153978
rect 224274 136294 224330 136350
rect 224398 136294 224454 136350
rect 224522 136294 224578 136350
rect 224646 136294 224702 136350
rect 224274 136170 224330 136226
rect 224398 136170 224454 136226
rect 224522 136170 224578 136226
rect 224646 136170 224702 136226
rect 224274 136046 224330 136102
rect 224398 136046 224454 136102
rect 224522 136046 224578 136102
rect 224646 136046 224702 136102
rect 224274 135922 224330 135978
rect 224398 135922 224454 135978
rect 224522 135922 224578 135978
rect 224646 135922 224702 135978
rect 224274 118294 224330 118350
rect 224398 118294 224454 118350
rect 224522 118294 224578 118350
rect 224646 118294 224702 118350
rect 224274 118170 224330 118226
rect 224398 118170 224454 118226
rect 224522 118170 224578 118226
rect 224646 118170 224702 118226
rect 224274 118046 224330 118102
rect 224398 118046 224454 118102
rect 224522 118046 224578 118102
rect 224646 118046 224702 118102
rect 224274 117922 224330 117978
rect 224398 117922 224454 117978
rect 224522 117922 224578 117978
rect 224646 117922 224702 117978
rect 224274 100294 224330 100350
rect 224398 100294 224454 100350
rect 224522 100294 224578 100350
rect 224646 100294 224702 100350
rect 224274 100170 224330 100226
rect 224398 100170 224454 100226
rect 224522 100170 224578 100226
rect 224646 100170 224702 100226
rect 224274 100046 224330 100102
rect 224398 100046 224454 100102
rect 224522 100046 224578 100102
rect 224646 100046 224702 100102
rect 224274 99922 224330 99978
rect 224398 99922 224454 99978
rect 224522 99922 224578 99978
rect 224646 99922 224702 99978
rect 224274 82294 224330 82350
rect 224398 82294 224454 82350
rect 224522 82294 224578 82350
rect 224646 82294 224702 82350
rect 224274 82170 224330 82226
rect 224398 82170 224454 82226
rect 224522 82170 224578 82226
rect 224646 82170 224702 82226
rect 224274 82046 224330 82102
rect 224398 82046 224454 82102
rect 224522 82046 224578 82102
rect 224646 82046 224702 82102
rect 224274 81922 224330 81978
rect 224398 81922 224454 81978
rect 224522 81922 224578 81978
rect 224646 81922 224702 81978
rect 220554 58294 220610 58350
rect 220678 58294 220734 58350
rect 220802 58294 220858 58350
rect 220926 58294 220982 58350
rect 220554 58170 220610 58226
rect 220678 58170 220734 58226
rect 220802 58170 220858 58226
rect 220926 58170 220982 58226
rect 220554 58046 220610 58102
rect 220678 58046 220734 58102
rect 220802 58046 220858 58102
rect 220926 58046 220982 58102
rect 220554 57922 220610 57978
rect 220678 57922 220734 57978
rect 220802 57922 220858 57978
rect 220926 57922 220982 57978
rect 220108 40922 220164 40978
rect 223468 67922 223524 67978
rect 220554 40294 220610 40350
rect 220678 40294 220734 40350
rect 220802 40294 220858 40350
rect 220926 40294 220982 40350
rect 220554 40170 220610 40226
rect 220678 40170 220734 40226
rect 220802 40170 220858 40226
rect 220926 40170 220982 40226
rect 220554 40046 220610 40102
rect 220678 40046 220734 40102
rect 220802 40046 220858 40102
rect 220926 40046 220982 40102
rect 220554 39922 220610 39978
rect 220678 39922 220734 39978
rect 220802 39922 220858 39978
rect 220926 39922 220982 39978
rect 220554 22294 220610 22350
rect 220678 22294 220734 22350
rect 220802 22294 220858 22350
rect 220926 22294 220982 22350
rect 220554 22170 220610 22226
rect 220678 22170 220734 22226
rect 220802 22170 220858 22226
rect 220926 22170 220982 22226
rect 220554 22046 220610 22102
rect 220678 22046 220734 22102
rect 220802 22046 220858 22102
rect 220926 22046 220982 22102
rect 220554 21922 220610 21978
rect 220678 21922 220734 21978
rect 220802 21922 220858 21978
rect 220926 21922 220982 21978
rect 220554 4294 220610 4350
rect 220678 4294 220734 4350
rect 220802 4294 220858 4350
rect 220926 4294 220982 4350
rect 220554 4170 220610 4226
rect 220678 4170 220734 4226
rect 220802 4170 220858 4226
rect 220926 4170 220982 4226
rect 221788 47582 221844 47638
rect 251274 597156 251330 597212
rect 251398 597156 251454 597212
rect 251522 597156 251578 597212
rect 251646 597156 251702 597212
rect 251274 597032 251330 597088
rect 251398 597032 251454 597088
rect 251522 597032 251578 597088
rect 251646 597032 251702 597088
rect 251274 596908 251330 596964
rect 251398 596908 251454 596964
rect 251522 596908 251578 596964
rect 251646 596908 251702 596964
rect 251274 596784 251330 596840
rect 251398 596784 251454 596840
rect 251522 596784 251578 596840
rect 251646 596784 251702 596840
rect 251274 580294 251330 580350
rect 251398 580294 251454 580350
rect 251522 580294 251578 580350
rect 251646 580294 251702 580350
rect 251274 580170 251330 580226
rect 251398 580170 251454 580226
rect 251522 580170 251578 580226
rect 251646 580170 251702 580226
rect 251274 580046 251330 580102
rect 251398 580046 251454 580102
rect 251522 580046 251578 580102
rect 251646 580046 251702 580102
rect 251274 579922 251330 579978
rect 251398 579922 251454 579978
rect 251522 579922 251578 579978
rect 251646 579922 251702 579978
rect 251274 562294 251330 562350
rect 251398 562294 251454 562350
rect 251522 562294 251578 562350
rect 251646 562294 251702 562350
rect 251274 562170 251330 562226
rect 251398 562170 251454 562226
rect 251522 562170 251578 562226
rect 251646 562170 251702 562226
rect 251274 562046 251330 562102
rect 251398 562046 251454 562102
rect 251522 562046 251578 562102
rect 251646 562046 251702 562102
rect 251274 561922 251330 561978
rect 251398 561922 251454 561978
rect 251522 561922 251578 561978
rect 251646 561922 251702 561978
rect 251274 544294 251330 544350
rect 251398 544294 251454 544350
rect 251522 544294 251578 544350
rect 251646 544294 251702 544350
rect 251274 544170 251330 544226
rect 251398 544170 251454 544226
rect 251522 544170 251578 544226
rect 251646 544170 251702 544226
rect 251274 544046 251330 544102
rect 251398 544046 251454 544102
rect 251522 544046 251578 544102
rect 251646 544046 251702 544102
rect 251274 543922 251330 543978
rect 251398 543922 251454 543978
rect 251522 543922 251578 543978
rect 251646 543922 251702 543978
rect 251274 526294 251330 526350
rect 251398 526294 251454 526350
rect 251522 526294 251578 526350
rect 251646 526294 251702 526350
rect 251274 526170 251330 526226
rect 251398 526170 251454 526226
rect 251522 526170 251578 526226
rect 251646 526170 251702 526226
rect 251274 526046 251330 526102
rect 251398 526046 251454 526102
rect 251522 526046 251578 526102
rect 251646 526046 251702 526102
rect 251274 525922 251330 525978
rect 251398 525922 251454 525978
rect 251522 525922 251578 525978
rect 251646 525922 251702 525978
rect 251274 508294 251330 508350
rect 251398 508294 251454 508350
rect 251522 508294 251578 508350
rect 251646 508294 251702 508350
rect 251274 508170 251330 508226
rect 251398 508170 251454 508226
rect 251522 508170 251578 508226
rect 251646 508170 251702 508226
rect 251274 508046 251330 508102
rect 251398 508046 251454 508102
rect 251522 508046 251578 508102
rect 251646 508046 251702 508102
rect 251274 507922 251330 507978
rect 251398 507922 251454 507978
rect 251522 507922 251578 507978
rect 251646 507922 251702 507978
rect 251274 490294 251330 490350
rect 251398 490294 251454 490350
rect 251522 490294 251578 490350
rect 251646 490294 251702 490350
rect 251274 490170 251330 490226
rect 251398 490170 251454 490226
rect 251522 490170 251578 490226
rect 251646 490170 251702 490226
rect 251274 490046 251330 490102
rect 251398 490046 251454 490102
rect 251522 490046 251578 490102
rect 251646 490046 251702 490102
rect 251274 489922 251330 489978
rect 251398 489922 251454 489978
rect 251522 489922 251578 489978
rect 251646 489922 251702 489978
rect 251274 472294 251330 472350
rect 251398 472294 251454 472350
rect 251522 472294 251578 472350
rect 251646 472294 251702 472350
rect 251274 472170 251330 472226
rect 251398 472170 251454 472226
rect 251522 472170 251578 472226
rect 251646 472170 251702 472226
rect 251274 472046 251330 472102
rect 251398 472046 251454 472102
rect 251522 472046 251578 472102
rect 251646 472046 251702 472102
rect 251274 471922 251330 471978
rect 251398 471922 251454 471978
rect 251522 471922 251578 471978
rect 251646 471922 251702 471978
rect 251274 454294 251330 454350
rect 251398 454294 251454 454350
rect 251522 454294 251578 454350
rect 251646 454294 251702 454350
rect 251274 454170 251330 454226
rect 251398 454170 251454 454226
rect 251522 454170 251578 454226
rect 251646 454170 251702 454226
rect 251274 454046 251330 454102
rect 251398 454046 251454 454102
rect 251522 454046 251578 454102
rect 251646 454046 251702 454102
rect 251274 453922 251330 453978
rect 251398 453922 251454 453978
rect 251522 453922 251578 453978
rect 251646 453922 251702 453978
rect 251274 436294 251330 436350
rect 251398 436294 251454 436350
rect 251522 436294 251578 436350
rect 251646 436294 251702 436350
rect 251274 436170 251330 436226
rect 251398 436170 251454 436226
rect 251522 436170 251578 436226
rect 251646 436170 251702 436226
rect 251274 436046 251330 436102
rect 251398 436046 251454 436102
rect 251522 436046 251578 436102
rect 251646 436046 251702 436102
rect 251274 435922 251330 435978
rect 251398 435922 251454 435978
rect 251522 435922 251578 435978
rect 251646 435922 251702 435978
rect 251274 418294 251330 418350
rect 251398 418294 251454 418350
rect 251522 418294 251578 418350
rect 251646 418294 251702 418350
rect 251274 418170 251330 418226
rect 251398 418170 251454 418226
rect 251522 418170 251578 418226
rect 251646 418170 251702 418226
rect 251274 418046 251330 418102
rect 251398 418046 251454 418102
rect 251522 418046 251578 418102
rect 251646 418046 251702 418102
rect 251274 417922 251330 417978
rect 251398 417922 251454 417978
rect 251522 417922 251578 417978
rect 251646 417922 251702 417978
rect 251274 400294 251330 400350
rect 251398 400294 251454 400350
rect 251522 400294 251578 400350
rect 251646 400294 251702 400350
rect 251274 400170 251330 400226
rect 251398 400170 251454 400226
rect 251522 400170 251578 400226
rect 251646 400170 251702 400226
rect 251274 400046 251330 400102
rect 251398 400046 251454 400102
rect 251522 400046 251578 400102
rect 251646 400046 251702 400102
rect 251274 399922 251330 399978
rect 251398 399922 251454 399978
rect 251522 399922 251578 399978
rect 251646 399922 251702 399978
rect 251274 382294 251330 382350
rect 251398 382294 251454 382350
rect 251522 382294 251578 382350
rect 251646 382294 251702 382350
rect 251274 382170 251330 382226
rect 251398 382170 251454 382226
rect 251522 382170 251578 382226
rect 251646 382170 251702 382226
rect 251274 382046 251330 382102
rect 251398 382046 251454 382102
rect 251522 382046 251578 382102
rect 251646 382046 251702 382102
rect 251274 381922 251330 381978
rect 251398 381922 251454 381978
rect 251522 381922 251578 381978
rect 251646 381922 251702 381978
rect 251274 364294 251330 364350
rect 251398 364294 251454 364350
rect 251522 364294 251578 364350
rect 251646 364294 251702 364350
rect 251274 364170 251330 364226
rect 251398 364170 251454 364226
rect 251522 364170 251578 364226
rect 251646 364170 251702 364226
rect 251274 364046 251330 364102
rect 251398 364046 251454 364102
rect 251522 364046 251578 364102
rect 251646 364046 251702 364102
rect 251274 363922 251330 363978
rect 251398 363922 251454 363978
rect 251522 363922 251578 363978
rect 251646 363922 251702 363978
rect 251274 346294 251330 346350
rect 251398 346294 251454 346350
rect 251522 346294 251578 346350
rect 251646 346294 251702 346350
rect 251274 346170 251330 346226
rect 251398 346170 251454 346226
rect 251522 346170 251578 346226
rect 251646 346170 251702 346226
rect 251274 346046 251330 346102
rect 251398 346046 251454 346102
rect 251522 346046 251578 346102
rect 251646 346046 251702 346102
rect 251274 345922 251330 345978
rect 251398 345922 251454 345978
rect 251522 345922 251578 345978
rect 251646 345922 251702 345978
rect 251274 328294 251330 328350
rect 251398 328294 251454 328350
rect 251522 328294 251578 328350
rect 251646 328294 251702 328350
rect 251274 328170 251330 328226
rect 251398 328170 251454 328226
rect 251522 328170 251578 328226
rect 251646 328170 251702 328226
rect 251274 328046 251330 328102
rect 251398 328046 251454 328102
rect 251522 328046 251578 328102
rect 251646 328046 251702 328102
rect 251274 327922 251330 327978
rect 251398 327922 251454 327978
rect 251522 327922 251578 327978
rect 251646 327922 251702 327978
rect 251274 310294 251330 310350
rect 251398 310294 251454 310350
rect 251522 310294 251578 310350
rect 251646 310294 251702 310350
rect 251274 310170 251330 310226
rect 251398 310170 251454 310226
rect 251522 310170 251578 310226
rect 251646 310170 251702 310226
rect 251274 310046 251330 310102
rect 251398 310046 251454 310102
rect 251522 310046 251578 310102
rect 251646 310046 251702 310102
rect 251274 309922 251330 309978
rect 251398 309922 251454 309978
rect 251522 309922 251578 309978
rect 251646 309922 251702 309978
rect 251274 292294 251330 292350
rect 251398 292294 251454 292350
rect 251522 292294 251578 292350
rect 251646 292294 251702 292350
rect 251274 292170 251330 292226
rect 251398 292170 251454 292226
rect 251522 292170 251578 292226
rect 251646 292170 251702 292226
rect 251274 292046 251330 292102
rect 251398 292046 251454 292102
rect 251522 292046 251578 292102
rect 251646 292046 251702 292102
rect 251274 291922 251330 291978
rect 251398 291922 251454 291978
rect 251522 291922 251578 291978
rect 251646 291922 251702 291978
rect 251274 274294 251330 274350
rect 251398 274294 251454 274350
rect 251522 274294 251578 274350
rect 251646 274294 251702 274350
rect 251274 274170 251330 274226
rect 251398 274170 251454 274226
rect 251522 274170 251578 274226
rect 251646 274170 251702 274226
rect 251274 274046 251330 274102
rect 251398 274046 251454 274102
rect 251522 274046 251578 274102
rect 251646 274046 251702 274102
rect 251274 273922 251330 273978
rect 251398 273922 251454 273978
rect 251522 273922 251578 273978
rect 251646 273922 251702 273978
rect 251274 256294 251330 256350
rect 251398 256294 251454 256350
rect 251522 256294 251578 256350
rect 251646 256294 251702 256350
rect 251274 256170 251330 256226
rect 251398 256170 251454 256226
rect 251522 256170 251578 256226
rect 251646 256170 251702 256226
rect 251274 256046 251330 256102
rect 251398 256046 251454 256102
rect 251522 256046 251578 256102
rect 251646 256046 251702 256102
rect 251274 255922 251330 255978
rect 251398 255922 251454 255978
rect 251522 255922 251578 255978
rect 251646 255922 251702 255978
rect 251274 238294 251330 238350
rect 251398 238294 251454 238350
rect 251522 238294 251578 238350
rect 251646 238294 251702 238350
rect 251274 238170 251330 238226
rect 251398 238170 251454 238226
rect 251522 238170 251578 238226
rect 251646 238170 251702 238226
rect 251274 238046 251330 238102
rect 251398 238046 251454 238102
rect 251522 238046 251578 238102
rect 251646 238046 251702 238102
rect 251274 237922 251330 237978
rect 251398 237922 251454 237978
rect 251522 237922 251578 237978
rect 251646 237922 251702 237978
rect 251274 220294 251330 220350
rect 251398 220294 251454 220350
rect 251522 220294 251578 220350
rect 251646 220294 251702 220350
rect 251274 220170 251330 220226
rect 251398 220170 251454 220226
rect 251522 220170 251578 220226
rect 251646 220170 251702 220226
rect 251274 220046 251330 220102
rect 251398 220046 251454 220102
rect 251522 220046 251578 220102
rect 251646 220046 251702 220102
rect 251274 219922 251330 219978
rect 251398 219922 251454 219978
rect 251522 219922 251578 219978
rect 251646 219922 251702 219978
rect 251274 202294 251330 202350
rect 251398 202294 251454 202350
rect 251522 202294 251578 202350
rect 251646 202294 251702 202350
rect 251274 202170 251330 202226
rect 251398 202170 251454 202226
rect 251522 202170 251578 202226
rect 251646 202170 251702 202226
rect 251274 202046 251330 202102
rect 251398 202046 251454 202102
rect 251522 202046 251578 202102
rect 251646 202046 251702 202102
rect 251274 201922 251330 201978
rect 251398 201922 251454 201978
rect 251522 201922 251578 201978
rect 251646 201922 251702 201978
rect 251274 184294 251330 184350
rect 251398 184294 251454 184350
rect 251522 184294 251578 184350
rect 251646 184294 251702 184350
rect 251274 184170 251330 184226
rect 251398 184170 251454 184226
rect 251522 184170 251578 184226
rect 251646 184170 251702 184226
rect 251274 184046 251330 184102
rect 251398 184046 251454 184102
rect 251522 184046 251578 184102
rect 251646 184046 251702 184102
rect 251274 183922 251330 183978
rect 251398 183922 251454 183978
rect 251522 183922 251578 183978
rect 251646 183922 251702 183978
rect 251274 166294 251330 166350
rect 251398 166294 251454 166350
rect 251522 166294 251578 166350
rect 251646 166294 251702 166350
rect 251274 166170 251330 166226
rect 251398 166170 251454 166226
rect 251522 166170 251578 166226
rect 251646 166170 251702 166226
rect 251274 166046 251330 166102
rect 251398 166046 251454 166102
rect 251522 166046 251578 166102
rect 251646 166046 251702 166102
rect 251274 165922 251330 165978
rect 251398 165922 251454 165978
rect 251522 165922 251578 165978
rect 251646 165922 251702 165978
rect 251274 148294 251330 148350
rect 251398 148294 251454 148350
rect 251522 148294 251578 148350
rect 251646 148294 251702 148350
rect 251274 148170 251330 148226
rect 251398 148170 251454 148226
rect 251522 148170 251578 148226
rect 251646 148170 251702 148226
rect 251274 148046 251330 148102
rect 251398 148046 251454 148102
rect 251522 148046 251578 148102
rect 251646 148046 251702 148102
rect 251274 147922 251330 147978
rect 251398 147922 251454 147978
rect 251522 147922 251578 147978
rect 251646 147922 251702 147978
rect 251274 130294 251330 130350
rect 251398 130294 251454 130350
rect 251522 130294 251578 130350
rect 251646 130294 251702 130350
rect 251274 130170 251330 130226
rect 251398 130170 251454 130226
rect 251522 130170 251578 130226
rect 251646 130170 251702 130226
rect 251274 130046 251330 130102
rect 251398 130046 251454 130102
rect 251522 130046 251578 130102
rect 251646 130046 251702 130102
rect 251274 129922 251330 129978
rect 251398 129922 251454 129978
rect 251522 129922 251578 129978
rect 251646 129922 251702 129978
rect 251274 112294 251330 112350
rect 251398 112294 251454 112350
rect 251522 112294 251578 112350
rect 251646 112294 251702 112350
rect 251274 112170 251330 112226
rect 251398 112170 251454 112226
rect 251522 112170 251578 112226
rect 251646 112170 251702 112226
rect 251274 112046 251330 112102
rect 251398 112046 251454 112102
rect 251522 112046 251578 112102
rect 251646 112046 251702 112102
rect 251274 111922 251330 111978
rect 251398 111922 251454 111978
rect 251522 111922 251578 111978
rect 251646 111922 251702 111978
rect 251274 94294 251330 94350
rect 251398 94294 251454 94350
rect 251522 94294 251578 94350
rect 251646 94294 251702 94350
rect 251274 94170 251330 94226
rect 251398 94170 251454 94226
rect 251522 94170 251578 94226
rect 251646 94170 251702 94226
rect 251274 94046 251330 94102
rect 251398 94046 251454 94102
rect 251522 94046 251578 94102
rect 251646 94046 251702 94102
rect 251274 93922 251330 93978
rect 251398 93922 251454 93978
rect 251522 93922 251578 93978
rect 251646 93922 251702 93978
rect 251274 76294 251330 76350
rect 251398 76294 251454 76350
rect 251522 76294 251578 76350
rect 251646 76294 251702 76350
rect 251274 76170 251330 76226
rect 251398 76170 251454 76226
rect 251522 76170 251578 76226
rect 251646 76170 251702 76226
rect 251274 76046 251330 76102
rect 251398 76046 251454 76102
rect 251522 76046 251578 76102
rect 251646 76046 251702 76102
rect 251274 75922 251330 75978
rect 251398 75922 251454 75978
rect 251522 75922 251578 75978
rect 251646 75922 251702 75978
rect 248668 71162 248724 71218
rect 238588 69362 238644 69418
rect 224274 64294 224330 64350
rect 224398 64294 224454 64350
rect 224522 64294 224578 64350
rect 224646 64294 224702 64350
rect 224274 64170 224330 64226
rect 224398 64170 224454 64226
rect 224522 64170 224578 64226
rect 224646 64170 224702 64226
rect 224274 64046 224330 64102
rect 224398 64046 224454 64102
rect 224522 64046 224578 64102
rect 224646 64046 224702 64102
rect 224274 63922 224330 63978
rect 224398 63922 224454 63978
rect 224522 63922 224578 63978
rect 224646 63922 224702 63978
rect 224274 46294 224330 46350
rect 224398 46294 224454 46350
rect 224522 46294 224578 46350
rect 224646 46294 224702 46350
rect 224274 46170 224330 46226
rect 224398 46170 224454 46226
rect 224522 46170 224578 46226
rect 224646 46170 224702 46226
rect 224274 46046 224330 46102
rect 224398 46046 224454 46102
rect 224522 46046 224578 46102
rect 224646 46046 224702 46102
rect 224274 45922 224330 45978
rect 224398 45922 224454 45978
rect 224522 45922 224578 45978
rect 224646 45922 224702 45978
rect 235228 66302 235284 66358
rect 231868 37322 231924 37378
rect 224274 28294 224330 28350
rect 224398 28294 224454 28350
rect 224522 28294 224578 28350
rect 224646 28294 224702 28350
rect 224274 28170 224330 28226
rect 224398 28170 224454 28226
rect 224522 28170 224578 28226
rect 224646 28170 224702 28226
rect 224274 28046 224330 28102
rect 224398 28046 224454 28102
rect 224522 28046 224578 28102
rect 224646 28046 224702 28102
rect 224274 27922 224330 27978
rect 224398 27922 224454 27978
rect 224522 27922 224578 27978
rect 224646 27922 224702 27978
rect 224274 10294 224330 10350
rect 224398 10294 224454 10350
rect 224522 10294 224578 10350
rect 224646 10294 224702 10350
rect 224274 10170 224330 10226
rect 224398 10170 224454 10226
rect 224522 10170 224578 10226
rect 224646 10170 224702 10226
rect 224274 10046 224330 10102
rect 224398 10046 224454 10102
rect 224522 10046 224578 10102
rect 224646 10046 224702 10102
rect 224274 9922 224330 9978
rect 224398 9922 224454 9978
rect 224522 9922 224578 9978
rect 224646 9922 224702 9978
rect 220554 4046 220610 4102
rect 220678 4046 220734 4102
rect 220802 4046 220858 4102
rect 220926 4046 220982 4102
rect 220554 3922 220610 3978
rect 220678 3922 220734 3978
rect 220802 3922 220858 3978
rect 220926 3922 220982 3978
rect 197932 2942 197988 2998
rect 211260 62 211316 118
rect 193554 -1176 193610 -1120
rect 193678 -1176 193734 -1120
rect 193802 -1176 193858 -1120
rect 193926 -1176 193982 -1120
rect 193554 -1300 193610 -1244
rect 193678 -1300 193734 -1244
rect 193802 -1300 193858 -1244
rect 193926 -1300 193982 -1244
rect 193554 -1424 193610 -1368
rect 193678 -1424 193734 -1368
rect 193802 -1424 193858 -1368
rect 193926 -1424 193982 -1368
rect 193554 -1548 193610 -1492
rect 193678 -1548 193734 -1492
rect 193802 -1548 193858 -1492
rect 193926 -1548 193982 -1492
rect 220554 -216 220610 -160
rect 220678 -216 220734 -160
rect 220802 -216 220858 -160
rect 220926 -216 220982 -160
rect 220554 -340 220610 -284
rect 220678 -340 220734 -284
rect 220802 -340 220858 -284
rect 220926 -340 220982 -284
rect 220554 -464 220610 -408
rect 220678 -464 220734 -408
rect 220802 -464 220858 -408
rect 220926 -464 220982 -408
rect 220554 -588 220610 -532
rect 220678 -588 220734 -532
rect 220802 -588 220858 -532
rect 220926 -588 220982 -532
rect 228508 36062 228564 36118
rect 233548 32282 233604 32338
rect 236908 25802 236964 25858
rect 243628 35882 243684 35938
rect 245532 18602 245588 18658
rect 254994 598116 255050 598172
rect 255118 598116 255174 598172
rect 255242 598116 255298 598172
rect 255366 598116 255422 598172
rect 254994 597992 255050 598048
rect 255118 597992 255174 598048
rect 255242 597992 255298 598048
rect 255366 597992 255422 598048
rect 254994 597868 255050 597924
rect 255118 597868 255174 597924
rect 255242 597868 255298 597924
rect 255366 597868 255422 597924
rect 254994 597744 255050 597800
rect 255118 597744 255174 597800
rect 255242 597744 255298 597800
rect 255366 597744 255422 597800
rect 254994 586294 255050 586350
rect 255118 586294 255174 586350
rect 255242 586294 255298 586350
rect 255366 586294 255422 586350
rect 254994 586170 255050 586226
rect 255118 586170 255174 586226
rect 255242 586170 255298 586226
rect 255366 586170 255422 586226
rect 254994 586046 255050 586102
rect 255118 586046 255174 586102
rect 255242 586046 255298 586102
rect 255366 586046 255422 586102
rect 254994 585922 255050 585978
rect 255118 585922 255174 585978
rect 255242 585922 255298 585978
rect 255366 585922 255422 585978
rect 254994 568294 255050 568350
rect 255118 568294 255174 568350
rect 255242 568294 255298 568350
rect 255366 568294 255422 568350
rect 254994 568170 255050 568226
rect 255118 568170 255174 568226
rect 255242 568170 255298 568226
rect 255366 568170 255422 568226
rect 254994 568046 255050 568102
rect 255118 568046 255174 568102
rect 255242 568046 255298 568102
rect 255366 568046 255422 568102
rect 254994 567922 255050 567978
rect 255118 567922 255174 567978
rect 255242 567922 255298 567978
rect 255366 567922 255422 567978
rect 254994 550294 255050 550350
rect 255118 550294 255174 550350
rect 255242 550294 255298 550350
rect 255366 550294 255422 550350
rect 254994 550170 255050 550226
rect 255118 550170 255174 550226
rect 255242 550170 255298 550226
rect 255366 550170 255422 550226
rect 254994 550046 255050 550102
rect 255118 550046 255174 550102
rect 255242 550046 255298 550102
rect 255366 550046 255422 550102
rect 254994 549922 255050 549978
rect 255118 549922 255174 549978
rect 255242 549922 255298 549978
rect 255366 549922 255422 549978
rect 254994 532294 255050 532350
rect 255118 532294 255174 532350
rect 255242 532294 255298 532350
rect 255366 532294 255422 532350
rect 254994 532170 255050 532226
rect 255118 532170 255174 532226
rect 255242 532170 255298 532226
rect 255366 532170 255422 532226
rect 254994 532046 255050 532102
rect 255118 532046 255174 532102
rect 255242 532046 255298 532102
rect 255366 532046 255422 532102
rect 254994 531922 255050 531978
rect 255118 531922 255174 531978
rect 255242 531922 255298 531978
rect 255366 531922 255422 531978
rect 254994 514294 255050 514350
rect 255118 514294 255174 514350
rect 255242 514294 255298 514350
rect 255366 514294 255422 514350
rect 254994 514170 255050 514226
rect 255118 514170 255174 514226
rect 255242 514170 255298 514226
rect 255366 514170 255422 514226
rect 254994 514046 255050 514102
rect 255118 514046 255174 514102
rect 255242 514046 255298 514102
rect 255366 514046 255422 514102
rect 254994 513922 255050 513978
rect 255118 513922 255174 513978
rect 255242 513922 255298 513978
rect 255366 513922 255422 513978
rect 254994 496294 255050 496350
rect 255118 496294 255174 496350
rect 255242 496294 255298 496350
rect 255366 496294 255422 496350
rect 254994 496170 255050 496226
rect 255118 496170 255174 496226
rect 255242 496170 255298 496226
rect 255366 496170 255422 496226
rect 254994 496046 255050 496102
rect 255118 496046 255174 496102
rect 255242 496046 255298 496102
rect 255366 496046 255422 496102
rect 254994 495922 255050 495978
rect 255118 495922 255174 495978
rect 255242 495922 255298 495978
rect 255366 495922 255422 495978
rect 254994 478294 255050 478350
rect 255118 478294 255174 478350
rect 255242 478294 255298 478350
rect 255366 478294 255422 478350
rect 254994 478170 255050 478226
rect 255118 478170 255174 478226
rect 255242 478170 255298 478226
rect 255366 478170 255422 478226
rect 254994 478046 255050 478102
rect 255118 478046 255174 478102
rect 255242 478046 255298 478102
rect 255366 478046 255422 478102
rect 254994 477922 255050 477978
rect 255118 477922 255174 477978
rect 255242 477922 255298 477978
rect 255366 477922 255422 477978
rect 254994 460294 255050 460350
rect 255118 460294 255174 460350
rect 255242 460294 255298 460350
rect 255366 460294 255422 460350
rect 254994 460170 255050 460226
rect 255118 460170 255174 460226
rect 255242 460170 255298 460226
rect 255366 460170 255422 460226
rect 254994 460046 255050 460102
rect 255118 460046 255174 460102
rect 255242 460046 255298 460102
rect 255366 460046 255422 460102
rect 254994 459922 255050 459978
rect 255118 459922 255174 459978
rect 255242 459922 255298 459978
rect 255366 459922 255422 459978
rect 254994 442294 255050 442350
rect 255118 442294 255174 442350
rect 255242 442294 255298 442350
rect 255366 442294 255422 442350
rect 254994 442170 255050 442226
rect 255118 442170 255174 442226
rect 255242 442170 255298 442226
rect 255366 442170 255422 442226
rect 254994 442046 255050 442102
rect 255118 442046 255174 442102
rect 255242 442046 255298 442102
rect 255366 442046 255422 442102
rect 254994 441922 255050 441978
rect 255118 441922 255174 441978
rect 255242 441922 255298 441978
rect 255366 441922 255422 441978
rect 254994 424294 255050 424350
rect 255118 424294 255174 424350
rect 255242 424294 255298 424350
rect 255366 424294 255422 424350
rect 254994 424170 255050 424226
rect 255118 424170 255174 424226
rect 255242 424170 255298 424226
rect 255366 424170 255422 424226
rect 254994 424046 255050 424102
rect 255118 424046 255174 424102
rect 255242 424046 255298 424102
rect 255366 424046 255422 424102
rect 254994 423922 255050 423978
rect 255118 423922 255174 423978
rect 255242 423922 255298 423978
rect 255366 423922 255422 423978
rect 254994 406294 255050 406350
rect 255118 406294 255174 406350
rect 255242 406294 255298 406350
rect 255366 406294 255422 406350
rect 254994 406170 255050 406226
rect 255118 406170 255174 406226
rect 255242 406170 255298 406226
rect 255366 406170 255422 406226
rect 254994 406046 255050 406102
rect 255118 406046 255174 406102
rect 255242 406046 255298 406102
rect 255366 406046 255422 406102
rect 254994 405922 255050 405978
rect 255118 405922 255174 405978
rect 255242 405922 255298 405978
rect 255366 405922 255422 405978
rect 254994 388294 255050 388350
rect 255118 388294 255174 388350
rect 255242 388294 255298 388350
rect 255366 388294 255422 388350
rect 254994 388170 255050 388226
rect 255118 388170 255174 388226
rect 255242 388170 255298 388226
rect 255366 388170 255422 388226
rect 254994 388046 255050 388102
rect 255118 388046 255174 388102
rect 255242 388046 255298 388102
rect 255366 388046 255422 388102
rect 254994 387922 255050 387978
rect 255118 387922 255174 387978
rect 255242 387922 255298 387978
rect 255366 387922 255422 387978
rect 254994 370294 255050 370350
rect 255118 370294 255174 370350
rect 255242 370294 255298 370350
rect 255366 370294 255422 370350
rect 254994 370170 255050 370226
rect 255118 370170 255174 370226
rect 255242 370170 255298 370226
rect 255366 370170 255422 370226
rect 254994 370046 255050 370102
rect 255118 370046 255174 370102
rect 255242 370046 255298 370102
rect 255366 370046 255422 370102
rect 254994 369922 255050 369978
rect 255118 369922 255174 369978
rect 255242 369922 255298 369978
rect 255366 369922 255422 369978
rect 254994 352294 255050 352350
rect 255118 352294 255174 352350
rect 255242 352294 255298 352350
rect 255366 352294 255422 352350
rect 254994 352170 255050 352226
rect 255118 352170 255174 352226
rect 255242 352170 255298 352226
rect 255366 352170 255422 352226
rect 254994 352046 255050 352102
rect 255118 352046 255174 352102
rect 255242 352046 255298 352102
rect 255366 352046 255422 352102
rect 254994 351922 255050 351978
rect 255118 351922 255174 351978
rect 255242 351922 255298 351978
rect 255366 351922 255422 351978
rect 254994 334294 255050 334350
rect 255118 334294 255174 334350
rect 255242 334294 255298 334350
rect 255366 334294 255422 334350
rect 254994 334170 255050 334226
rect 255118 334170 255174 334226
rect 255242 334170 255298 334226
rect 255366 334170 255422 334226
rect 254994 334046 255050 334102
rect 255118 334046 255174 334102
rect 255242 334046 255298 334102
rect 255366 334046 255422 334102
rect 254994 333922 255050 333978
rect 255118 333922 255174 333978
rect 255242 333922 255298 333978
rect 255366 333922 255422 333978
rect 254994 316294 255050 316350
rect 255118 316294 255174 316350
rect 255242 316294 255298 316350
rect 255366 316294 255422 316350
rect 254994 316170 255050 316226
rect 255118 316170 255174 316226
rect 255242 316170 255298 316226
rect 255366 316170 255422 316226
rect 254994 316046 255050 316102
rect 255118 316046 255174 316102
rect 255242 316046 255298 316102
rect 255366 316046 255422 316102
rect 254994 315922 255050 315978
rect 255118 315922 255174 315978
rect 255242 315922 255298 315978
rect 255366 315922 255422 315978
rect 254994 298294 255050 298350
rect 255118 298294 255174 298350
rect 255242 298294 255298 298350
rect 255366 298294 255422 298350
rect 254994 298170 255050 298226
rect 255118 298170 255174 298226
rect 255242 298170 255298 298226
rect 255366 298170 255422 298226
rect 254994 298046 255050 298102
rect 255118 298046 255174 298102
rect 255242 298046 255298 298102
rect 255366 298046 255422 298102
rect 254994 297922 255050 297978
rect 255118 297922 255174 297978
rect 255242 297922 255298 297978
rect 255366 297922 255422 297978
rect 254994 280294 255050 280350
rect 255118 280294 255174 280350
rect 255242 280294 255298 280350
rect 255366 280294 255422 280350
rect 254994 280170 255050 280226
rect 255118 280170 255174 280226
rect 255242 280170 255298 280226
rect 255366 280170 255422 280226
rect 254994 280046 255050 280102
rect 255118 280046 255174 280102
rect 255242 280046 255298 280102
rect 255366 280046 255422 280102
rect 254994 279922 255050 279978
rect 255118 279922 255174 279978
rect 255242 279922 255298 279978
rect 255366 279922 255422 279978
rect 254994 262294 255050 262350
rect 255118 262294 255174 262350
rect 255242 262294 255298 262350
rect 255366 262294 255422 262350
rect 254994 262170 255050 262226
rect 255118 262170 255174 262226
rect 255242 262170 255298 262226
rect 255366 262170 255422 262226
rect 254994 262046 255050 262102
rect 255118 262046 255174 262102
rect 255242 262046 255298 262102
rect 255366 262046 255422 262102
rect 254994 261922 255050 261978
rect 255118 261922 255174 261978
rect 255242 261922 255298 261978
rect 255366 261922 255422 261978
rect 254994 244294 255050 244350
rect 255118 244294 255174 244350
rect 255242 244294 255298 244350
rect 255366 244294 255422 244350
rect 254994 244170 255050 244226
rect 255118 244170 255174 244226
rect 255242 244170 255298 244226
rect 255366 244170 255422 244226
rect 254994 244046 255050 244102
rect 255118 244046 255174 244102
rect 255242 244046 255298 244102
rect 255366 244046 255422 244102
rect 254994 243922 255050 243978
rect 255118 243922 255174 243978
rect 255242 243922 255298 243978
rect 255366 243922 255422 243978
rect 254994 226294 255050 226350
rect 255118 226294 255174 226350
rect 255242 226294 255298 226350
rect 255366 226294 255422 226350
rect 254994 226170 255050 226226
rect 255118 226170 255174 226226
rect 255242 226170 255298 226226
rect 255366 226170 255422 226226
rect 254994 226046 255050 226102
rect 255118 226046 255174 226102
rect 255242 226046 255298 226102
rect 255366 226046 255422 226102
rect 254994 225922 255050 225978
rect 255118 225922 255174 225978
rect 255242 225922 255298 225978
rect 255366 225922 255422 225978
rect 254994 208294 255050 208350
rect 255118 208294 255174 208350
rect 255242 208294 255298 208350
rect 255366 208294 255422 208350
rect 254994 208170 255050 208226
rect 255118 208170 255174 208226
rect 255242 208170 255298 208226
rect 255366 208170 255422 208226
rect 254994 208046 255050 208102
rect 255118 208046 255174 208102
rect 255242 208046 255298 208102
rect 255366 208046 255422 208102
rect 254994 207922 255050 207978
rect 255118 207922 255174 207978
rect 255242 207922 255298 207978
rect 255366 207922 255422 207978
rect 254994 190294 255050 190350
rect 255118 190294 255174 190350
rect 255242 190294 255298 190350
rect 255366 190294 255422 190350
rect 254994 190170 255050 190226
rect 255118 190170 255174 190226
rect 255242 190170 255298 190226
rect 255366 190170 255422 190226
rect 254994 190046 255050 190102
rect 255118 190046 255174 190102
rect 255242 190046 255298 190102
rect 255366 190046 255422 190102
rect 254994 189922 255050 189978
rect 255118 189922 255174 189978
rect 255242 189922 255298 189978
rect 255366 189922 255422 189978
rect 254994 172294 255050 172350
rect 255118 172294 255174 172350
rect 255242 172294 255298 172350
rect 255366 172294 255422 172350
rect 254994 172170 255050 172226
rect 255118 172170 255174 172226
rect 255242 172170 255298 172226
rect 255366 172170 255422 172226
rect 254994 172046 255050 172102
rect 255118 172046 255174 172102
rect 255242 172046 255298 172102
rect 255366 172046 255422 172102
rect 254994 171922 255050 171978
rect 255118 171922 255174 171978
rect 255242 171922 255298 171978
rect 255366 171922 255422 171978
rect 254994 154294 255050 154350
rect 255118 154294 255174 154350
rect 255242 154294 255298 154350
rect 255366 154294 255422 154350
rect 254994 154170 255050 154226
rect 255118 154170 255174 154226
rect 255242 154170 255298 154226
rect 255366 154170 255422 154226
rect 254994 154046 255050 154102
rect 255118 154046 255174 154102
rect 255242 154046 255298 154102
rect 255366 154046 255422 154102
rect 254994 153922 255050 153978
rect 255118 153922 255174 153978
rect 255242 153922 255298 153978
rect 255366 153922 255422 153978
rect 254994 136294 255050 136350
rect 255118 136294 255174 136350
rect 255242 136294 255298 136350
rect 255366 136294 255422 136350
rect 254994 136170 255050 136226
rect 255118 136170 255174 136226
rect 255242 136170 255298 136226
rect 255366 136170 255422 136226
rect 254994 136046 255050 136102
rect 255118 136046 255174 136102
rect 255242 136046 255298 136102
rect 255366 136046 255422 136102
rect 254994 135922 255050 135978
rect 255118 135922 255174 135978
rect 255242 135922 255298 135978
rect 255366 135922 255422 135978
rect 254994 118294 255050 118350
rect 255118 118294 255174 118350
rect 255242 118294 255298 118350
rect 255366 118294 255422 118350
rect 254994 118170 255050 118226
rect 255118 118170 255174 118226
rect 255242 118170 255298 118226
rect 255366 118170 255422 118226
rect 254994 118046 255050 118102
rect 255118 118046 255174 118102
rect 255242 118046 255298 118102
rect 255366 118046 255422 118102
rect 254994 117922 255050 117978
rect 255118 117922 255174 117978
rect 255242 117922 255298 117978
rect 255366 117922 255422 117978
rect 254994 100294 255050 100350
rect 255118 100294 255174 100350
rect 255242 100294 255298 100350
rect 255366 100294 255422 100350
rect 254994 100170 255050 100226
rect 255118 100170 255174 100226
rect 255242 100170 255298 100226
rect 255366 100170 255422 100226
rect 254994 100046 255050 100102
rect 255118 100046 255174 100102
rect 255242 100046 255298 100102
rect 255366 100046 255422 100102
rect 254994 99922 255050 99978
rect 255118 99922 255174 99978
rect 255242 99922 255298 99978
rect 255366 99922 255422 99978
rect 254994 82294 255050 82350
rect 255118 82294 255174 82350
rect 255242 82294 255298 82350
rect 255366 82294 255422 82350
rect 254994 82170 255050 82226
rect 255118 82170 255174 82226
rect 255242 82170 255298 82226
rect 255366 82170 255422 82226
rect 254994 82046 255050 82102
rect 255118 82046 255174 82102
rect 255242 82046 255298 82102
rect 255366 82046 255422 82102
rect 254994 81922 255050 81978
rect 255118 81922 255174 81978
rect 255242 81922 255298 81978
rect 255366 81922 255422 81978
rect 251274 58294 251330 58350
rect 251398 58294 251454 58350
rect 251522 58294 251578 58350
rect 251646 58294 251702 58350
rect 251274 58170 251330 58226
rect 251398 58170 251454 58226
rect 251522 58170 251578 58226
rect 251646 58170 251702 58226
rect 251274 58046 251330 58102
rect 251398 58046 251454 58102
rect 251522 58046 251578 58102
rect 251646 58046 251702 58102
rect 251274 57922 251330 57978
rect 251398 57922 251454 57978
rect 251522 57922 251578 57978
rect 251646 57922 251702 57978
rect 251274 40294 251330 40350
rect 251398 40294 251454 40350
rect 251522 40294 251578 40350
rect 251646 40294 251702 40350
rect 251274 40170 251330 40226
rect 251398 40170 251454 40226
rect 251522 40170 251578 40226
rect 251646 40170 251702 40226
rect 251274 40046 251330 40102
rect 251398 40046 251454 40102
rect 251522 40046 251578 40102
rect 251646 40046 251702 40102
rect 251274 39922 251330 39978
rect 251398 39922 251454 39978
rect 251522 39922 251578 39978
rect 251646 39922 251702 39978
rect 251274 22294 251330 22350
rect 251398 22294 251454 22350
rect 251522 22294 251578 22350
rect 251646 22294 251702 22350
rect 251274 22170 251330 22226
rect 251398 22170 251454 22226
rect 251522 22170 251578 22226
rect 251646 22170 251702 22226
rect 251274 22046 251330 22102
rect 251398 22046 251454 22102
rect 251522 22046 251578 22102
rect 251646 22046 251702 22102
rect 251274 21922 251330 21978
rect 251398 21922 251454 21978
rect 251522 21922 251578 21978
rect 251646 21922 251702 21978
rect 250348 13742 250404 13798
rect 251274 4294 251330 4350
rect 251398 4294 251454 4350
rect 251522 4294 251578 4350
rect 251646 4294 251702 4350
rect 251274 4170 251330 4226
rect 251398 4170 251454 4226
rect 251522 4170 251578 4226
rect 251646 4170 251702 4226
rect 224274 -1176 224330 -1120
rect 224398 -1176 224454 -1120
rect 224522 -1176 224578 -1120
rect 224646 -1176 224702 -1120
rect 224274 -1300 224330 -1244
rect 224398 -1300 224454 -1244
rect 224522 -1300 224578 -1244
rect 224646 -1300 224702 -1244
rect 224274 -1424 224330 -1368
rect 224398 -1424 224454 -1368
rect 224522 -1424 224578 -1368
rect 224646 -1424 224702 -1368
rect 224274 -1548 224330 -1492
rect 224398 -1548 224454 -1492
rect 224522 -1548 224578 -1492
rect 224646 -1548 224702 -1492
rect 252028 64862 252084 64918
rect 253708 64682 253764 64738
rect 281994 597156 282050 597212
rect 282118 597156 282174 597212
rect 282242 597156 282298 597212
rect 282366 597156 282422 597212
rect 281994 597032 282050 597088
rect 282118 597032 282174 597088
rect 282242 597032 282298 597088
rect 282366 597032 282422 597088
rect 281994 596908 282050 596964
rect 282118 596908 282174 596964
rect 282242 596908 282298 596964
rect 282366 596908 282422 596964
rect 281994 596784 282050 596840
rect 282118 596784 282174 596840
rect 282242 596784 282298 596840
rect 282366 596784 282422 596840
rect 281994 580294 282050 580350
rect 282118 580294 282174 580350
rect 282242 580294 282298 580350
rect 282366 580294 282422 580350
rect 281994 580170 282050 580226
rect 282118 580170 282174 580226
rect 282242 580170 282298 580226
rect 282366 580170 282422 580226
rect 281994 580046 282050 580102
rect 282118 580046 282174 580102
rect 282242 580046 282298 580102
rect 282366 580046 282422 580102
rect 281994 579922 282050 579978
rect 282118 579922 282174 579978
rect 282242 579922 282298 579978
rect 282366 579922 282422 579978
rect 281994 562294 282050 562350
rect 282118 562294 282174 562350
rect 282242 562294 282298 562350
rect 282366 562294 282422 562350
rect 281994 562170 282050 562226
rect 282118 562170 282174 562226
rect 282242 562170 282298 562226
rect 282366 562170 282422 562226
rect 281994 562046 282050 562102
rect 282118 562046 282174 562102
rect 282242 562046 282298 562102
rect 282366 562046 282422 562102
rect 281994 561922 282050 561978
rect 282118 561922 282174 561978
rect 282242 561922 282298 561978
rect 282366 561922 282422 561978
rect 281994 544294 282050 544350
rect 282118 544294 282174 544350
rect 282242 544294 282298 544350
rect 282366 544294 282422 544350
rect 281994 544170 282050 544226
rect 282118 544170 282174 544226
rect 282242 544170 282298 544226
rect 282366 544170 282422 544226
rect 281994 544046 282050 544102
rect 282118 544046 282174 544102
rect 282242 544046 282298 544102
rect 282366 544046 282422 544102
rect 281994 543922 282050 543978
rect 282118 543922 282174 543978
rect 282242 543922 282298 543978
rect 282366 543922 282422 543978
rect 281994 526294 282050 526350
rect 282118 526294 282174 526350
rect 282242 526294 282298 526350
rect 282366 526294 282422 526350
rect 281994 526170 282050 526226
rect 282118 526170 282174 526226
rect 282242 526170 282298 526226
rect 282366 526170 282422 526226
rect 281994 526046 282050 526102
rect 282118 526046 282174 526102
rect 282242 526046 282298 526102
rect 282366 526046 282422 526102
rect 281994 525922 282050 525978
rect 282118 525922 282174 525978
rect 282242 525922 282298 525978
rect 282366 525922 282422 525978
rect 281994 508294 282050 508350
rect 282118 508294 282174 508350
rect 282242 508294 282298 508350
rect 282366 508294 282422 508350
rect 281994 508170 282050 508226
rect 282118 508170 282174 508226
rect 282242 508170 282298 508226
rect 282366 508170 282422 508226
rect 281994 508046 282050 508102
rect 282118 508046 282174 508102
rect 282242 508046 282298 508102
rect 282366 508046 282422 508102
rect 281994 507922 282050 507978
rect 282118 507922 282174 507978
rect 282242 507922 282298 507978
rect 282366 507922 282422 507978
rect 281994 490294 282050 490350
rect 282118 490294 282174 490350
rect 282242 490294 282298 490350
rect 282366 490294 282422 490350
rect 281994 490170 282050 490226
rect 282118 490170 282174 490226
rect 282242 490170 282298 490226
rect 282366 490170 282422 490226
rect 281994 490046 282050 490102
rect 282118 490046 282174 490102
rect 282242 490046 282298 490102
rect 282366 490046 282422 490102
rect 281994 489922 282050 489978
rect 282118 489922 282174 489978
rect 282242 489922 282298 489978
rect 282366 489922 282422 489978
rect 281994 472294 282050 472350
rect 282118 472294 282174 472350
rect 282242 472294 282298 472350
rect 282366 472294 282422 472350
rect 281994 472170 282050 472226
rect 282118 472170 282174 472226
rect 282242 472170 282298 472226
rect 282366 472170 282422 472226
rect 281994 472046 282050 472102
rect 282118 472046 282174 472102
rect 282242 472046 282298 472102
rect 282366 472046 282422 472102
rect 281994 471922 282050 471978
rect 282118 471922 282174 471978
rect 282242 471922 282298 471978
rect 282366 471922 282422 471978
rect 281994 454294 282050 454350
rect 282118 454294 282174 454350
rect 282242 454294 282298 454350
rect 282366 454294 282422 454350
rect 281994 454170 282050 454226
rect 282118 454170 282174 454226
rect 282242 454170 282298 454226
rect 282366 454170 282422 454226
rect 281994 454046 282050 454102
rect 282118 454046 282174 454102
rect 282242 454046 282298 454102
rect 282366 454046 282422 454102
rect 281994 453922 282050 453978
rect 282118 453922 282174 453978
rect 282242 453922 282298 453978
rect 282366 453922 282422 453978
rect 281994 436294 282050 436350
rect 282118 436294 282174 436350
rect 282242 436294 282298 436350
rect 282366 436294 282422 436350
rect 281994 436170 282050 436226
rect 282118 436170 282174 436226
rect 282242 436170 282298 436226
rect 282366 436170 282422 436226
rect 281994 436046 282050 436102
rect 282118 436046 282174 436102
rect 282242 436046 282298 436102
rect 282366 436046 282422 436102
rect 281994 435922 282050 435978
rect 282118 435922 282174 435978
rect 282242 435922 282298 435978
rect 282366 435922 282422 435978
rect 281994 418294 282050 418350
rect 282118 418294 282174 418350
rect 282242 418294 282298 418350
rect 282366 418294 282422 418350
rect 281994 418170 282050 418226
rect 282118 418170 282174 418226
rect 282242 418170 282298 418226
rect 282366 418170 282422 418226
rect 281994 418046 282050 418102
rect 282118 418046 282174 418102
rect 282242 418046 282298 418102
rect 282366 418046 282422 418102
rect 281994 417922 282050 417978
rect 282118 417922 282174 417978
rect 282242 417922 282298 417978
rect 282366 417922 282422 417978
rect 281994 400294 282050 400350
rect 282118 400294 282174 400350
rect 282242 400294 282298 400350
rect 282366 400294 282422 400350
rect 281994 400170 282050 400226
rect 282118 400170 282174 400226
rect 282242 400170 282298 400226
rect 282366 400170 282422 400226
rect 281994 400046 282050 400102
rect 282118 400046 282174 400102
rect 282242 400046 282298 400102
rect 282366 400046 282422 400102
rect 281994 399922 282050 399978
rect 282118 399922 282174 399978
rect 282242 399922 282298 399978
rect 282366 399922 282422 399978
rect 281994 382294 282050 382350
rect 282118 382294 282174 382350
rect 282242 382294 282298 382350
rect 282366 382294 282422 382350
rect 281994 382170 282050 382226
rect 282118 382170 282174 382226
rect 282242 382170 282298 382226
rect 282366 382170 282422 382226
rect 281994 382046 282050 382102
rect 282118 382046 282174 382102
rect 282242 382046 282298 382102
rect 282366 382046 282422 382102
rect 281994 381922 282050 381978
rect 282118 381922 282174 381978
rect 282242 381922 282298 381978
rect 282366 381922 282422 381978
rect 281994 364294 282050 364350
rect 282118 364294 282174 364350
rect 282242 364294 282298 364350
rect 282366 364294 282422 364350
rect 281994 364170 282050 364226
rect 282118 364170 282174 364226
rect 282242 364170 282298 364226
rect 282366 364170 282422 364226
rect 281994 364046 282050 364102
rect 282118 364046 282174 364102
rect 282242 364046 282298 364102
rect 282366 364046 282422 364102
rect 281994 363922 282050 363978
rect 282118 363922 282174 363978
rect 282242 363922 282298 363978
rect 282366 363922 282422 363978
rect 281994 346294 282050 346350
rect 282118 346294 282174 346350
rect 282242 346294 282298 346350
rect 282366 346294 282422 346350
rect 281994 346170 282050 346226
rect 282118 346170 282174 346226
rect 282242 346170 282298 346226
rect 282366 346170 282422 346226
rect 281994 346046 282050 346102
rect 282118 346046 282174 346102
rect 282242 346046 282298 346102
rect 282366 346046 282422 346102
rect 281994 345922 282050 345978
rect 282118 345922 282174 345978
rect 282242 345922 282298 345978
rect 282366 345922 282422 345978
rect 281994 328294 282050 328350
rect 282118 328294 282174 328350
rect 282242 328294 282298 328350
rect 282366 328294 282422 328350
rect 281994 328170 282050 328226
rect 282118 328170 282174 328226
rect 282242 328170 282298 328226
rect 282366 328170 282422 328226
rect 281994 328046 282050 328102
rect 282118 328046 282174 328102
rect 282242 328046 282298 328102
rect 282366 328046 282422 328102
rect 281994 327922 282050 327978
rect 282118 327922 282174 327978
rect 282242 327922 282298 327978
rect 282366 327922 282422 327978
rect 281994 310294 282050 310350
rect 282118 310294 282174 310350
rect 282242 310294 282298 310350
rect 282366 310294 282422 310350
rect 281994 310170 282050 310226
rect 282118 310170 282174 310226
rect 282242 310170 282298 310226
rect 282366 310170 282422 310226
rect 281994 310046 282050 310102
rect 282118 310046 282174 310102
rect 282242 310046 282298 310102
rect 282366 310046 282422 310102
rect 281994 309922 282050 309978
rect 282118 309922 282174 309978
rect 282242 309922 282298 309978
rect 282366 309922 282422 309978
rect 281994 292294 282050 292350
rect 282118 292294 282174 292350
rect 282242 292294 282298 292350
rect 282366 292294 282422 292350
rect 281994 292170 282050 292226
rect 282118 292170 282174 292226
rect 282242 292170 282298 292226
rect 282366 292170 282422 292226
rect 281994 292046 282050 292102
rect 282118 292046 282174 292102
rect 282242 292046 282298 292102
rect 282366 292046 282422 292102
rect 281994 291922 282050 291978
rect 282118 291922 282174 291978
rect 282242 291922 282298 291978
rect 282366 291922 282422 291978
rect 281994 274294 282050 274350
rect 282118 274294 282174 274350
rect 282242 274294 282298 274350
rect 282366 274294 282422 274350
rect 281994 274170 282050 274226
rect 282118 274170 282174 274226
rect 282242 274170 282298 274226
rect 282366 274170 282422 274226
rect 281994 274046 282050 274102
rect 282118 274046 282174 274102
rect 282242 274046 282298 274102
rect 282366 274046 282422 274102
rect 281994 273922 282050 273978
rect 282118 273922 282174 273978
rect 282242 273922 282298 273978
rect 282366 273922 282422 273978
rect 281994 256294 282050 256350
rect 282118 256294 282174 256350
rect 282242 256294 282298 256350
rect 282366 256294 282422 256350
rect 281994 256170 282050 256226
rect 282118 256170 282174 256226
rect 282242 256170 282298 256226
rect 282366 256170 282422 256226
rect 281994 256046 282050 256102
rect 282118 256046 282174 256102
rect 282242 256046 282298 256102
rect 282366 256046 282422 256102
rect 281994 255922 282050 255978
rect 282118 255922 282174 255978
rect 282242 255922 282298 255978
rect 282366 255922 282422 255978
rect 281994 238294 282050 238350
rect 282118 238294 282174 238350
rect 282242 238294 282298 238350
rect 282366 238294 282422 238350
rect 281994 238170 282050 238226
rect 282118 238170 282174 238226
rect 282242 238170 282298 238226
rect 282366 238170 282422 238226
rect 281994 238046 282050 238102
rect 282118 238046 282174 238102
rect 282242 238046 282298 238102
rect 282366 238046 282422 238102
rect 281994 237922 282050 237978
rect 282118 237922 282174 237978
rect 282242 237922 282298 237978
rect 282366 237922 282422 237978
rect 281994 220294 282050 220350
rect 282118 220294 282174 220350
rect 282242 220294 282298 220350
rect 282366 220294 282422 220350
rect 281994 220170 282050 220226
rect 282118 220170 282174 220226
rect 282242 220170 282298 220226
rect 282366 220170 282422 220226
rect 281994 220046 282050 220102
rect 282118 220046 282174 220102
rect 282242 220046 282298 220102
rect 282366 220046 282422 220102
rect 281994 219922 282050 219978
rect 282118 219922 282174 219978
rect 282242 219922 282298 219978
rect 282366 219922 282422 219978
rect 281994 202294 282050 202350
rect 282118 202294 282174 202350
rect 282242 202294 282298 202350
rect 282366 202294 282422 202350
rect 281994 202170 282050 202226
rect 282118 202170 282174 202226
rect 282242 202170 282298 202226
rect 282366 202170 282422 202226
rect 281994 202046 282050 202102
rect 282118 202046 282174 202102
rect 282242 202046 282298 202102
rect 282366 202046 282422 202102
rect 281994 201922 282050 201978
rect 282118 201922 282174 201978
rect 282242 201922 282298 201978
rect 282366 201922 282422 201978
rect 281994 184294 282050 184350
rect 282118 184294 282174 184350
rect 282242 184294 282298 184350
rect 282366 184294 282422 184350
rect 281994 184170 282050 184226
rect 282118 184170 282174 184226
rect 282242 184170 282298 184226
rect 282366 184170 282422 184226
rect 281994 184046 282050 184102
rect 282118 184046 282174 184102
rect 282242 184046 282298 184102
rect 282366 184046 282422 184102
rect 281994 183922 282050 183978
rect 282118 183922 282174 183978
rect 282242 183922 282298 183978
rect 282366 183922 282422 183978
rect 281994 166294 282050 166350
rect 282118 166294 282174 166350
rect 282242 166294 282298 166350
rect 282366 166294 282422 166350
rect 281994 166170 282050 166226
rect 282118 166170 282174 166226
rect 282242 166170 282298 166226
rect 282366 166170 282422 166226
rect 281994 166046 282050 166102
rect 282118 166046 282174 166102
rect 282242 166046 282298 166102
rect 282366 166046 282422 166102
rect 281994 165922 282050 165978
rect 282118 165922 282174 165978
rect 282242 165922 282298 165978
rect 282366 165922 282422 165978
rect 281994 148294 282050 148350
rect 282118 148294 282174 148350
rect 282242 148294 282298 148350
rect 282366 148294 282422 148350
rect 281994 148170 282050 148226
rect 282118 148170 282174 148226
rect 282242 148170 282298 148226
rect 282366 148170 282422 148226
rect 281994 148046 282050 148102
rect 282118 148046 282174 148102
rect 282242 148046 282298 148102
rect 282366 148046 282422 148102
rect 281994 147922 282050 147978
rect 282118 147922 282174 147978
rect 282242 147922 282298 147978
rect 282366 147922 282422 147978
rect 281994 130294 282050 130350
rect 282118 130294 282174 130350
rect 282242 130294 282298 130350
rect 282366 130294 282422 130350
rect 281994 130170 282050 130226
rect 282118 130170 282174 130226
rect 282242 130170 282298 130226
rect 282366 130170 282422 130226
rect 281994 130046 282050 130102
rect 282118 130046 282174 130102
rect 282242 130046 282298 130102
rect 282366 130046 282422 130102
rect 281994 129922 282050 129978
rect 282118 129922 282174 129978
rect 282242 129922 282298 129978
rect 282366 129922 282422 129978
rect 281994 112294 282050 112350
rect 282118 112294 282174 112350
rect 282242 112294 282298 112350
rect 282366 112294 282422 112350
rect 281994 112170 282050 112226
rect 282118 112170 282174 112226
rect 282242 112170 282298 112226
rect 282366 112170 282422 112226
rect 281994 112046 282050 112102
rect 282118 112046 282174 112102
rect 282242 112046 282298 112102
rect 282366 112046 282422 112102
rect 281994 111922 282050 111978
rect 282118 111922 282174 111978
rect 282242 111922 282298 111978
rect 282366 111922 282422 111978
rect 281994 94294 282050 94350
rect 282118 94294 282174 94350
rect 282242 94294 282298 94350
rect 282366 94294 282422 94350
rect 281994 94170 282050 94226
rect 282118 94170 282174 94226
rect 282242 94170 282298 94226
rect 282366 94170 282422 94226
rect 281994 94046 282050 94102
rect 282118 94046 282174 94102
rect 282242 94046 282298 94102
rect 282366 94046 282422 94102
rect 281994 93922 282050 93978
rect 282118 93922 282174 93978
rect 282242 93922 282298 93978
rect 282366 93922 282422 93978
rect 281994 76294 282050 76350
rect 282118 76294 282174 76350
rect 282242 76294 282298 76350
rect 282366 76294 282422 76350
rect 281994 76170 282050 76226
rect 282118 76170 282174 76226
rect 282242 76170 282298 76226
rect 282366 76170 282422 76226
rect 281994 76046 282050 76102
rect 282118 76046 282174 76102
rect 282242 76046 282298 76102
rect 282366 76046 282422 76102
rect 281994 75922 282050 75978
rect 282118 75922 282174 75978
rect 282242 75922 282298 75978
rect 282366 75922 282422 75978
rect 263788 70982 263844 71038
rect 254994 64294 255050 64350
rect 255118 64294 255174 64350
rect 255242 64294 255298 64350
rect 255366 64294 255422 64350
rect 254994 64170 255050 64226
rect 255118 64170 255174 64226
rect 255242 64170 255298 64226
rect 255366 64170 255422 64226
rect 254994 64046 255050 64102
rect 255118 64046 255174 64102
rect 255242 64046 255298 64102
rect 255366 64046 255422 64102
rect 254994 63922 255050 63978
rect 255118 63922 255174 63978
rect 255242 63922 255298 63978
rect 255366 63922 255422 63978
rect 254994 46294 255050 46350
rect 255118 46294 255174 46350
rect 255242 46294 255298 46350
rect 255366 46294 255422 46350
rect 254994 46170 255050 46226
rect 255118 46170 255174 46226
rect 255242 46170 255298 46226
rect 255366 46170 255422 46226
rect 254994 46046 255050 46102
rect 255118 46046 255174 46102
rect 255242 46046 255298 46102
rect 255366 46046 255422 46102
rect 254994 45922 255050 45978
rect 255118 45922 255174 45978
rect 255242 45922 255298 45978
rect 255366 45922 255422 45978
rect 254994 28294 255050 28350
rect 255118 28294 255174 28350
rect 255242 28294 255298 28350
rect 255366 28294 255422 28350
rect 254994 28170 255050 28226
rect 255118 28170 255174 28226
rect 255242 28170 255298 28226
rect 255366 28170 255422 28226
rect 254994 28046 255050 28102
rect 255118 28046 255174 28102
rect 255242 28046 255298 28102
rect 255366 28046 255422 28102
rect 254994 27922 255050 27978
rect 255118 27922 255174 27978
rect 255242 27922 255298 27978
rect 255366 27922 255422 27978
rect 258748 66122 258804 66178
rect 260428 42362 260484 42418
rect 254994 10294 255050 10350
rect 255118 10294 255174 10350
rect 255242 10294 255298 10350
rect 255366 10294 255422 10350
rect 254994 10170 255050 10226
rect 255118 10170 255174 10226
rect 255242 10170 255298 10226
rect 255366 10170 255422 10226
rect 254994 10046 255050 10102
rect 255118 10046 255174 10102
rect 255242 10046 255298 10102
rect 255366 10046 255422 10102
rect 254994 9922 255050 9978
rect 255118 9922 255174 9978
rect 255242 9922 255298 9978
rect 255366 9922 255422 9978
rect 251274 4046 251330 4102
rect 251398 4046 251454 4102
rect 251522 4046 251578 4102
rect 251646 4046 251702 4102
rect 251274 3922 251330 3978
rect 251398 3922 251454 3978
rect 251522 3922 251578 3978
rect 251646 3922 251702 3978
rect 251274 -216 251330 -160
rect 251398 -216 251454 -160
rect 251522 -216 251578 -160
rect 251646 -216 251702 -160
rect 251274 -340 251330 -284
rect 251398 -340 251454 -284
rect 251522 -340 251578 -284
rect 251646 -340 251702 -284
rect 251274 -464 251330 -408
rect 251398 -464 251454 -408
rect 251522 -464 251578 -408
rect 251646 -464 251702 -408
rect 251274 -588 251330 -532
rect 251398 -588 251454 -532
rect 251522 -588 251578 -532
rect 251646 -588 251702 -532
rect 257068 7082 257124 7138
rect 262108 15542 262164 15598
rect 273868 59642 273924 59698
rect 265468 56042 265524 56098
rect 281994 58294 282050 58350
rect 282118 58294 282174 58350
rect 282242 58294 282298 58350
rect 282366 58294 282422 58350
rect 281994 58170 282050 58226
rect 282118 58170 282174 58226
rect 282242 58170 282298 58226
rect 282366 58170 282422 58226
rect 281994 58046 282050 58102
rect 282118 58046 282174 58102
rect 282242 58046 282298 58102
rect 282366 58046 282422 58102
rect 281994 57922 282050 57978
rect 282118 57922 282174 57978
rect 282242 57922 282298 57978
rect 282366 57922 282422 57978
rect 285714 598116 285770 598172
rect 285838 598116 285894 598172
rect 285962 598116 286018 598172
rect 286086 598116 286142 598172
rect 285714 597992 285770 598048
rect 285838 597992 285894 598048
rect 285962 597992 286018 598048
rect 286086 597992 286142 598048
rect 285714 597868 285770 597924
rect 285838 597868 285894 597924
rect 285962 597868 286018 597924
rect 286086 597868 286142 597924
rect 285714 597744 285770 597800
rect 285838 597744 285894 597800
rect 285962 597744 286018 597800
rect 286086 597744 286142 597800
rect 312714 597156 312770 597212
rect 312838 597156 312894 597212
rect 312962 597156 313018 597212
rect 313086 597156 313142 597212
rect 312714 597032 312770 597088
rect 312838 597032 312894 597088
rect 312962 597032 313018 597088
rect 313086 597032 313142 597088
rect 312714 596908 312770 596964
rect 312838 596908 312894 596964
rect 312962 596908 313018 596964
rect 313086 596908 313142 596964
rect 312714 596784 312770 596840
rect 312838 596784 312894 596840
rect 312962 596784 313018 596840
rect 313086 596784 313142 596840
rect 285714 586294 285770 586350
rect 285838 586294 285894 586350
rect 285962 586294 286018 586350
rect 286086 586294 286142 586350
rect 285714 586170 285770 586226
rect 285838 586170 285894 586226
rect 285962 586170 286018 586226
rect 286086 586170 286142 586226
rect 285714 586046 285770 586102
rect 285838 586046 285894 586102
rect 285962 586046 286018 586102
rect 286086 586046 286142 586102
rect 285714 585922 285770 585978
rect 285838 585922 285894 585978
rect 285962 585922 286018 585978
rect 286086 585922 286142 585978
rect 285714 568294 285770 568350
rect 285838 568294 285894 568350
rect 285962 568294 286018 568350
rect 286086 568294 286142 568350
rect 285714 568170 285770 568226
rect 285838 568170 285894 568226
rect 285962 568170 286018 568226
rect 286086 568170 286142 568226
rect 285714 568046 285770 568102
rect 285838 568046 285894 568102
rect 285962 568046 286018 568102
rect 286086 568046 286142 568102
rect 285714 567922 285770 567978
rect 285838 567922 285894 567978
rect 285962 567922 286018 567978
rect 286086 567922 286142 567978
rect 285714 550294 285770 550350
rect 285838 550294 285894 550350
rect 285962 550294 286018 550350
rect 286086 550294 286142 550350
rect 285714 550170 285770 550226
rect 285838 550170 285894 550226
rect 285962 550170 286018 550226
rect 286086 550170 286142 550226
rect 285714 550046 285770 550102
rect 285838 550046 285894 550102
rect 285962 550046 286018 550102
rect 286086 550046 286142 550102
rect 285714 549922 285770 549978
rect 285838 549922 285894 549978
rect 285962 549922 286018 549978
rect 286086 549922 286142 549978
rect 285714 532294 285770 532350
rect 285838 532294 285894 532350
rect 285962 532294 286018 532350
rect 286086 532294 286142 532350
rect 285714 532170 285770 532226
rect 285838 532170 285894 532226
rect 285962 532170 286018 532226
rect 286086 532170 286142 532226
rect 285714 532046 285770 532102
rect 285838 532046 285894 532102
rect 285962 532046 286018 532102
rect 286086 532046 286142 532102
rect 285714 531922 285770 531978
rect 285838 531922 285894 531978
rect 285962 531922 286018 531978
rect 286086 531922 286142 531978
rect 285714 514294 285770 514350
rect 285838 514294 285894 514350
rect 285962 514294 286018 514350
rect 286086 514294 286142 514350
rect 285714 514170 285770 514226
rect 285838 514170 285894 514226
rect 285962 514170 286018 514226
rect 286086 514170 286142 514226
rect 285714 514046 285770 514102
rect 285838 514046 285894 514102
rect 285962 514046 286018 514102
rect 286086 514046 286142 514102
rect 285714 513922 285770 513978
rect 285838 513922 285894 513978
rect 285962 513922 286018 513978
rect 286086 513922 286142 513978
rect 285714 496294 285770 496350
rect 285838 496294 285894 496350
rect 285962 496294 286018 496350
rect 286086 496294 286142 496350
rect 285714 496170 285770 496226
rect 285838 496170 285894 496226
rect 285962 496170 286018 496226
rect 286086 496170 286142 496226
rect 285714 496046 285770 496102
rect 285838 496046 285894 496102
rect 285962 496046 286018 496102
rect 286086 496046 286142 496102
rect 285714 495922 285770 495978
rect 285838 495922 285894 495978
rect 285962 495922 286018 495978
rect 286086 495922 286142 495978
rect 285714 478294 285770 478350
rect 285838 478294 285894 478350
rect 285962 478294 286018 478350
rect 286086 478294 286142 478350
rect 285714 478170 285770 478226
rect 285838 478170 285894 478226
rect 285962 478170 286018 478226
rect 286086 478170 286142 478226
rect 285714 478046 285770 478102
rect 285838 478046 285894 478102
rect 285962 478046 286018 478102
rect 286086 478046 286142 478102
rect 285714 477922 285770 477978
rect 285838 477922 285894 477978
rect 285962 477922 286018 477978
rect 286086 477922 286142 477978
rect 285714 460294 285770 460350
rect 285838 460294 285894 460350
rect 285962 460294 286018 460350
rect 286086 460294 286142 460350
rect 285714 460170 285770 460226
rect 285838 460170 285894 460226
rect 285962 460170 286018 460226
rect 286086 460170 286142 460226
rect 285714 460046 285770 460102
rect 285838 460046 285894 460102
rect 285962 460046 286018 460102
rect 286086 460046 286142 460102
rect 285714 459922 285770 459978
rect 285838 459922 285894 459978
rect 285962 459922 286018 459978
rect 286086 459922 286142 459978
rect 285714 442294 285770 442350
rect 285838 442294 285894 442350
rect 285962 442294 286018 442350
rect 286086 442294 286142 442350
rect 285714 442170 285770 442226
rect 285838 442170 285894 442226
rect 285962 442170 286018 442226
rect 286086 442170 286142 442226
rect 285714 442046 285770 442102
rect 285838 442046 285894 442102
rect 285962 442046 286018 442102
rect 286086 442046 286142 442102
rect 285714 441922 285770 441978
rect 285838 441922 285894 441978
rect 285962 441922 286018 441978
rect 286086 441922 286142 441978
rect 285714 424294 285770 424350
rect 285838 424294 285894 424350
rect 285962 424294 286018 424350
rect 286086 424294 286142 424350
rect 285714 424170 285770 424226
rect 285838 424170 285894 424226
rect 285962 424170 286018 424226
rect 286086 424170 286142 424226
rect 285714 424046 285770 424102
rect 285838 424046 285894 424102
rect 285962 424046 286018 424102
rect 286086 424046 286142 424102
rect 285714 423922 285770 423978
rect 285838 423922 285894 423978
rect 285962 423922 286018 423978
rect 286086 423922 286142 423978
rect 285714 406294 285770 406350
rect 285838 406294 285894 406350
rect 285962 406294 286018 406350
rect 286086 406294 286142 406350
rect 285714 406170 285770 406226
rect 285838 406170 285894 406226
rect 285962 406170 286018 406226
rect 286086 406170 286142 406226
rect 285714 406046 285770 406102
rect 285838 406046 285894 406102
rect 285962 406046 286018 406102
rect 286086 406046 286142 406102
rect 285714 405922 285770 405978
rect 285838 405922 285894 405978
rect 285962 405922 286018 405978
rect 286086 405922 286142 405978
rect 285714 388294 285770 388350
rect 285838 388294 285894 388350
rect 285962 388294 286018 388350
rect 286086 388294 286142 388350
rect 285714 388170 285770 388226
rect 285838 388170 285894 388226
rect 285962 388170 286018 388226
rect 286086 388170 286142 388226
rect 285714 388046 285770 388102
rect 285838 388046 285894 388102
rect 285962 388046 286018 388102
rect 286086 388046 286142 388102
rect 285714 387922 285770 387978
rect 285838 387922 285894 387978
rect 285962 387922 286018 387978
rect 286086 387922 286142 387978
rect 285714 370294 285770 370350
rect 285838 370294 285894 370350
rect 285962 370294 286018 370350
rect 286086 370294 286142 370350
rect 285714 370170 285770 370226
rect 285838 370170 285894 370226
rect 285962 370170 286018 370226
rect 286086 370170 286142 370226
rect 285714 370046 285770 370102
rect 285838 370046 285894 370102
rect 285962 370046 286018 370102
rect 286086 370046 286142 370102
rect 285714 369922 285770 369978
rect 285838 369922 285894 369978
rect 285962 369922 286018 369978
rect 286086 369922 286142 369978
rect 285714 352294 285770 352350
rect 285838 352294 285894 352350
rect 285962 352294 286018 352350
rect 286086 352294 286142 352350
rect 285714 352170 285770 352226
rect 285838 352170 285894 352226
rect 285962 352170 286018 352226
rect 286086 352170 286142 352226
rect 285714 352046 285770 352102
rect 285838 352046 285894 352102
rect 285962 352046 286018 352102
rect 286086 352046 286142 352102
rect 285714 351922 285770 351978
rect 285838 351922 285894 351978
rect 285962 351922 286018 351978
rect 286086 351922 286142 351978
rect 285714 334294 285770 334350
rect 285838 334294 285894 334350
rect 285962 334294 286018 334350
rect 286086 334294 286142 334350
rect 285714 334170 285770 334226
rect 285838 334170 285894 334226
rect 285962 334170 286018 334226
rect 286086 334170 286142 334226
rect 285714 334046 285770 334102
rect 285838 334046 285894 334102
rect 285962 334046 286018 334102
rect 286086 334046 286142 334102
rect 285714 333922 285770 333978
rect 285838 333922 285894 333978
rect 285962 333922 286018 333978
rect 286086 333922 286142 333978
rect 285714 316294 285770 316350
rect 285838 316294 285894 316350
rect 285962 316294 286018 316350
rect 286086 316294 286142 316350
rect 285714 316170 285770 316226
rect 285838 316170 285894 316226
rect 285962 316170 286018 316226
rect 286086 316170 286142 316226
rect 285714 316046 285770 316102
rect 285838 316046 285894 316102
rect 285962 316046 286018 316102
rect 286086 316046 286142 316102
rect 285714 315922 285770 315978
rect 285838 315922 285894 315978
rect 285962 315922 286018 315978
rect 286086 315922 286142 315978
rect 285714 298294 285770 298350
rect 285838 298294 285894 298350
rect 285962 298294 286018 298350
rect 286086 298294 286142 298350
rect 285714 298170 285770 298226
rect 285838 298170 285894 298226
rect 285962 298170 286018 298226
rect 286086 298170 286142 298226
rect 285714 298046 285770 298102
rect 285838 298046 285894 298102
rect 285962 298046 286018 298102
rect 286086 298046 286142 298102
rect 285714 297922 285770 297978
rect 285838 297922 285894 297978
rect 285962 297922 286018 297978
rect 286086 297922 286142 297978
rect 285714 280294 285770 280350
rect 285838 280294 285894 280350
rect 285962 280294 286018 280350
rect 286086 280294 286142 280350
rect 285714 280170 285770 280226
rect 285838 280170 285894 280226
rect 285962 280170 286018 280226
rect 286086 280170 286142 280226
rect 285714 280046 285770 280102
rect 285838 280046 285894 280102
rect 285962 280046 286018 280102
rect 286086 280046 286142 280102
rect 285714 279922 285770 279978
rect 285838 279922 285894 279978
rect 285962 279922 286018 279978
rect 286086 279922 286142 279978
rect 285714 262294 285770 262350
rect 285838 262294 285894 262350
rect 285962 262294 286018 262350
rect 286086 262294 286142 262350
rect 285714 262170 285770 262226
rect 285838 262170 285894 262226
rect 285962 262170 286018 262226
rect 286086 262170 286142 262226
rect 285714 262046 285770 262102
rect 285838 262046 285894 262102
rect 285962 262046 286018 262102
rect 286086 262046 286142 262102
rect 285714 261922 285770 261978
rect 285838 261922 285894 261978
rect 285962 261922 286018 261978
rect 286086 261922 286142 261978
rect 285714 244294 285770 244350
rect 285838 244294 285894 244350
rect 285962 244294 286018 244350
rect 286086 244294 286142 244350
rect 285714 244170 285770 244226
rect 285838 244170 285894 244226
rect 285962 244170 286018 244226
rect 286086 244170 286142 244226
rect 285714 244046 285770 244102
rect 285838 244046 285894 244102
rect 285962 244046 286018 244102
rect 286086 244046 286142 244102
rect 285714 243922 285770 243978
rect 285838 243922 285894 243978
rect 285962 243922 286018 243978
rect 286086 243922 286142 243978
rect 285714 226294 285770 226350
rect 285838 226294 285894 226350
rect 285962 226294 286018 226350
rect 286086 226294 286142 226350
rect 285714 226170 285770 226226
rect 285838 226170 285894 226226
rect 285962 226170 286018 226226
rect 286086 226170 286142 226226
rect 285714 226046 285770 226102
rect 285838 226046 285894 226102
rect 285962 226046 286018 226102
rect 286086 226046 286142 226102
rect 285714 225922 285770 225978
rect 285838 225922 285894 225978
rect 285962 225922 286018 225978
rect 286086 225922 286142 225978
rect 285714 208294 285770 208350
rect 285838 208294 285894 208350
rect 285962 208294 286018 208350
rect 286086 208294 286142 208350
rect 285714 208170 285770 208226
rect 285838 208170 285894 208226
rect 285962 208170 286018 208226
rect 286086 208170 286142 208226
rect 285714 208046 285770 208102
rect 285838 208046 285894 208102
rect 285962 208046 286018 208102
rect 286086 208046 286142 208102
rect 285714 207922 285770 207978
rect 285838 207922 285894 207978
rect 285962 207922 286018 207978
rect 286086 207922 286142 207978
rect 285714 190294 285770 190350
rect 285838 190294 285894 190350
rect 285962 190294 286018 190350
rect 286086 190294 286142 190350
rect 285714 190170 285770 190226
rect 285838 190170 285894 190226
rect 285962 190170 286018 190226
rect 286086 190170 286142 190226
rect 285714 190046 285770 190102
rect 285838 190046 285894 190102
rect 285962 190046 286018 190102
rect 286086 190046 286142 190102
rect 285714 189922 285770 189978
rect 285838 189922 285894 189978
rect 285962 189922 286018 189978
rect 286086 189922 286142 189978
rect 285714 172294 285770 172350
rect 285838 172294 285894 172350
rect 285962 172294 286018 172350
rect 286086 172294 286142 172350
rect 285714 172170 285770 172226
rect 285838 172170 285894 172226
rect 285962 172170 286018 172226
rect 286086 172170 286142 172226
rect 285714 172046 285770 172102
rect 285838 172046 285894 172102
rect 285962 172046 286018 172102
rect 286086 172046 286142 172102
rect 285714 171922 285770 171978
rect 285838 171922 285894 171978
rect 285962 171922 286018 171978
rect 286086 171922 286142 171978
rect 285714 154294 285770 154350
rect 285838 154294 285894 154350
rect 285962 154294 286018 154350
rect 286086 154294 286142 154350
rect 285714 154170 285770 154226
rect 285838 154170 285894 154226
rect 285962 154170 286018 154226
rect 286086 154170 286142 154226
rect 285714 154046 285770 154102
rect 285838 154046 285894 154102
rect 285962 154046 286018 154102
rect 286086 154046 286142 154102
rect 285714 153922 285770 153978
rect 285838 153922 285894 153978
rect 285962 153922 286018 153978
rect 286086 153922 286142 153978
rect 285714 136294 285770 136350
rect 285838 136294 285894 136350
rect 285962 136294 286018 136350
rect 286086 136294 286142 136350
rect 285714 136170 285770 136226
rect 285838 136170 285894 136226
rect 285962 136170 286018 136226
rect 286086 136170 286142 136226
rect 285714 136046 285770 136102
rect 285838 136046 285894 136102
rect 285962 136046 286018 136102
rect 286086 136046 286142 136102
rect 285714 135922 285770 135978
rect 285838 135922 285894 135978
rect 285962 135922 286018 135978
rect 286086 135922 286142 135978
rect 285714 118294 285770 118350
rect 285838 118294 285894 118350
rect 285962 118294 286018 118350
rect 286086 118294 286142 118350
rect 285714 118170 285770 118226
rect 285838 118170 285894 118226
rect 285962 118170 286018 118226
rect 286086 118170 286142 118226
rect 285714 118046 285770 118102
rect 285838 118046 285894 118102
rect 285962 118046 286018 118102
rect 286086 118046 286142 118102
rect 285714 117922 285770 117978
rect 285838 117922 285894 117978
rect 285962 117922 286018 117978
rect 286086 117922 286142 117978
rect 285714 100294 285770 100350
rect 285838 100294 285894 100350
rect 285962 100294 286018 100350
rect 286086 100294 286142 100350
rect 285714 100170 285770 100226
rect 285838 100170 285894 100226
rect 285962 100170 286018 100226
rect 286086 100170 286142 100226
rect 285714 100046 285770 100102
rect 285838 100046 285894 100102
rect 285962 100046 286018 100102
rect 286086 100046 286142 100102
rect 285714 99922 285770 99978
rect 285838 99922 285894 99978
rect 285962 99922 286018 99978
rect 286086 99922 286142 99978
rect 285714 82294 285770 82350
rect 285838 82294 285894 82350
rect 285962 82294 286018 82350
rect 286086 82294 286142 82350
rect 285714 82170 285770 82226
rect 285838 82170 285894 82226
rect 285962 82170 286018 82226
rect 286086 82170 286142 82226
rect 285714 82046 285770 82102
rect 285838 82046 285894 82102
rect 285962 82046 286018 82102
rect 286086 82046 286142 82102
rect 285714 81922 285770 81978
rect 285838 81922 285894 81978
rect 285962 81922 286018 81978
rect 286086 81922 286142 81978
rect 297388 78182 297444 78238
rect 312714 580294 312770 580350
rect 312838 580294 312894 580350
rect 312962 580294 313018 580350
rect 313086 580294 313142 580350
rect 312714 580170 312770 580226
rect 312838 580170 312894 580226
rect 312962 580170 313018 580226
rect 313086 580170 313142 580226
rect 312714 580046 312770 580102
rect 312838 580046 312894 580102
rect 312962 580046 313018 580102
rect 313086 580046 313142 580102
rect 312714 579922 312770 579978
rect 312838 579922 312894 579978
rect 312962 579922 313018 579978
rect 313086 579922 313142 579978
rect 312714 562294 312770 562350
rect 312838 562294 312894 562350
rect 312962 562294 313018 562350
rect 313086 562294 313142 562350
rect 312714 562170 312770 562226
rect 312838 562170 312894 562226
rect 312962 562170 313018 562226
rect 313086 562170 313142 562226
rect 312714 562046 312770 562102
rect 312838 562046 312894 562102
rect 312962 562046 313018 562102
rect 313086 562046 313142 562102
rect 312714 561922 312770 561978
rect 312838 561922 312894 561978
rect 312962 561922 313018 561978
rect 313086 561922 313142 561978
rect 312714 544294 312770 544350
rect 312838 544294 312894 544350
rect 312962 544294 313018 544350
rect 313086 544294 313142 544350
rect 312714 544170 312770 544226
rect 312838 544170 312894 544226
rect 312962 544170 313018 544226
rect 313086 544170 313142 544226
rect 312714 544046 312770 544102
rect 312838 544046 312894 544102
rect 312962 544046 313018 544102
rect 313086 544046 313142 544102
rect 312714 543922 312770 543978
rect 312838 543922 312894 543978
rect 312962 543922 313018 543978
rect 313086 543922 313142 543978
rect 312714 526294 312770 526350
rect 312838 526294 312894 526350
rect 312962 526294 313018 526350
rect 313086 526294 313142 526350
rect 312714 526170 312770 526226
rect 312838 526170 312894 526226
rect 312962 526170 313018 526226
rect 313086 526170 313142 526226
rect 312714 526046 312770 526102
rect 312838 526046 312894 526102
rect 312962 526046 313018 526102
rect 313086 526046 313142 526102
rect 312714 525922 312770 525978
rect 312838 525922 312894 525978
rect 312962 525922 313018 525978
rect 313086 525922 313142 525978
rect 312714 508294 312770 508350
rect 312838 508294 312894 508350
rect 312962 508294 313018 508350
rect 313086 508294 313142 508350
rect 312714 508170 312770 508226
rect 312838 508170 312894 508226
rect 312962 508170 313018 508226
rect 313086 508170 313142 508226
rect 312714 508046 312770 508102
rect 312838 508046 312894 508102
rect 312962 508046 313018 508102
rect 313086 508046 313142 508102
rect 312714 507922 312770 507978
rect 312838 507922 312894 507978
rect 312962 507922 313018 507978
rect 313086 507922 313142 507978
rect 312714 490294 312770 490350
rect 312838 490294 312894 490350
rect 312962 490294 313018 490350
rect 313086 490294 313142 490350
rect 312714 490170 312770 490226
rect 312838 490170 312894 490226
rect 312962 490170 313018 490226
rect 313086 490170 313142 490226
rect 312714 490046 312770 490102
rect 312838 490046 312894 490102
rect 312962 490046 313018 490102
rect 313086 490046 313142 490102
rect 312714 489922 312770 489978
rect 312838 489922 312894 489978
rect 312962 489922 313018 489978
rect 313086 489922 313142 489978
rect 312714 472294 312770 472350
rect 312838 472294 312894 472350
rect 312962 472294 313018 472350
rect 313086 472294 313142 472350
rect 312714 472170 312770 472226
rect 312838 472170 312894 472226
rect 312962 472170 313018 472226
rect 313086 472170 313142 472226
rect 312714 472046 312770 472102
rect 312838 472046 312894 472102
rect 312962 472046 313018 472102
rect 313086 472046 313142 472102
rect 312714 471922 312770 471978
rect 312838 471922 312894 471978
rect 312962 471922 313018 471978
rect 313086 471922 313142 471978
rect 312714 454294 312770 454350
rect 312838 454294 312894 454350
rect 312962 454294 313018 454350
rect 313086 454294 313142 454350
rect 312714 454170 312770 454226
rect 312838 454170 312894 454226
rect 312962 454170 313018 454226
rect 313086 454170 313142 454226
rect 312714 454046 312770 454102
rect 312838 454046 312894 454102
rect 312962 454046 313018 454102
rect 313086 454046 313142 454102
rect 312714 453922 312770 453978
rect 312838 453922 312894 453978
rect 312962 453922 313018 453978
rect 313086 453922 313142 453978
rect 312714 436294 312770 436350
rect 312838 436294 312894 436350
rect 312962 436294 313018 436350
rect 313086 436294 313142 436350
rect 312714 436170 312770 436226
rect 312838 436170 312894 436226
rect 312962 436170 313018 436226
rect 313086 436170 313142 436226
rect 312714 436046 312770 436102
rect 312838 436046 312894 436102
rect 312962 436046 313018 436102
rect 313086 436046 313142 436102
rect 312714 435922 312770 435978
rect 312838 435922 312894 435978
rect 312962 435922 313018 435978
rect 313086 435922 313142 435978
rect 312714 418294 312770 418350
rect 312838 418294 312894 418350
rect 312962 418294 313018 418350
rect 313086 418294 313142 418350
rect 312714 418170 312770 418226
rect 312838 418170 312894 418226
rect 312962 418170 313018 418226
rect 313086 418170 313142 418226
rect 312714 418046 312770 418102
rect 312838 418046 312894 418102
rect 312962 418046 313018 418102
rect 313086 418046 313142 418102
rect 312714 417922 312770 417978
rect 312838 417922 312894 417978
rect 312962 417922 313018 417978
rect 313086 417922 313142 417978
rect 312714 400294 312770 400350
rect 312838 400294 312894 400350
rect 312962 400294 313018 400350
rect 313086 400294 313142 400350
rect 312714 400170 312770 400226
rect 312838 400170 312894 400226
rect 312962 400170 313018 400226
rect 313086 400170 313142 400226
rect 312714 400046 312770 400102
rect 312838 400046 312894 400102
rect 312962 400046 313018 400102
rect 313086 400046 313142 400102
rect 312714 399922 312770 399978
rect 312838 399922 312894 399978
rect 312962 399922 313018 399978
rect 313086 399922 313142 399978
rect 312714 382294 312770 382350
rect 312838 382294 312894 382350
rect 312962 382294 313018 382350
rect 313086 382294 313142 382350
rect 312714 382170 312770 382226
rect 312838 382170 312894 382226
rect 312962 382170 313018 382226
rect 313086 382170 313142 382226
rect 312714 382046 312770 382102
rect 312838 382046 312894 382102
rect 312962 382046 313018 382102
rect 313086 382046 313142 382102
rect 312714 381922 312770 381978
rect 312838 381922 312894 381978
rect 312962 381922 313018 381978
rect 313086 381922 313142 381978
rect 312714 364294 312770 364350
rect 312838 364294 312894 364350
rect 312962 364294 313018 364350
rect 313086 364294 313142 364350
rect 312714 364170 312770 364226
rect 312838 364170 312894 364226
rect 312962 364170 313018 364226
rect 313086 364170 313142 364226
rect 312714 364046 312770 364102
rect 312838 364046 312894 364102
rect 312962 364046 313018 364102
rect 313086 364046 313142 364102
rect 312714 363922 312770 363978
rect 312838 363922 312894 363978
rect 312962 363922 313018 363978
rect 313086 363922 313142 363978
rect 312714 346294 312770 346350
rect 312838 346294 312894 346350
rect 312962 346294 313018 346350
rect 313086 346294 313142 346350
rect 312714 346170 312770 346226
rect 312838 346170 312894 346226
rect 312962 346170 313018 346226
rect 313086 346170 313142 346226
rect 312714 346046 312770 346102
rect 312838 346046 312894 346102
rect 312962 346046 313018 346102
rect 313086 346046 313142 346102
rect 312714 345922 312770 345978
rect 312838 345922 312894 345978
rect 312962 345922 313018 345978
rect 313086 345922 313142 345978
rect 312714 328294 312770 328350
rect 312838 328294 312894 328350
rect 312962 328294 313018 328350
rect 313086 328294 313142 328350
rect 312714 328170 312770 328226
rect 312838 328170 312894 328226
rect 312962 328170 313018 328226
rect 313086 328170 313142 328226
rect 312714 328046 312770 328102
rect 312838 328046 312894 328102
rect 312962 328046 313018 328102
rect 313086 328046 313142 328102
rect 312714 327922 312770 327978
rect 312838 327922 312894 327978
rect 312962 327922 313018 327978
rect 313086 327922 313142 327978
rect 312714 310294 312770 310350
rect 312838 310294 312894 310350
rect 312962 310294 313018 310350
rect 313086 310294 313142 310350
rect 312714 310170 312770 310226
rect 312838 310170 312894 310226
rect 312962 310170 313018 310226
rect 313086 310170 313142 310226
rect 312714 310046 312770 310102
rect 312838 310046 312894 310102
rect 312962 310046 313018 310102
rect 313086 310046 313142 310102
rect 312714 309922 312770 309978
rect 312838 309922 312894 309978
rect 312962 309922 313018 309978
rect 313086 309922 313142 309978
rect 312714 292294 312770 292350
rect 312838 292294 312894 292350
rect 312962 292294 313018 292350
rect 313086 292294 313142 292350
rect 312714 292170 312770 292226
rect 312838 292170 312894 292226
rect 312962 292170 313018 292226
rect 313086 292170 313142 292226
rect 312714 292046 312770 292102
rect 312838 292046 312894 292102
rect 312962 292046 313018 292102
rect 313086 292046 313142 292102
rect 312714 291922 312770 291978
rect 312838 291922 312894 291978
rect 312962 291922 313018 291978
rect 313086 291922 313142 291978
rect 312714 274294 312770 274350
rect 312838 274294 312894 274350
rect 312962 274294 313018 274350
rect 313086 274294 313142 274350
rect 312714 274170 312770 274226
rect 312838 274170 312894 274226
rect 312962 274170 313018 274226
rect 313086 274170 313142 274226
rect 312714 274046 312770 274102
rect 312838 274046 312894 274102
rect 312962 274046 313018 274102
rect 313086 274046 313142 274102
rect 312714 273922 312770 273978
rect 312838 273922 312894 273978
rect 312962 273922 313018 273978
rect 313086 273922 313142 273978
rect 312714 256294 312770 256350
rect 312838 256294 312894 256350
rect 312962 256294 313018 256350
rect 313086 256294 313142 256350
rect 312714 256170 312770 256226
rect 312838 256170 312894 256226
rect 312962 256170 313018 256226
rect 313086 256170 313142 256226
rect 312714 256046 312770 256102
rect 312838 256046 312894 256102
rect 312962 256046 313018 256102
rect 313086 256046 313142 256102
rect 312714 255922 312770 255978
rect 312838 255922 312894 255978
rect 312962 255922 313018 255978
rect 313086 255922 313142 255978
rect 312714 238294 312770 238350
rect 312838 238294 312894 238350
rect 312962 238294 313018 238350
rect 313086 238294 313142 238350
rect 312714 238170 312770 238226
rect 312838 238170 312894 238226
rect 312962 238170 313018 238226
rect 313086 238170 313142 238226
rect 312714 238046 312770 238102
rect 312838 238046 312894 238102
rect 312962 238046 313018 238102
rect 313086 238046 313142 238102
rect 312714 237922 312770 237978
rect 312838 237922 312894 237978
rect 312962 237922 313018 237978
rect 313086 237922 313142 237978
rect 312714 220294 312770 220350
rect 312838 220294 312894 220350
rect 312962 220294 313018 220350
rect 313086 220294 313142 220350
rect 312714 220170 312770 220226
rect 312838 220170 312894 220226
rect 312962 220170 313018 220226
rect 313086 220170 313142 220226
rect 312714 220046 312770 220102
rect 312838 220046 312894 220102
rect 312962 220046 313018 220102
rect 313086 220046 313142 220102
rect 312714 219922 312770 219978
rect 312838 219922 312894 219978
rect 312962 219922 313018 219978
rect 313086 219922 313142 219978
rect 312714 202294 312770 202350
rect 312838 202294 312894 202350
rect 312962 202294 313018 202350
rect 313086 202294 313142 202350
rect 312714 202170 312770 202226
rect 312838 202170 312894 202226
rect 312962 202170 313018 202226
rect 313086 202170 313142 202226
rect 312714 202046 312770 202102
rect 312838 202046 312894 202102
rect 312962 202046 313018 202102
rect 313086 202046 313142 202102
rect 312714 201922 312770 201978
rect 312838 201922 312894 201978
rect 312962 201922 313018 201978
rect 313086 201922 313142 201978
rect 312714 184294 312770 184350
rect 312838 184294 312894 184350
rect 312962 184294 313018 184350
rect 313086 184294 313142 184350
rect 312714 184170 312770 184226
rect 312838 184170 312894 184226
rect 312962 184170 313018 184226
rect 313086 184170 313142 184226
rect 312714 184046 312770 184102
rect 312838 184046 312894 184102
rect 312962 184046 313018 184102
rect 313086 184046 313142 184102
rect 312714 183922 312770 183978
rect 312838 183922 312894 183978
rect 312962 183922 313018 183978
rect 313086 183922 313142 183978
rect 312714 166294 312770 166350
rect 312838 166294 312894 166350
rect 312962 166294 313018 166350
rect 313086 166294 313142 166350
rect 312714 166170 312770 166226
rect 312838 166170 312894 166226
rect 312962 166170 313018 166226
rect 313086 166170 313142 166226
rect 312714 166046 312770 166102
rect 312838 166046 312894 166102
rect 312962 166046 313018 166102
rect 313086 166046 313142 166102
rect 312714 165922 312770 165978
rect 312838 165922 312894 165978
rect 312962 165922 313018 165978
rect 313086 165922 313142 165978
rect 312714 148294 312770 148350
rect 312838 148294 312894 148350
rect 312962 148294 313018 148350
rect 313086 148294 313142 148350
rect 312714 148170 312770 148226
rect 312838 148170 312894 148226
rect 312962 148170 313018 148226
rect 313086 148170 313142 148226
rect 312714 148046 312770 148102
rect 312838 148046 312894 148102
rect 312962 148046 313018 148102
rect 313086 148046 313142 148102
rect 312714 147922 312770 147978
rect 312838 147922 312894 147978
rect 312962 147922 313018 147978
rect 313086 147922 313142 147978
rect 312714 130294 312770 130350
rect 312838 130294 312894 130350
rect 312962 130294 313018 130350
rect 313086 130294 313142 130350
rect 312714 130170 312770 130226
rect 312838 130170 312894 130226
rect 312962 130170 313018 130226
rect 313086 130170 313142 130226
rect 312714 130046 312770 130102
rect 312838 130046 312894 130102
rect 312962 130046 313018 130102
rect 313086 130046 313142 130102
rect 312714 129922 312770 129978
rect 312838 129922 312894 129978
rect 312962 129922 313018 129978
rect 313086 129922 313142 129978
rect 312714 112294 312770 112350
rect 312838 112294 312894 112350
rect 312962 112294 313018 112350
rect 313086 112294 313142 112350
rect 312714 112170 312770 112226
rect 312838 112170 312894 112226
rect 312962 112170 313018 112226
rect 313086 112170 313142 112226
rect 312714 112046 312770 112102
rect 312838 112046 312894 112102
rect 312962 112046 313018 112102
rect 313086 112046 313142 112102
rect 312714 111922 312770 111978
rect 312838 111922 312894 111978
rect 312962 111922 313018 111978
rect 313086 111922 313142 111978
rect 312714 94294 312770 94350
rect 312838 94294 312894 94350
rect 312962 94294 313018 94350
rect 313086 94294 313142 94350
rect 312714 94170 312770 94226
rect 312838 94170 312894 94226
rect 312962 94170 313018 94226
rect 313086 94170 313142 94226
rect 312714 94046 312770 94102
rect 312838 94046 312894 94102
rect 312962 94046 313018 94102
rect 313086 94046 313142 94102
rect 312714 93922 312770 93978
rect 312838 93922 312894 93978
rect 312962 93922 313018 93978
rect 313086 93922 313142 93978
rect 312714 76294 312770 76350
rect 312838 76294 312894 76350
rect 312962 76294 313018 76350
rect 313086 76294 313142 76350
rect 312714 76170 312770 76226
rect 312838 76170 312894 76226
rect 312962 76170 313018 76226
rect 313086 76170 313142 76226
rect 312714 76046 312770 76102
rect 312838 76046 312894 76102
rect 312962 76046 313018 76102
rect 313086 76046 313142 76102
rect 312714 75922 312770 75978
rect 312838 75922 312894 75978
rect 312962 75922 313018 75978
rect 313086 75922 313142 75978
rect 288988 70802 289044 70858
rect 285714 64294 285770 64350
rect 285838 64294 285894 64350
rect 285962 64294 286018 64350
rect 286086 64294 286142 64350
rect 285714 64170 285770 64226
rect 285838 64170 285894 64226
rect 285962 64170 286018 64226
rect 286086 64170 286142 64226
rect 285714 64046 285770 64102
rect 285838 64046 285894 64102
rect 285962 64046 286018 64102
rect 286086 64046 286142 64102
rect 285714 63922 285770 63978
rect 285838 63922 285894 63978
rect 285962 63922 286018 63978
rect 286086 63922 286142 63978
rect 281994 40294 282050 40350
rect 282118 40294 282174 40350
rect 282242 40294 282298 40350
rect 282366 40294 282422 40350
rect 281994 40170 282050 40226
rect 282118 40170 282174 40226
rect 282242 40170 282298 40226
rect 282366 40170 282422 40226
rect 281994 40046 282050 40102
rect 282118 40046 282174 40102
rect 282242 40046 282298 40102
rect 282366 40046 282422 40102
rect 281994 39922 282050 39978
rect 282118 39922 282174 39978
rect 282242 39922 282298 39978
rect 282366 39922 282422 39978
rect 278908 34262 278964 34318
rect 268380 5642 268436 5698
rect 281994 22294 282050 22350
rect 282118 22294 282174 22350
rect 282242 22294 282298 22350
rect 282366 22294 282422 22350
rect 281994 22170 282050 22226
rect 282118 22170 282174 22226
rect 282242 22170 282298 22226
rect 282366 22170 282422 22226
rect 281994 22046 282050 22102
rect 282118 22046 282174 22102
rect 282242 22046 282298 22102
rect 282366 22046 282422 22102
rect 281994 21922 282050 21978
rect 282118 21922 282174 21978
rect 282242 21922 282298 21978
rect 282366 21922 282422 21978
rect 281994 4294 282050 4350
rect 282118 4294 282174 4350
rect 282242 4294 282298 4350
rect 282366 4294 282422 4350
rect 281994 4170 282050 4226
rect 282118 4170 282174 4226
rect 282242 4170 282298 4226
rect 282366 4170 282422 4226
rect 282604 49562 282660 49618
rect 285714 46294 285770 46350
rect 285838 46294 285894 46350
rect 285962 46294 286018 46350
rect 286086 46294 286142 46350
rect 285714 46170 285770 46226
rect 285838 46170 285894 46226
rect 285962 46170 286018 46226
rect 286086 46170 286142 46226
rect 285714 46046 285770 46102
rect 285838 46046 285894 46102
rect 285962 46046 286018 46102
rect 286086 46046 286142 46102
rect 285714 45922 285770 45978
rect 285838 45922 285894 45978
rect 285962 45922 286018 45978
rect 286086 45922 286142 45978
rect 285714 28294 285770 28350
rect 285838 28294 285894 28350
rect 285962 28294 286018 28350
rect 286086 28294 286142 28350
rect 285714 28170 285770 28226
rect 285838 28170 285894 28226
rect 285962 28170 286018 28226
rect 286086 28170 286142 28226
rect 285714 28046 285770 28102
rect 285838 28046 285894 28102
rect 285962 28046 286018 28102
rect 286086 28046 286142 28102
rect 285714 27922 285770 27978
rect 285838 27922 285894 27978
rect 285962 27922 286018 27978
rect 286086 27922 286142 27978
rect 285714 10294 285770 10350
rect 285838 10294 285894 10350
rect 285962 10294 286018 10350
rect 286086 10294 286142 10350
rect 285714 10170 285770 10226
rect 285838 10170 285894 10226
rect 285962 10170 286018 10226
rect 286086 10170 286142 10226
rect 285714 10046 285770 10102
rect 285838 10046 285894 10102
rect 285962 10046 286018 10102
rect 286086 10046 286142 10102
rect 285714 9922 285770 9978
rect 285838 9922 285894 9978
rect 285962 9922 286018 9978
rect 286086 9922 286142 9978
rect 281994 4046 282050 4102
rect 282118 4046 282174 4102
rect 282242 4046 282298 4102
rect 282366 4046 282422 4102
rect 281994 3922 282050 3978
rect 282118 3922 282174 3978
rect 282242 3922 282298 3978
rect 282366 3922 282422 3978
rect 254994 -1176 255050 -1120
rect 255118 -1176 255174 -1120
rect 255242 -1176 255298 -1120
rect 255366 -1176 255422 -1120
rect 254994 -1300 255050 -1244
rect 255118 -1300 255174 -1244
rect 255242 -1300 255298 -1244
rect 255366 -1300 255422 -1244
rect 254994 -1424 255050 -1368
rect 255118 -1424 255174 -1368
rect 255242 -1424 255298 -1368
rect 255366 -1424 255422 -1368
rect 254994 -1548 255050 -1492
rect 255118 -1548 255174 -1492
rect 255242 -1548 255298 -1492
rect 255366 -1548 255422 -1492
rect 281994 -216 282050 -160
rect 282118 -216 282174 -160
rect 282242 -216 282298 -160
rect 282366 -216 282422 -160
rect 281994 -340 282050 -284
rect 282118 -340 282174 -284
rect 282242 -340 282298 -284
rect 282366 -340 282422 -284
rect 281994 -464 282050 -408
rect 282118 -464 282174 -408
rect 282242 -464 282298 -408
rect 282366 -464 282422 -408
rect 281994 -588 282050 -532
rect 282118 -588 282174 -532
rect 282242 -588 282298 -532
rect 282366 -588 282422 -532
rect 286300 69182 286356 69238
rect 295708 70622 295764 70678
rect 294028 67562 294084 67618
rect 290668 52622 290724 52678
rect 302428 69002 302484 69058
rect 300748 32102 300804 32158
rect 305788 67742 305844 67798
rect 312714 58294 312770 58350
rect 312838 58294 312894 58350
rect 312962 58294 313018 58350
rect 313086 58294 313142 58350
rect 312714 58170 312770 58226
rect 312838 58170 312894 58226
rect 312962 58170 313018 58226
rect 313086 58170 313142 58226
rect 312714 58046 312770 58102
rect 312838 58046 312894 58102
rect 312962 58046 313018 58102
rect 313086 58046 313142 58102
rect 312714 57922 312770 57978
rect 312838 57922 312894 57978
rect 312962 57922 313018 57978
rect 313086 57922 313142 57978
rect 312714 40294 312770 40350
rect 312838 40294 312894 40350
rect 312962 40294 313018 40350
rect 313086 40294 313142 40350
rect 312714 40170 312770 40226
rect 312838 40170 312894 40226
rect 312962 40170 313018 40226
rect 313086 40170 313142 40226
rect 312714 40046 312770 40102
rect 312838 40046 312894 40102
rect 312962 40046 313018 40102
rect 313086 40046 313142 40102
rect 312714 39922 312770 39978
rect 312838 39922 312894 39978
rect 312962 39922 313018 39978
rect 313086 39922 313142 39978
rect 310828 35702 310884 35758
rect 308364 5462 308420 5518
rect 316434 598116 316490 598172
rect 316558 598116 316614 598172
rect 316682 598116 316738 598172
rect 316806 598116 316862 598172
rect 316434 597992 316490 598048
rect 316558 597992 316614 598048
rect 316682 597992 316738 598048
rect 316806 597992 316862 598048
rect 316434 597868 316490 597924
rect 316558 597868 316614 597924
rect 316682 597868 316738 597924
rect 316806 597868 316862 597924
rect 316434 597744 316490 597800
rect 316558 597744 316614 597800
rect 316682 597744 316738 597800
rect 316806 597744 316862 597800
rect 343434 597156 343490 597212
rect 343558 597156 343614 597212
rect 343682 597156 343738 597212
rect 343806 597156 343862 597212
rect 343434 597032 343490 597088
rect 343558 597032 343614 597088
rect 343682 597032 343738 597088
rect 343806 597032 343862 597088
rect 343434 596908 343490 596964
rect 343558 596908 343614 596964
rect 343682 596908 343738 596964
rect 343806 596908 343862 596964
rect 343434 596784 343490 596840
rect 343558 596784 343614 596840
rect 343682 596784 343738 596840
rect 343806 596784 343862 596840
rect 316434 586294 316490 586350
rect 316558 586294 316614 586350
rect 316682 586294 316738 586350
rect 316806 586294 316862 586350
rect 316434 586170 316490 586226
rect 316558 586170 316614 586226
rect 316682 586170 316738 586226
rect 316806 586170 316862 586226
rect 316434 586046 316490 586102
rect 316558 586046 316614 586102
rect 316682 586046 316738 586102
rect 316806 586046 316862 586102
rect 316434 585922 316490 585978
rect 316558 585922 316614 585978
rect 316682 585922 316738 585978
rect 316806 585922 316862 585978
rect 316434 568294 316490 568350
rect 316558 568294 316614 568350
rect 316682 568294 316738 568350
rect 316806 568294 316862 568350
rect 316434 568170 316490 568226
rect 316558 568170 316614 568226
rect 316682 568170 316738 568226
rect 316806 568170 316862 568226
rect 316434 568046 316490 568102
rect 316558 568046 316614 568102
rect 316682 568046 316738 568102
rect 316806 568046 316862 568102
rect 316434 567922 316490 567978
rect 316558 567922 316614 567978
rect 316682 567922 316738 567978
rect 316806 567922 316862 567978
rect 316434 550294 316490 550350
rect 316558 550294 316614 550350
rect 316682 550294 316738 550350
rect 316806 550294 316862 550350
rect 316434 550170 316490 550226
rect 316558 550170 316614 550226
rect 316682 550170 316738 550226
rect 316806 550170 316862 550226
rect 316434 550046 316490 550102
rect 316558 550046 316614 550102
rect 316682 550046 316738 550102
rect 316806 550046 316862 550102
rect 316434 549922 316490 549978
rect 316558 549922 316614 549978
rect 316682 549922 316738 549978
rect 316806 549922 316862 549978
rect 316434 532294 316490 532350
rect 316558 532294 316614 532350
rect 316682 532294 316738 532350
rect 316806 532294 316862 532350
rect 316434 532170 316490 532226
rect 316558 532170 316614 532226
rect 316682 532170 316738 532226
rect 316806 532170 316862 532226
rect 316434 532046 316490 532102
rect 316558 532046 316614 532102
rect 316682 532046 316738 532102
rect 316806 532046 316862 532102
rect 316434 531922 316490 531978
rect 316558 531922 316614 531978
rect 316682 531922 316738 531978
rect 316806 531922 316862 531978
rect 316434 514294 316490 514350
rect 316558 514294 316614 514350
rect 316682 514294 316738 514350
rect 316806 514294 316862 514350
rect 316434 514170 316490 514226
rect 316558 514170 316614 514226
rect 316682 514170 316738 514226
rect 316806 514170 316862 514226
rect 316434 514046 316490 514102
rect 316558 514046 316614 514102
rect 316682 514046 316738 514102
rect 316806 514046 316862 514102
rect 316434 513922 316490 513978
rect 316558 513922 316614 513978
rect 316682 513922 316738 513978
rect 316806 513922 316862 513978
rect 316434 496294 316490 496350
rect 316558 496294 316614 496350
rect 316682 496294 316738 496350
rect 316806 496294 316862 496350
rect 316434 496170 316490 496226
rect 316558 496170 316614 496226
rect 316682 496170 316738 496226
rect 316806 496170 316862 496226
rect 316434 496046 316490 496102
rect 316558 496046 316614 496102
rect 316682 496046 316738 496102
rect 316806 496046 316862 496102
rect 316434 495922 316490 495978
rect 316558 495922 316614 495978
rect 316682 495922 316738 495978
rect 316806 495922 316862 495978
rect 316434 478294 316490 478350
rect 316558 478294 316614 478350
rect 316682 478294 316738 478350
rect 316806 478294 316862 478350
rect 316434 478170 316490 478226
rect 316558 478170 316614 478226
rect 316682 478170 316738 478226
rect 316806 478170 316862 478226
rect 316434 478046 316490 478102
rect 316558 478046 316614 478102
rect 316682 478046 316738 478102
rect 316806 478046 316862 478102
rect 316434 477922 316490 477978
rect 316558 477922 316614 477978
rect 316682 477922 316738 477978
rect 316806 477922 316862 477978
rect 316434 460294 316490 460350
rect 316558 460294 316614 460350
rect 316682 460294 316738 460350
rect 316806 460294 316862 460350
rect 316434 460170 316490 460226
rect 316558 460170 316614 460226
rect 316682 460170 316738 460226
rect 316806 460170 316862 460226
rect 316434 460046 316490 460102
rect 316558 460046 316614 460102
rect 316682 460046 316738 460102
rect 316806 460046 316862 460102
rect 316434 459922 316490 459978
rect 316558 459922 316614 459978
rect 316682 459922 316738 459978
rect 316806 459922 316862 459978
rect 316434 442294 316490 442350
rect 316558 442294 316614 442350
rect 316682 442294 316738 442350
rect 316806 442294 316862 442350
rect 316434 442170 316490 442226
rect 316558 442170 316614 442226
rect 316682 442170 316738 442226
rect 316806 442170 316862 442226
rect 316434 442046 316490 442102
rect 316558 442046 316614 442102
rect 316682 442046 316738 442102
rect 316806 442046 316862 442102
rect 316434 441922 316490 441978
rect 316558 441922 316614 441978
rect 316682 441922 316738 441978
rect 316806 441922 316862 441978
rect 316434 424294 316490 424350
rect 316558 424294 316614 424350
rect 316682 424294 316738 424350
rect 316806 424294 316862 424350
rect 316434 424170 316490 424226
rect 316558 424170 316614 424226
rect 316682 424170 316738 424226
rect 316806 424170 316862 424226
rect 316434 424046 316490 424102
rect 316558 424046 316614 424102
rect 316682 424046 316738 424102
rect 316806 424046 316862 424102
rect 316434 423922 316490 423978
rect 316558 423922 316614 423978
rect 316682 423922 316738 423978
rect 316806 423922 316862 423978
rect 316434 406294 316490 406350
rect 316558 406294 316614 406350
rect 316682 406294 316738 406350
rect 316806 406294 316862 406350
rect 316434 406170 316490 406226
rect 316558 406170 316614 406226
rect 316682 406170 316738 406226
rect 316806 406170 316862 406226
rect 316434 406046 316490 406102
rect 316558 406046 316614 406102
rect 316682 406046 316738 406102
rect 316806 406046 316862 406102
rect 316434 405922 316490 405978
rect 316558 405922 316614 405978
rect 316682 405922 316738 405978
rect 316806 405922 316862 405978
rect 316434 388294 316490 388350
rect 316558 388294 316614 388350
rect 316682 388294 316738 388350
rect 316806 388294 316862 388350
rect 316434 388170 316490 388226
rect 316558 388170 316614 388226
rect 316682 388170 316738 388226
rect 316806 388170 316862 388226
rect 316434 388046 316490 388102
rect 316558 388046 316614 388102
rect 316682 388046 316738 388102
rect 316806 388046 316862 388102
rect 316434 387922 316490 387978
rect 316558 387922 316614 387978
rect 316682 387922 316738 387978
rect 316806 387922 316862 387978
rect 316434 370294 316490 370350
rect 316558 370294 316614 370350
rect 316682 370294 316738 370350
rect 316806 370294 316862 370350
rect 316434 370170 316490 370226
rect 316558 370170 316614 370226
rect 316682 370170 316738 370226
rect 316806 370170 316862 370226
rect 316434 370046 316490 370102
rect 316558 370046 316614 370102
rect 316682 370046 316738 370102
rect 316806 370046 316862 370102
rect 316434 369922 316490 369978
rect 316558 369922 316614 369978
rect 316682 369922 316738 369978
rect 316806 369922 316862 369978
rect 316434 352294 316490 352350
rect 316558 352294 316614 352350
rect 316682 352294 316738 352350
rect 316806 352294 316862 352350
rect 316434 352170 316490 352226
rect 316558 352170 316614 352226
rect 316682 352170 316738 352226
rect 316806 352170 316862 352226
rect 316434 352046 316490 352102
rect 316558 352046 316614 352102
rect 316682 352046 316738 352102
rect 316806 352046 316862 352102
rect 316434 351922 316490 351978
rect 316558 351922 316614 351978
rect 316682 351922 316738 351978
rect 316806 351922 316862 351978
rect 316434 334294 316490 334350
rect 316558 334294 316614 334350
rect 316682 334294 316738 334350
rect 316806 334294 316862 334350
rect 316434 334170 316490 334226
rect 316558 334170 316614 334226
rect 316682 334170 316738 334226
rect 316806 334170 316862 334226
rect 316434 334046 316490 334102
rect 316558 334046 316614 334102
rect 316682 334046 316738 334102
rect 316806 334046 316862 334102
rect 316434 333922 316490 333978
rect 316558 333922 316614 333978
rect 316682 333922 316738 333978
rect 316806 333922 316862 333978
rect 316434 316294 316490 316350
rect 316558 316294 316614 316350
rect 316682 316294 316738 316350
rect 316806 316294 316862 316350
rect 316434 316170 316490 316226
rect 316558 316170 316614 316226
rect 316682 316170 316738 316226
rect 316806 316170 316862 316226
rect 316434 316046 316490 316102
rect 316558 316046 316614 316102
rect 316682 316046 316738 316102
rect 316806 316046 316862 316102
rect 316434 315922 316490 315978
rect 316558 315922 316614 315978
rect 316682 315922 316738 315978
rect 316806 315922 316862 315978
rect 316434 298294 316490 298350
rect 316558 298294 316614 298350
rect 316682 298294 316738 298350
rect 316806 298294 316862 298350
rect 316434 298170 316490 298226
rect 316558 298170 316614 298226
rect 316682 298170 316738 298226
rect 316806 298170 316862 298226
rect 316434 298046 316490 298102
rect 316558 298046 316614 298102
rect 316682 298046 316738 298102
rect 316806 298046 316862 298102
rect 316434 297922 316490 297978
rect 316558 297922 316614 297978
rect 316682 297922 316738 297978
rect 316806 297922 316862 297978
rect 316434 280294 316490 280350
rect 316558 280294 316614 280350
rect 316682 280294 316738 280350
rect 316806 280294 316862 280350
rect 316434 280170 316490 280226
rect 316558 280170 316614 280226
rect 316682 280170 316738 280226
rect 316806 280170 316862 280226
rect 316434 280046 316490 280102
rect 316558 280046 316614 280102
rect 316682 280046 316738 280102
rect 316806 280046 316862 280102
rect 316434 279922 316490 279978
rect 316558 279922 316614 279978
rect 316682 279922 316738 279978
rect 316806 279922 316862 279978
rect 316434 262294 316490 262350
rect 316558 262294 316614 262350
rect 316682 262294 316738 262350
rect 316806 262294 316862 262350
rect 316434 262170 316490 262226
rect 316558 262170 316614 262226
rect 316682 262170 316738 262226
rect 316806 262170 316862 262226
rect 316434 262046 316490 262102
rect 316558 262046 316614 262102
rect 316682 262046 316738 262102
rect 316806 262046 316862 262102
rect 316434 261922 316490 261978
rect 316558 261922 316614 261978
rect 316682 261922 316738 261978
rect 316806 261922 316862 261978
rect 316434 244294 316490 244350
rect 316558 244294 316614 244350
rect 316682 244294 316738 244350
rect 316806 244294 316862 244350
rect 316434 244170 316490 244226
rect 316558 244170 316614 244226
rect 316682 244170 316738 244226
rect 316806 244170 316862 244226
rect 316434 244046 316490 244102
rect 316558 244046 316614 244102
rect 316682 244046 316738 244102
rect 316806 244046 316862 244102
rect 316434 243922 316490 243978
rect 316558 243922 316614 243978
rect 316682 243922 316738 243978
rect 316806 243922 316862 243978
rect 316434 226294 316490 226350
rect 316558 226294 316614 226350
rect 316682 226294 316738 226350
rect 316806 226294 316862 226350
rect 316434 226170 316490 226226
rect 316558 226170 316614 226226
rect 316682 226170 316738 226226
rect 316806 226170 316862 226226
rect 316434 226046 316490 226102
rect 316558 226046 316614 226102
rect 316682 226046 316738 226102
rect 316806 226046 316862 226102
rect 316434 225922 316490 225978
rect 316558 225922 316614 225978
rect 316682 225922 316738 225978
rect 316806 225922 316862 225978
rect 316434 208294 316490 208350
rect 316558 208294 316614 208350
rect 316682 208294 316738 208350
rect 316806 208294 316862 208350
rect 316434 208170 316490 208226
rect 316558 208170 316614 208226
rect 316682 208170 316738 208226
rect 316806 208170 316862 208226
rect 316434 208046 316490 208102
rect 316558 208046 316614 208102
rect 316682 208046 316738 208102
rect 316806 208046 316862 208102
rect 316434 207922 316490 207978
rect 316558 207922 316614 207978
rect 316682 207922 316738 207978
rect 316806 207922 316862 207978
rect 316434 190294 316490 190350
rect 316558 190294 316614 190350
rect 316682 190294 316738 190350
rect 316806 190294 316862 190350
rect 316434 190170 316490 190226
rect 316558 190170 316614 190226
rect 316682 190170 316738 190226
rect 316806 190170 316862 190226
rect 316434 190046 316490 190102
rect 316558 190046 316614 190102
rect 316682 190046 316738 190102
rect 316806 190046 316862 190102
rect 316434 189922 316490 189978
rect 316558 189922 316614 189978
rect 316682 189922 316738 189978
rect 316806 189922 316862 189978
rect 316434 172294 316490 172350
rect 316558 172294 316614 172350
rect 316682 172294 316738 172350
rect 316806 172294 316862 172350
rect 316434 172170 316490 172226
rect 316558 172170 316614 172226
rect 316682 172170 316738 172226
rect 316806 172170 316862 172226
rect 316434 172046 316490 172102
rect 316558 172046 316614 172102
rect 316682 172046 316738 172102
rect 316806 172046 316862 172102
rect 316434 171922 316490 171978
rect 316558 171922 316614 171978
rect 316682 171922 316738 171978
rect 316806 171922 316862 171978
rect 316434 154294 316490 154350
rect 316558 154294 316614 154350
rect 316682 154294 316738 154350
rect 316806 154294 316862 154350
rect 316434 154170 316490 154226
rect 316558 154170 316614 154226
rect 316682 154170 316738 154226
rect 316806 154170 316862 154226
rect 316434 154046 316490 154102
rect 316558 154046 316614 154102
rect 316682 154046 316738 154102
rect 316806 154046 316862 154102
rect 316434 153922 316490 153978
rect 316558 153922 316614 153978
rect 316682 153922 316738 153978
rect 316806 153922 316862 153978
rect 316434 136294 316490 136350
rect 316558 136294 316614 136350
rect 316682 136294 316738 136350
rect 316806 136294 316862 136350
rect 316434 136170 316490 136226
rect 316558 136170 316614 136226
rect 316682 136170 316738 136226
rect 316806 136170 316862 136226
rect 316434 136046 316490 136102
rect 316558 136046 316614 136102
rect 316682 136046 316738 136102
rect 316806 136046 316862 136102
rect 316434 135922 316490 135978
rect 316558 135922 316614 135978
rect 316682 135922 316738 135978
rect 316806 135922 316862 135978
rect 316434 118294 316490 118350
rect 316558 118294 316614 118350
rect 316682 118294 316738 118350
rect 316806 118294 316862 118350
rect 316434 118170 316490 118226
rect 316558 118170 316614 118226
rect 316682 118170 316738 118226
rect 316806 118170 316862 118226
rect 316434 118046 316490 118102
rect 316558 118046 316614 118102
rect 316682 118046 316738 118102
rect 316806 118046 316862 118102
rect 316434 117922 316490 117978
rect 316558 117922 316614 117978
rect 316682 117922 316738 117978
rect 316806 117922 316862 117978
rect 316434 100294 316490 100350
rect 316558 100294 316614 100350
rect 316682 100294 316738 100350
rect 316806 100294 316862 100350
rect 316434 100170 316490 100226
rect 316558 100170 316614 100226
rect 316682 100170 316738 100226
rect 316806 100170 316862 100226
rect 316434 100046 316490 100102
rect 316558 100046 316614 100102
rect 316682 100046 316738 100102
rect 316806 100046 316862 100102
rect 316434 99922 316490 99978
rect 316558 99922 316614 99978
rect 316682 99922 316738 99978
rect 316806 99922 316862 99978
rect 316434 82294 316490 82350
rect 316558 82294 316614 82350
rect 316682 82294 316738 82350
rect 316806 82294 316862 82350
rect 316434 82170 316490 82226
rect 316558 82170 316614 82226
rect 316682 82170 316738 82226
rect 316806 82170 316862 82226
rect 316434 82046 316490 82102
rect 316558 82046 316614 82102
rect 316682 82046 316738 82102
rect 316806 82046 316862 82102
rect 316434 81922 316490 81978
rect 316558 81922 316614 81978
rect 316682 81922 316738 81978
rect 316806 81922 316862 81978
rect 341068 79802 341124 79858
rect 343434 580294 343490 580350
rect 343558 580294 343614 580350
rect 343682 580294 343738 580350
rect 343806 580294 343862 580350
rect 343434 580170 343490 580226
rect 343558 580170 343614 580226
rect 343682 580170 343738 580226
rect 343806 580170 343862 580226
rect 343434 580046 343490 580102
rect 343558 580046 343614 580102
rect 343682 580046 343738 580102
rect 343806 580046 343862 580102
rect 343434 579922 343490 579978
rect 343558 579922 343614 579978
rect 343682 579922 343738 579978
rect 343806 579922 343862 579978
rect 343434 562294 343490 562350
rect 343558 562294 343614 562350
rect 343682 562294 343738 562350
rect 343806 562294 343862 562350
rect 343434 562170 343490 562226
rect 343558 562170 343614 562226
rect 343682 562170 343738 562226
rect 343806 562170 343862 562226
rect 343434 562046 343490 562102
rect 343558 562046 343614 562102
rect 343682 562046 343738 562102
rect 343806 562046 343862 562102
rect 343434 561922 343490 561978
rect 343558 561922 343614 561978
rect 343682 561922 343738 561978
rect 343806 561922 343862 561978
rect 343434 544294 343490 544350
rect 343558 544294 343614 544350
rect 343682 544294 343738 544350
rect 343806 544294 343862 544350
rect 343434 544170 343490 544226
rect 343558 544170 343614 544226
rect 343682 544170 343738 544226
rect 343806 544170 343862 544226
rect 343434 544046 343490 544102
rect 343558 544046 343614 544102
rect 343682 544046 343738 544102
rect 343806 544046 343862 544102
rect 343434 543922 343490 543978
rect 343558 543922 343614 543978
rect 343682 543922 343738 543978
rect 343806 543922 343862 543978
rect 343434 526294 343490 526350
rect 343558 526294 343614 526350
rect 343682 526294 343738 526350
rect 343806 526294 343862 526350
rect 343434 526170 343490 526226
rect 343558 526170 343614 526226
rect 343682 526170 343738 526226
rect 343806 526170 343862 526226
rect 343434 526046 343490 526102
rect 343558 526046 343614 526102
rect 343682 526046 343738 526102
rect 343806 526046 343862 526102
rect 343434 525922 343490 525978
rect 343558 525922 343614 525978
rect 343682 525922 343738 525978
rect 343806 525922 343862 525978
rect 343434 508294 343490 508350
rect 343558 508294 343614 508350
rect 343682 508294 343738 508350
rect 343806 508294 343862 508350
rect 343434 508170 343490 508226
rect 343558 508170 343614 508226
rect 343682 508170 343738 508226
rect 343806 508170 343862 508226
rect 343434 508046 343490 508102
rect 343558 508046 343614 508102
rect 343682 508046 343738 508102
rect 343806 508046 343862 508102
rect 343434 507922 343490 507978
rect 343558 507922 343614 507978
rect 343682 507922 343738 507978
rect 343806 507922 343862 507978
rect 343434 490294 343490 490350
rect 343558 490294 343614 490350
rect 343682 490294 343738 490350
rect 343806 490294 343862 490350
rect 343434 490170 343490 490226
rect 343558 490170 343614 490226
rect 343682 490170 343738 490226
rect 343806 490170 343862 490226
rect 343434 490046 343490 490102
rect 343558 490046 343614 490102
rect 343682 490046 343738 490102
rect 343806 490046 343862 490102
rect 343434 489922 343490 489978
rect 343558 489922 343614 489978
rect 343682 489922 343738 489978
rect 343806 489922 343862 489978
rect 343434 472294 343490 472350
rect 343558 472294 343614 472350
rect 343682 472294 343738 472350
rect 343806 472294 343862 472350
rect 343434 472170 343490 472226
rect 343558 472170 343614 472226
rect 343682 472170 343738 472226
rect 343806 472170 343862 472226
rect 343434 472046 343490 472102
rect 343558 472046 343614 472102
rect 343682 472046 343738 472102
rect 343806 472046 343862 472102
rect 343434 471922 343490 471978
rect 343558 471922 343614 471978
rect 343682 471922 343738 471978
rect 343806 471922 343862 471978
rect 343434 454294 343490 454350
rect 343558 454294 343614 454350
rect 343682 454294 343738 454350
rect 343806 454294 343862 454350
rect 343434 454170 343490 454226
rect 343558 454170 343614 454226
rect 343682 454170 343738 454226
rect 343806 454170 343862 454226
rect 343434 454046 343490 454102
rect 343558 454046 343614 454102
rect 343682 454046 343738 454102
rect 343806 454046 343862 454102
rect 343434 453922 343490 453978
rect 343558 453922 343614 453978
rect 343682 453922 343738 453978
rect 343806 453922 343862 453978
rect 343434 436294 343490 436350
rect 343558 436294 343614 436350
rect 343682 436294 343738 436350
rect 343806 436294 343862 436350
rect 343434 436170 343490 436226
rect 343558 436170 343614 436226
rect 343682 436170 343738 436226
rect 343806 436170 343862 436226
rect 343434 436046 343490 436102
rect 343558 436046 343614 436102
rect 343682 436046 343738 436102
rect 343806 436046 343862 436102
rect 343434 435922 343490 435978
rect 343558 435922 343614 435978
rect 343682 435922 343738 435978
rect 343806 435922 343862 435978
rect 343434 418294 343490 418350
rect 343558 418294 343614 418350
rect 343682 418294 343738 418350
rect 343806 418294 343862 418350
rect 343434 418170 343490 418226
rect 343558 418170 343614 418226
rect 343682 418170 343738 418226
rect 343806 418170 343862 418226
rect 343434 418046 343490 418102
rect 343558 418046 343614 418102
rect 343682 418046 343738 418102
rect 343806 418046 343862 418102
rect 343434 417922 343490 417978
rect 343558 417922 343614 417978
rect 343682 417922 343738 417978
rect 343806 417922 343862 417978
rect 343434 400294 343490 400350
rect 343558 400294 343614 400350
rect 343682 400294 343738 400350
rect 343806 400294 343862 400350
rect 343434 400170 343490 400226
rect 343558 400170 343614 400226
rect 343682 400170 343738 400226
rect 343806 400170 343862 400226
rect 343434 400046 343490 400102
rect 343558 400046 343614 400102
rect 343682 400046 343738 400102
rect 343806 400046 343862 400102
rect 343434 399922 343490 399978
rect 343558 399922 343614 399978
rect 343682 399922 343738 399978
rect 343806 399922 343862 399978
rect 343434 382294 343490 382350
rect 343558 382294 343614 382350
rect 343682 382294 343738 382350
rect 343806 382294 343862 382350
rect 343434 382170 343490 382226
rect 343558 382170 343614 382226
rect 343682 382170 343738 382226
rect 343806 382170 343862 382226
rect 343434 382046 343490 382102
rect 343558 382046 343614 382102
rect 343682 382046 343738 382102
rect 343806 382046 343862 382102
rect 343434 381922 343490 381978
rect 343558 381922 343614 381978
rect 343682 381922 343738 381978
rect 343806 381922 343862 381978
rect 343434 364294 343490 364350
rect 343558 364294 343614 364350
rect 343682 364294 343738 364350
rect 343806 364294 343862 364350
rect 343434 364170 343490 364226
rect 343558 364170 343614 364226
rect 343682 364170 343738 364226
rect 343806 364170 343862 364226
rect 343434 364046 343490 364102
rect 343558 364046 343614 364102
rect 343682 364046 343738 364102
rect 343806 364046 343862 364102
rect 343434 363922 343490 363978
rect 343558 363922 343614 363978
rect 343682 363922 343738 363978
rect 343806 363922 343862 363978
rect 343434 346294 343490 346350
rect 343558 346294 343614 346350
rect 343682 346294 343738 346350
rect 343806 346294 343862 346350
rect 343434 346170 343490 346226
rect 343558 346170 343614 346226
rect 343682 346170 343738 346226
rect 343806 346170 343862 346226
rect 343434 346046 343490 346102
rect 343558 346046 343614 346102
rect 343682 346046 343738 346102
rect 343806 346046 343862 346102
rect 343434 345922 343490 345978
rect 343558 345922 343614 345978
rect 343682 345922 343738 345978
rect 343806 345922 343862 345978
rect 343434 328294 343490 328350
rect 343558 328294 343614 328350
rect 343682 328294 343738 328350
rect 343806 328294 343862 328350
rect 343434 328170 343490 328226
rect 343558 328170 343614 328226
rect 343682 328170 343738 328226
rect 343806 328170 343862 328226
rect 343434 328046 343490 328102
rect 343558 328046 343614 328102
rect 343682 328046 343738 328102
rect 343806 328046 343862 328102
rect 343434 327922 343490 327978
rect 343558 327922 343614 327978
rect 343682 327922 343738 327978
rect 343806 327922 343862 327978
rect 343434 310294 343490 310350
rect 343558 310294 343614 310350
rect 343682 310294 343738 310350
rect 343806 310294 343862 310350
rect 343434 310170 343490 310226
rect 343558 310170 343614 310226
rect 343682 310170 343738 310226
rect 343806 310170 343862 310226
rect 343434 310046 343490 310102
rect 343558 310046 343614 310102
rect 343682 310046 343738 310102
rect 343806 310046 343862 310102
rect 343434 309922 343490 309978
rect 343558 309922 343614 309978
rect 343682 309922 343738 309978
rect 343806 309922 343862 309978
rect 343434 292294 343490 292350
rect 343558 292294 343614 292350
rect 343682 292294 343738 292350
rect 343806 292294 343862 292350
rect 343434 292170 343490 292226
rect 343558 292170 343614 292226
rect 343682 292170 343738 292226
rect 343806 292170 343862 292226
rect 343434 292046 343490 292102
rect 343558 292046 343614 292102
rect 343682 292046 343738 292102
rect 343806 292046 343862 292102
rect 343434 291922 343490 291978
rect 343558 291922 343614 291978
rect 343682 291922 343738 291978
rect 343806 291922 343862 291978
rect 343434 274294 343490 274350
rect 343558 274294 343614 274350
rect 343682 274294 343738 274350
rect 343806 274294 343862 274350
rect 343434 274170 343490 274226
rect 343558 274170 343614 274226
rect 343682 274170 343738 274226
rect 343806 274170 343862 274226
rect 343434 274046 343490 274102
rect 343558 274046 343614 274102
rect 343682 274046 343738 274102
rect 343806 274046 343862 274102
rect 343434 273922 343490 273978
rect 343558 273922 343614 273978
rect 343682 273922 343738 273978
rect 343806 273922 343862 273978
rect 343434 256294 343490 256350
rect 343558 256294 343614 256350
rect 343682 256294 343738 256350
rect 343806 256294 343862 256350
rect 343434 256170 343490 256226
rect 343558 256170 343614 256226
rect 343682 256170 343738 256226
rect 343806 256170 343862 256226
rect 343434 256046 343490 256102
rect 343558 256046 343614 256102
rect 343682 256046 343738 256102
rect 343806 256046 343862 256102
rect 343434 255922 343490 255978
rect 343558 255922 343614 255978
rect 343682 255922 343738 255978
rect 343806 255922 343862 255978
rect 343434 238294 343490 238350
rect 343558 238294 343614 238350
rect 343682 238294 343738 238350
rect 343806 238294 343862 238350
rect 343434 238170 343490 238226
rect 343558 238170 343614 238226
rect 343682 238170 343738 238226
rect 343806 238170 343862 238226
rect 343434 238046 343490 238102
rect 343558 238046 343614 238102
rect 343682 238046 343738 238102
rect 343806 238046 343862 238102
rect 343434 237922 343490 237978
rect 343558 237922 343614 237978
rect 343682 237922 343738 237978
rect 343806 237922 343862 237978
rect 343434 220294 343490 220350
rect 343558 220294 343614 220350
rect 343682 220294 343738 220350
rect 343806 220294 343862 220350
rect 343434 220170 343490 220226
rect 343558 220170 343614 220226
rect 343682 220170 343738 220226
rect 343806 220170 343862 220226
rect 343434 220046 343490 220102
rect 343558 220046 343614 220102
rect 343682 220046 343738 220102
rect 343806 220046 343862 220102
rect 343434 219922 343490 219978
rect 343558 219922 343614 219978
rect 343682 219922 343738 219978
rect 343806 219922 343862 219978
rect 343434 202294 343490 202350
rect 343558 202294 343614 202350
rect 343682 202294 343738 202350
rect 343806 202294 343862 202350
rect 343434 202170 343490 202226
rect 343558 202170 343614 202226
rect 343682 202170 343738 202226
rect 343806 202170 343862 202226
rect 343434 202046 343490 202102
rect 343558 202046 343614 202102
rect 343682 202046 343738 202102
rect 343806 202046 343862 202102
rect 343434 201922 343490 201978
rect 343558 201922 343614 201978
rect 343682 201922 343738 201978
rect 343806 201922 343862 201978
rect 343434 184294 343490 184350
rect 343558 184294 343614 184350
rect 343682 184294 343738 184350
rect 343806 184294 343862 184350
rect 343434 184170 343490 184226
rect 343558 184170 343614 184226
rect 343682 184170 343738 184226
rect 343806 184170 343862 184226
rect 343434 184046 343490 184102
rect 343558 184046 343614 184102
rect 343682 184046 343738 184102
rect 343806 184046 343862 184102
rect 343434 183922 343490 183978
rect 343558 183922 343614 183978
rect 343682 183922 343738 183978
rect 343806 183922 343862 183978
rect 343434 166294 343490 166350
rect 343558 166294 343614 166350
rect 343682 166294 343738 166350
rect 343806 166294 343862 166350
rect 343434 166170 343490 166226
rect 343558 166170 343614 166226
rect 343682 166170 343738 166226
rect 343806 166170 343862 166226
rect 343434 166046 343490 166102
rect 343558 166046 343614 166102
rect 343682 166046 343738 166102
rect 343806 166046 343862 166102
rect 343434 165922 343490 165978
rect 343558 165922 343614 165978
rect 343682 165922 343738 165978
rect 343806 165922 343862 165978
rect 343434 148294 343490 148350
rect 343558 148294 343614 148350
rect 343682 148294 343738 148350
rect 343806 148294 343862 148350
rect 343434 148170 343490 148226
rect 343558 148170 343614 148226
rect 343682 148170 343738 148226
rect 343806 148170 343862 148226
rect 343434 148046 343490 148102
rect 343558 148046 343614 148102
rect 343682 148046 343738 148102
rect 343806 148046 343862 148102
rect 343434 147922 343490 147978
rect 343558 147922 343614 147978
rect 343682 147922 343738 147978
rect 343806 147922 343862 147978
rect 343434 130294 343490 130350
rect 343558 130294 343614 130350
rect 343682 130294 343738 130350
rect 343806 130294 343862 130350
rect 343434 130170 343490 130226
rect 343558 130170 343614 130226
rect 343682 130170 343738 130226
rect 343806 130170 343862 130226
rect 343434 130046 343490 130102
rect 343558 130046 343614 130102
rect 343682 130046 343738 130102
rect 343806 130046 343862 130102
rect 343434 129922 343490 129978
rect 343558 129922 343614 129978
rect 343682 129922 343738 129978
rect 343806 129922 343862 129978
rect 343434 112294 343490 112350
rect 343558 112294 343614 112350
rect 343682 112294 343738 112350
rect 343806 112294 343862 112350
rect 343434 112170 343490 112226
rect 343558 112170 343614 112226
rect 343682 112170 343738 112226
rect 343806 112170 343862 112226
rect 343434 112046 343490 112102
rect 343558 112046 343614 112102
rect 343682 112046 343738 112102
rect 343806 112046 343862 112102
rect 343434 111922 343490 111978
rect 343558 111922 343614 111978
rect 343682 111922 343738 111978
rect 343806 111922 343862 111978
rect 343434 94294 343490 94350
rect 343558 94294 343614 94350
rect 343682 94294 343738 94350
rect 343806 94294 343862 94350
rect 343434 94170 343490 94226
rect 343558 94170 343614 94226
rect 343682 94170 343738 94226
rect 343806 94170 343862 94226
rect 343434 94046 343490 94102
rect 343558 94046 343614 94102
rect 343682 94046 343738 94102
rect 343806 94046 343862 94102
rect 343434 93922 343490 93978
rect 343558 93922 343614 93978
rect 343682 93922 343738 93978
rect 343806 93922 343862 93978
rect 343434 76294 343490 76350
rect 343558 76294 343614 76350
rect 343682 76294 343738 76350
rect 343806 76294 343862 76350
rect 343434 76170 343490 76226
rect 343558 76170 343614 76226
rect 343682 76170 343738 76226
rect 343806 76170 343862 76226
rect 343434 76046 343490 76102
rect 343558 76046 343614 76102
rect 343682 76046 343738 76102
rect 343806 76046 343862 76102
rect 343434 75922 343490 75978
rect 343558 75922 343614 75978
rect 343682 75922 343738 75978
rect 343806 75922 343862 75978
rect 316434 64294 316490 64350
rect 316558 64294 316614 64350
rect 316682 64294 316738 64350
rect 316806 64294 316862 64350
rect 316434 64170 316490 64226
rect 316558 64170 316614 64226
rect 316682 64170 316738 64226
rect 316806 64170 316862 64226
rect 316434 64046 316490 64102
rect 316558 64046 316614 64102
rect 316682 64046 316738 64102
rect 316806 64046 316862 64102
rect 316434 63922 316490 63978
rect 316558 63922 316614 63978
rect 316682 63922 316738 63978
rect 316806 63922 316862 63978
rect 316434 46294 316490 46350
rect 316558 46294 316614 46350
rect 316682 46294 316738 46350
rect 316806 46294 316862 46350
rect 316434 46170 316490 46226
rect 316558 46170 316614 46226
rect 316682 46170 316738 46226
rect 316806 46170 316862 46226
rect 316434 46046 316490 46102
rect 316558 46046 316614 46102
rect 316682 46046 316738 46102
rect 316806 46046 316862 46102
rect 316434 45922 316490 45978
rect 316558 45922 316614 45978
rect 316682 45922 316738 45978
rect 316806 45922 316862 45978
rect 316434 28294 316490 28350
rect 316558 28294 316614 28350
rect 316682 28294 316738 28350
rect 316806 28294 316862 28350
rect 316434 28170 316490 28226
rect 316558 28170 316614 28226
rect 316682 28170 316738 28226
rect 316806 28170 316862 28226
rect 316434 28046 316490 28102
rect 316558 28046 316614 28102
rect 316682 28046 316738 28102
rect 316806 28046 316862 28102
rect 316434 27922 316490 27978
rect 316558 27922 316614 27978
rect 316682 27922 316738 27978
rect 316806 27922 316862 27978
rect 312714 22294 312770 22350
rect 312838 22294 312894 22350
rect 312962 22294 313018 22350
rect 313086 22294 313142 22350
rect 312714 22170 312770 22226
rect 312838 22170 312894 22226
rect 312962 22170 313018 22226
rect 313086 22170 313142 22226
rect 312714 22046 312770 22102
rect 312838 22046 312894 22102
rect 312962 22046 313018 22102
rect 313086 22046 313142 22102
rect 312714 21922 312770 21978
rect 312838 21922 312894 21978
rect 312962 21922 313018 21978
rect 313086 21922 313142 21978
rect 312714 4294 312770 4350
rect 312838 4294 312894 4350
rect 312962 4294 313018 4350
rect 313086 4294 313142 4350
rect 312714 4170 312770 4226
rect 312838 4170 312894 4226
rect 312962 4170 313018 4226
rect 313086 4170 313142 4226
rect 314188 22742 314244 22798
rect 316434 10294 316490 10350
rect 316558 10294 316614 10350
rect 316682 10294 316738 10350
rect 316806 10294 316862 10350
rect 316434 10170 316490 10226
rect 316558 10170 316614 10226
rect 316682 10170 316738 10226
rect 316806 10170 316862 10226
rect 316434 10046 316490 10102
rect 316558 10046 316614 10102
rect 316682 10046 316738 10102
rect 316806 10046 316862 10102
rect 316434 9922 316490 9978
rect 316558 9922 316614 9978
rect 316682 9922 316738 9978
rect 316806 9922 316862 9978
rect 312714 4046 312770 4102
rect 312838 4046 312894 4102
rect 312962 4046 313018 4102
rect 313086 4046 313142 4102
rect 312714 3922 312770 3978
rect 312838 3922 312894 3978
rect 312962 3922 313018 3978
rect 313086 3922 313142 3978
rect 285714 -1176 285770 -1120
rect 285838 -1176 285894 -1120
rect 285962 -1176 286018 -1120
rect 286086 -1176 286142 -1120
rect 285714 -1300 285770 -1244
rect 285838 -1300 285894 -1244
rect 285962 -1300 286018 -1244
rect 286086 -1300 286142 -1244
rect 285714 -1424 285770 -1368
rect 285838 -1424 285894 -1368
rect 285962 -1424 286018 -1368
rect 286086 -1424 286142 -1368
rect 285714 -1548 285770 -1492
rect 285838 -1548 285894 -1492
rect 285962 -1548 286018 -1492
rect 286086 -1548 286142 -1492
rect 312714 -216 312770 -160
rect 312838 -216 312894 -160
rect 312962 -216 313018 -160
rect 313086 -216 313142 -160
rect 312714 -340 312770 -284
rect 312838 -340 312894 -284
rect 312962 -340 313018 -284
rect 313086 -340 313142 -284
rect 312714 -464 312770 -408
rect 312838 -464 312894 -408
rect 312962 -464 313018 -408
rect 313086 -464 313142 -408
rect 312714 -588 312770 -532
rect 312838 -588 312894 -532
rect 312962 -588 313018 -532
rect 313086 -588 313142 -532
rect 317548 65942 317604 65998
rect 324268 62522 324324 62578
rect 322588 59462 322644 59518
rect 319228 44342 319284 44398
rect 343434 58294 343490 58350
rect 343558 58294 343614 58350
rect 343682 58294 343738 58350
rect 343806 58294 343862 58350
rect 343434 58170 343490 58226
rect 343558 58170 343614 58226
rect 343682 58170 343738 58226
rect 343806 58170 343862 58226
rect 343434 58046 343490 58102
rect 343558 58046 343614 58102
rect 343682 58046 343738 58102
rect 343806 58046 343862 58102
rect 343434 57922 343490 57978
rect 343558 57922 343614 57978
rect 343682 57922 343738 57978
rect 343806 57922 343862 57978
rect 330988 40742 331044 40798
rect 347154 598116 347210 598172
rect 347278 598116 347334 598172
rect 347402 598116 347458 598172
rect 347526 598116 347582 598172
rect 347154 597992 347210 598048
rect 347278 597992 347334 598048
rect 347402 597992 347458 598048
rect 347526 597992 347582 598048
rect 347154 597868 347210 597924
rect 347278 597868 347334 597924
rect 347402 597868 347458 597924
rect 347526 597868 347582 597924
rect 347154 597744 347210 597800
rect 347278 597744 347334 597800
rect 347402 597744 347458 597800
rect 347526 597744 347582 597800
rect 347154 586294 347210 586350
rect 347278 586294 347334 586350
rect 347402 586294 347458 586350
rect 347526 586294 347582 586350
rect 347154 586170 347210 586226
rect 347278 586170 347334 586226
rect 347402 586170 347458 586226
rect 347526 586170 347582 586226
rect 347154 586046 347210 586102
rect 347278 586046 347334 586102
rect 347402 586046 347458 586102
rect 347526 586046 347582 586102
rect 347154 585922 347210 585978
rect 347278 585922 347334 585978
rect 347402 585922 347458 585978
rect 347526 585922 347582 585978
rect 347154 568294 347210 568350
rect 347278 568294 347334 568350
rect 347402 568294 347458 568350
rect 347526 568294 347582 568350
rect 347154 568170 347210 568226
rect 347278 568170 347334 568226
rect 347402 568170 347458 568226
rect 347526 568170 347582 568226
rect 347154 568046 347210 568102
rect 347278 568046 347334 568102
rect 347402 568046 347458 568102
rect 347526 568046 347582 568102
rect 347154 567922 347210 567978
rect 347278 567922 347334 567978
rect 347402 567922 347458 567978
rect 347526 567922 347582 567978
rect 347154 550294 347210 550350
rect 347278 550294 347334 550350
rect 347402 550294 347458 550350
rect 347526 550294 347582 550350
rect 347154 550170 347210 550226
rect 347278 550170 347334 550226
rect 347402 550170 347458 550226
rect 347526 550170 347582 550226
rect 347154 550046 347210 550102
rect 347278 550046 347334 550102
rect 347402 550046 347458 550102
rect 347526 550046 347582 550102
rect 347154 549922 347210 549978
rect 347278 549922 347334 549978
rect 347402 549922 347458 549978
rect 347526 549922 347582 549978
rect 347154 532294 347210 532350
rect 347278 532294 347334 532350
rect 347402 532294 347458 532350
rect 347526 532294 347582 532350
rect 347154 532170 347210 532226
rect 347278 532170 347334 532226
rect 347402 532170 347458 532226
rect 347526 532170 347582 532226
rect 347154 532046 347210 532102
rect 347278 532046 347334 532102
rect 347402 532046 347458 532102
rect 347526 532046 347582 532102
rect 347154 531922 347210 531978
rect 347278 531922 347334 531978
rect 347402 531922 347458 531978
rect 347526 531922 347582 531978
rect 347154 514294 347210 514350
rect 347278 514294 347334 514350
rect 347402 514294 347458 514350
rect 347526 514294 347582 514350
rect 347154 514170 347210 514226
rect 347278 514170 347334 514226
rect 347402 514170 347458 514226
rect 347526 514170 347582 514226
rect 347154 514046 347210 514102
rect 347278 514046 347334 514102
rect 347402 514046 347458 514102
rect 347526 514046 347582 514102
rect 347154 513922 347210 513978
rect 347278 513922 347334 513978
rect 347402 513922 347458 513978
rect 347526 513922 347582 513978
rect 347154 496294 347210 496350
rect 347278 496294 347334 496350
rect 347402 496294 347458 496350
rect 347526 496294 347582 496350
rect 347154 496170 347210 496226
rect 347278 496170 347334 496226
rect 347402 496170 347458 496226
rect 347526 496170 347582 496226
rect 347154 496046 347210 496102
rect 347278 496046 347334 496102
rect 347402 496046 347458 496102
rect 347526 496046 347582 496102
rect 347154 495922 347210 495978
rect 347278 495922 347334 495978
rect 347402 495922 347458 495978
rect 347526 495922 347582 495978
rect 347154 478294 347210 478350
rect 347278 478294 347334 478350
rect 347402 478294 347458 478350
rect 347526 478294 347582 478350
rect 347154 478170 347210 478226
rect 347278 478170 347334 478226
rect 347402 478170 347458 478226
rect 347526 478170 347582 478226
rect 347154 478046 347210 478102
rect 347278 478046 347334 478102
rect 347402 478046 347458 478102
rect 347526 478046 347582 478102
rect 347154 477922 347210 477978
rect 347278 477922 347334 477978
rect 347402 477922 347458 477978
rect 347526 477922 347582 477978
rect 347154 460294 347210 460350
rect 347278 460294 347334 460350
rect 347402 460294 347458 460350
rect 347526 460294 347582 460350
rect 347154 460170 347210 460226
rect 347278 460170 347334 460226
rect 347402 460170 347458 460226
rect 347526 460170 347582 460226
rect 347154 460046 347210 460102
rect 347278 460046 347334 460102
rect 347402 460046 347458 460102
rect 347526 460046 347582 460102
rect 347154 459922 347210 459978
rect 347278 459922 347334 459978
rect 347402 459922 347458 459978
rect 347526 459922 347582 459978
rect 347154 442294 347210 442350
rect 347278 442294 347334 442350
rect 347402 442294 347458 442350
rect 347526 442294 347582 442350
rect 347154 442170 347210 442226
rect 347278 442170 347334 442226
rect 347402 442170 347458 442226
rect 347526 442170 347582 442226
rect 347154 442046 347210 442102
rect 347278 442046 347334 442102
rect 347402 442046 347458 442102
rect 347526 442046 347582 442102
rect 347154 441922 347210 441978
rect 347278 441922 347334 441978
rect 347402 441922 347458 441978
rect 347526 441922 347582 441978
rect 347154 424294 347210 424350
rect 347278 424294 347334 424350
rect 347402 424294 347458 424350
rect 347526 424294 347582 424350
rect 347154 424170 347210 424226
rect 347278 424170 347334 424226
rect 347402 424170 347458 424226
rect 347526 424170 347582 424226
rect 347154 424046 347210 424102
rect 347278 424046 347334 424102
rect 347402 424046 347458 424102
rect 347526 424046 347582 424102
rect 347154 423922 347210 423978
rect 347278 423922 347334 423978
rect 347402 423922 347458 423978
rect 347526 423922 347582 423978
rect 347154 406294 347210 406350
rect 347278 406294 347334 406350
rect 347402 406294 347458 406350
rect 347526 406294 347582 406350
rect 347154 406170 347210 406226
rect 347278 406170 347334 406226
rect 347402 406170 347458 406226
rect 347526 406170 347582 406226
rect 347154 406046 347210 406102
rect 347278 406046 347334 406102
rect 347402 406046 347458 406102
rect 347526 406046 347582 406102
rect 347154 405922 347210 405978
rect 347278 405922 347334 405978
rect 347402 405922 347458 405978
rect 347526 405922 347582 405978
rect 347154 388294 347210 388350
rect 347278 388294 347334 388350
rect 347402 388294 347458 388350
rect 347526 388294 347582 388350
rect 347154 388170 347210 388226
rect 347278 388170 347334 388226
rect 347402 388170 347458 388226
rect 347526 388170 347582 388226
rect 347154 388046 347210 388102
rect 347278 388046 347334 388102
rect 347402 388046 347458 388102
rect 347526 388046 347582 388102
rect 347154 387922 347210 387978
rect 347278 387922 347334 387978
rect 347402 387922 347458 387978
rect 347526 387922 347582 387978
rect 347154 370294 347210 370350
rect 347278 370294 347334 370350
rect 347402 370294 347458 370350
rect 347526 370294 347582 370350
rect 347154 370170 347210 370226
rect 347278 370170 347334 370226
rect 347402 370170 347458 370226
rect 347526 370170 347582 370226
rect 347154 370046 347210 370102
rect 347278 370046 347334 370102
rect 347402 370046 347458 370102
rect 347526 370046 347582 370102
rect 347154 369922 347210 369978
rect 347278 369922 347334 369978
rect 347402 369922 347458 369978
rect 347526 369922 347582 369978
rect 347154 352294 347210 352350
rect 347278 352294 347334 352350
rect 347402 352294 347458 352350
rect 347526 352294 347582 352350
rect 347154 352170 347210 352226
rect 347278 352170 347334 352226
rect 347402 352170 347458 352226
rect 347526 352170 347582 352226
rect 347154 352046 347210 352102
rect 347278 352046 347334 352102
rect 347402 352046 347458 352102
rect 347526 352046 347582 352102
rect 347154 351922 347210 351978
rect 347278 351922 347334 351978
rect 347402 351922 347458 351978
rect 347526 351922 347582 351978
rect 347154 334294 347210 334350
rect 347278 334294 347334 334350
rect 347402 334294 347458 334350
rect 347526 334294 347582 334350
rect 347154 334170 347210 334226
rect 347278 334170 347334 334226
rect 347402 334170 347458 334226
rect 347526 334170 347582 334226
rect 347154 334046 347210 334102
rect 347278 334046 347334 334102
rect 347402 334046 347458 334102
rect 347526 334046 347582 334102
rect 347154 333922 347210 333978
rect 347278 333922 347334 333978
rect 347402 333922 347458 333978
rect 347526 333922 347582 333978
rect 347154 316294 347210 316350
rect 347278 316294 347334 316350
rect 347402 316294 347458 316350
rect 347526 316294 347582 316350
rect 347154 316170 347210 316226
rect 347278 316170 347334 316226
rect 347402 316170 347458 316226
rect 347526 316170 347582 316226
rect 347154 316046 347210 316102
rect 347278 316046 347334 316102
rect 347402 316046 347458 316102
rect 347526 316046 347582 316102
rect 347154 315922 347210 315978
rect 347278 315922 347334 315978
rect 347402 315922 347458 315978
rect 347526 315922 347582 315978
rect 347154 298294 347210 298350
rect 347278 298294 347334 298350
rect 347402 298294 347458 298350
rect 347526 298294 347582 298350
rect 347154 298170 347210 298226
rect 347278 298170 347334 298226
rect 347402 298170 347458 298226
rect 347526 298170 347582 298226
rect 347154 298046 347210 298102
rect 347278 298046 347334 298102
rect 347402 298046 347458 298102
rect 347526 298046 347582 298102
rect 347154 297922 347210 297978
rect 347278 297922 347334 297978
rect 347402 297922 347458 297978
rect 347526 297922 347582 297978
rect 347154 280294 347210 280350
rect 347278 280294 347334 280350
rect 347402 280294 347458 280350
rect 347526 280294 347582 280350
rect 347154 280170 347210 280226
rect 347278 280170 347334 280226
rect 347402 280170 347458 280226
rect 347526 280170 347582 280226
rect 347154 280046 347210 280102
rect 347278 280046 347334 280102
rect 347402 280046 347458 280102
rect 347526 280046 347582 280102
rect 347154 279922 347210 279978
rect 347278 279922 347334 279978
rect 347402 279922 347458 279978
rect 347526 279922 347582 279978
rect 347154 262294 347210 262350
rect 347278 262294 347334 262350
rect 347402 262294 347458 262350
rect 347526 262294 347582 262350
rect 347154 262170 347210 262226
rect 347278 262170 347334 262226
rect 347402 262170 347458 262226
rect 347526 262170 347582 262226
rect 347154 262046 347210 262102
rect 347278 262046 347334 262102
rect 347402 262046 347458 262102
rect 347526 262046 347582 262102
rect 347154 261922 347210 261978
rect 347278 261922 347334 261978
rect 347402 261922 347458 261978
rect 347526 261922 347582 261978
rect 347154 244294 347210 244350
rect 347278 244294 347334 244350
rect 347402 244294 347458 244350
rect 347526 244294 347582 244350
rect 347154 244170 347210 244226
rect 347278 244170 347334 244226
rect 347402 244170 347458 244226
rect 347526 244170 347582 244226
rect 347154 244046 347210 244102
rect 347278 244046 347334 244102
rect 347402 244046 347458 244102
rect 347526 244046 347582 244102
rect 347154 243922 347210 243978
rect 347278 243922 347334 243978
rect 347402 243922 347458 243978
rect 347526 243922 347582 243978
rect 347154 226294 347210 226350
rect 347278 226294 347334 226350
rect 347402 226294 347458 226350
rect 347526 226294 347582 226350
rect 347154 226170 347210 226226
rect 347278 226170 347334 226226
rect 347402 226170 347458 226226
rect 347526 226170 347582 226226
rect 347154 226046 347210 226102
rect 347278 226046 347334 226102
rect 347402 226046 347458 226102
rect 347526 226046 347582 226102
rect 347154 225922 347210 225978
rect 347278 225922 347334 225978
rect 347402 225922 347458 225978
rect 347526 225922 347582 225978
rect 347154 208294 347210 208350
rect 347278 208294 347334 208350
rect 347402 208294 347458 208350
rect 347526 208294 347582 208350
rect 347154 208170 347210 208226
rect 347278 208170 347334 208226
rect 347402 208170 347458 208226
rect 347526 208170 347582 208226
rect 347154 208046 347210 208102
rect 347278 208046 347334 208102
rect 347402 208046 347458 208102
rect 347526 208046 347582 208102
rect 347154 207922 347210 207978
rect 347278 207922 347334 207978
rect 347402 207922 347458 207978
rect 347526 207922 347582 207978
rect 347154 190294 347210 190350
rect 347278 190294 347334 190350
rect 347402 190294 347458 190350
rect 347526 190294 347582 190350
rect 347154 190170 347210 190226
rect 347278 190170 347334 190226
rect 347402 190170 347458 190226
rect 347526 190170 347582 190226
rect 347154 190046 347210 190102
rect 347278 190046 347334 190102
rect 347402 190046 347458 190102
rect 347526 190046 347582 190102
rect 347154 189922 347210 189978
rect 347278 189922 347334 189978
rect 347402 189922 347458 189978
rect 347526 189922 347582 189978
rect 347154 172294 347210 172350
rect 347278 172294 347334 172350
rect 347402 172294 347458 172350
rect 347526 172294 347582 172350
rect 347154 172170 347210 172226
rect 347278 172170 347334 172226
rect 347402 172170 347458 172226
rect 347526 172170 347582 172226
rect 347154 172046 347210 172102
rect 347278 172046 347334 172102
rect 347402 172046 347458 172102
rect 347526 172046 347582 172102
rect 347154 171922 347210 171978
rect 347278 171922 347334 171978
rect 347402 171922 347458 171978
rect 347526 171922 347582 171978
rect 347154 154294 347210 154350
rect 347278 154294 347334 154350
rect 347402 154294 347458 154350
rect 347526 154294 347582 154350
rect 347154 154170 347210 154226
rect 347278 154170 347334 154226
rect 347402 154170 347458 154226
rect 347526 154170 347582 154226
rect 347154 154046 347210 154102
rect 347278 154046 347334 154102
rect 347402 154046 347458 154102
rect 347526 154046 347582 154102
rect 347154 153922 347210 153978
rect 347278 153922 347334 153978
rect 347402 153922 347458 153978
rect 347526 153922 347582 153978
rect 347154 136294 347210 136350
rect 347278 136294 347334 136350
rect 347402 136294 347458 136350
rect 347526 136294 347582 136350
rect 347154 136170 347210 136226
rect 347278 136170 347334 136226
rect 347402 136170 347458 136226
rect 347526 136170 347582 136226
rect 347154 136046 347210 136102
rect 347278 136046 347334 136102
rect 347402 136046 347458 136102
rect 347526 136046 347582 136102
rect 347154 135922 347210 135978
rect 347278 135922 347334 135978
rect 347402 135922 347458 135978
rect 347526 135922 347582 135978
rect 347154 118294 347210 118350
rect 347278 118294 347334 118350
rect 347402 118294 347458 118350
rect 347526 118294 347582 118350
rect 347154 118170 347210 118226
rect 347278 118170 347334 118226
rect 347402 118170 347458 118226
rect 347526 118170 347582 118226
rect 347154 118046 347210 118102
rect 347278 118046 347334 118102
rect 347402 118046 347458 118102
rect 347526 118046 347582 118102
rect 347154 117922 347210 117978
rect 347278 117922 347334 117978
rect 347402 117922 347458 117978
rect 347526 117922 347582 117978
rect 347154 100294 347210 100350
rect 347278 100294 347334 100350
rect 347402 100294 347458 100350
rect 347526 100294 347582 100350
rect 347154 100170 347210 100226
rect 347278 100170 347334 100226
rect 347402 100170 347458 100226
rect 347526 100170 347582 100226
rect 347154 100046 347210 100102
rect 347278 100046 347334 100102
rect 347402 100046 347458 100102
rect 347526 100046 347582 100102
rect 347154 99922 347210 99978
rect 347278 99922 347334 99978
rect 347402 99922 347458 99978
rect 347526 99922 347582 99978
rect 347154 82294 347210 82350
rect 347278 82294 347334 82350
rect 347402 82294 347458 82350
rect 347526 82294 347582 82350
rect 347154 82170 347210 82226
rect 347278 82170 347334 82226
rect 347402 82170 347458 82226
rect 347526 82170 347582 82226
rect 347154 82046 347210 82102
rect 347278 82046 347334 82102
rect 347402 82046 347458 82102
rect 347526 82046 347582 82102
rect 347154 81922 347210 81978
rect 347278 81922 347334 81978
rect 347402 81922 347458 81978
rect 347526 81922 347582 81978
rect 347154 64294 347210 64350
rect 347278 64294 347334 64350
rect 347402 64294 347458 64350
rect 347526 64294 347582 64350
rect 347154 64170 347210 64226
rect 347278 64170 347334 64226
rect 347402 64170 347458 64226
rect 347526 64170 347582 64226
rect 347154 64046 347210 64102
rect 347278 64046 347334 64102
rect 347402 64046 347458 64102
rect 347526 64046 347582 64102
rect 347154 63922 347210 63978
rect 347278 63922 347334 63978
rect 347402 63922 347458 63978
rect 347526 63922 347582 63978
rect 347154 46294 347210 46350
rect 347278 46294 347334 46350
rect 347402 46294 347458 46350
rect 347526 46294 347582 46350
rect 347154 46170 347210 46226
rect 347278 46170 347334 46226
rect 347402 46170 347458 46226
rect 347526 46170 347582 46226
rect 347154 46046 347210 46102
rect 347278 46046 347334 46102
rect 347402 46046 347458 46102
rect 347526 46046 347582 46102
rect 347154 45922 347210 45978
rect 347278 45922 347334 45978
rect 347402 45922 347458 45978
rect 347526 45922 347582 45978
rect 343434 40294 343490 40350
rect 343558 40294 343614 40350
rect 343682 40294 343738 40350
rect 343806 40294 343862 40350
rect 343434 40170 343490 40226
rect 343558 40170 343614 40226
rect 343682 40170 343738 40226
rect 343806 40170 343862 40226
rect 343434 40046 343490 40102
rect 343558 40046 343614 40102
rect 343682 40046 343738 40102
rect 343806 40046 343862 40102
rect 343434 39922 343490 39978
rect 343558 39922 343614 39978
rect 343682 39922 343738 39978
rect 343806 39922 343862 39978
rect 342748 30662 342804 30718
rect 339388 30482 339444 30538
rect 336028 17162 336084 17218
rect 343434 22294 343490 22350
rect 343558 22294 343614 22350
rect 343682 22294 343738 22350
rect 343806 22294 343862 22350
rect 343434 22170 343490 22226
rect 343558 22170 343614 22226
rect 343682 22170 343738 22226
rect 343806 22170 343862 22226
rect 343434 22046 343490 22102
rect 343558 22046 343614 22102
rect 343682 22046 343738 22102
rect 343806 22046 343862 22102
rect 343434 21922 343490 21978
rect 343558 21922 343614 21978
rect 343682 21922 343738 21978
rect 343806 21922 343862 21978
rect 343434 4294 343490 4350
rect 343558 4294 343614 4350
rect 343682 4294 343738 4350
rect 343806 4294 343862 4350
rect 343434 4170 343490 4226
rect 343558 4170 343614 4226
rect 343682 4170 343738 4226
rect 343806 4170 343862 4226
rect 316434 -1176 316490 -1120
rect 316558 -1176 316614 -1120
rect 316682 -1176 316738 -1120
rect 316806 -1176 316862 -1120
rect 316434 -1300 316490 -1244
rect 316558 -1300 316614 -1244
rect 316682 -1300 316738 -1244
rect 316806 -1300 316862 -1244
rect 316434 -1424 316490 -1368
rect 316558 -1424 316614 -1368
rect 316682 -1424 316738 -1368
rect 316806 -1424 316862 -1368
rect 316434 -1548 316490 -1492
rect 316558 -1548 316614 -1492
rect 316682 -1548 316738 -1492
rect 316806 -1548 316862 -1492
rect 346108 42722 346164 42778
rect 374154 597156 374210 597212
rect 374278 597156 374334 597212
rect 374402 597156 374458 597212
rect 374526 597156 374582 597212
rect 374154 597032 374210 597088
rect 374278 597032 374334 597088
rect 374402 597032 374458 597088
rect 374526 597032 374582 597088
rect 374154 596908 374210 596964
rect 374278 596908 374334 596964
rect 374402 596908 374458 596964
rect 374526 596908 374582 596964
rect 374154 596784 374210 596840
rect 374278 596784 374334 596840
rect 374402 596784 374458 596840
rect 374526 596784 374582 596840
rect 374154 580294 374210 580350
rect 374278 580294 374334 580350
rect 374402 580294 374458 580350
rect 374526 580294 374582 580350
rect 374154 580170 374210 580226
rect 374278 580170 374334 580226
rect 374402 580170 374458 580226
rect 374526 580170 374582 580226
rect 374154 580046 374210 580102
rect 374278 580046 374334 580102
rect 374402 580046 374458 580102
rect 374526 580046 374582 580102
rect 374154 579922 374210 579978
rect 374278 579922 374334 579978
rect 374402 579922 374458 579978
rect 374526 579922 374582 579978
rect 374154 562294 374210 562350
rect 374278 562294 374334 562350
rect 374402 562294 374458 562350
rect 374526 562294 374582 562350
rect 374154 562170 374210 562226
rect 374278 562170 374334 562226
rect 374402 562170 374458 562226
rect 374526 562170 374582 562226
rect 374154 562046 374210 562102
rect 374278 562046 374334 562102
rect 374402 562046 374458 562102
rect 374526 562046 374582 562102
rect 374154 561922 374210 561978
rect 374278 561922 374334 561978
rect 374402 561922 374458 561978
rect 374526 561922 374582 561978
rect 374154 544294 374210 544350
rect 374278 544294 374334 544350
rect 374402 544294 374458 544350
rect 374526 544294 374582 544350
rect 374154 544170 374210 544226
rect 374278 544170 374334 544226
rect 374402 544170 374458 544226
rect 374526 544170 374582 544226
rect 374154 544046 374210 544102
rect 374278 544046 374334 544102
rect 374402 544046 374458 544102
rect 374526 544046 374582 544102
rect 374154 543922 374210 543978
rect 374278 543922 374334 543978
rect 374402 543922 374458 543978
rect 374526 543922 374582 543978
rect 374154 526294 374210 526350
rect 374278 526294 374334 526350
rect 374402 526294 374458 526350
rect 374526 526294 374582 526350
rect 374154 526170 374210 526226
rect 374278 526170 374334 526226
rect 374402 526170 374458 526226
rect 374526 526170 374582 526226
rect 374154 526046 374210 526102
rect 374278 526046 374334 526102
rect 374402 526046 374458 526102
rect 374526 526046 374582 526102
rect 374154 525922 374210 525978
rect 374278 525922 374334 525978
rect 374402 525922 374458 525978
rect 374526 525922 374582 525978
rect 374154 508294 374210 508350
rect 374278 508294 374334 508350
rect 374402 508294 374458 508350
rect 374526 508294 374582 508350
rect 374154 508170 374210 508226
rect 374278 508170 374334 508226
rect 374402 508170 374458 508226
rect 374526 508170 374582 508226
rect 374154 508046 374210 508102
rect 374278 508046 374334 508102
rect 374402 508046 374458 508102
rect 374526 508046 374582 508102
rect 374154 507922 374210 507978
rect 374278 507922 374334 507978
rect 374402 507922 374458 507978
rect 374526 507922 374582 507978
rect 374154 490294 374210 490350
rect 374278 490294 374334 490350
rect 374402 490294 374458 490350
rect 374526 490294 374582 490350
rect 374154 490170 374210 490226
rect 374278 490170 374334 490226
rect 374402 490170 374458 490226
rect 374526 490170 374582 490226
rect 374154 490046 374210 490102
rect 374278 490046 374334 490102
rect 374402 490046 374458 490102
rect 374526 490046 374582 490102
rect 374154 489922 374210 489978
rect 374278 489922 374334 489978
rect 374402 489922 374458 489978
rect 374526 489922 374582 489978
rect 374154 472294 374210 472350
rect 374278 472294 374334 472350
rect 374402 472294 374458 472350
rect 374526 472294 374582 472350
rect 374154 472170 374210 472226
rect 374278 472170 374334 472226
rect 374402 472170 374458 472226
rect 374526 472170 374582 472226
rect 374154 472046 374210 472102
rect 374278 472046 374334 472102
rect 374402 472046 374458 472102
rect 374526 472046 374582 472102
rect 374154 471922 374210 471978
rect 374278 471922 374334 471978
rect 374402 471922 374458 471978
rect 374526 471922 374582 471978
rect 374154 454294 374210 454350
rect 374278 454294 374334 454350
rect 374402 454294 374458 454350
rect 374526 454294 374582 454350
rect 374154 454170 374210 454226
rect 374278 454170 374334 454226
rect 374402 454170 374458 454226
rect 374526 454170 374582 454226
rect 374154 454046 374210 454102
rect 374278 454046 374334 454102
rect 374402 454046 374458 454102
rect 374526 454046 374582 454102
rect 374154 453922 374210 453978
rect 374278 453922 374334 453978
rect 374402 453922 374458 453978
rect 374526 453922 374582 453978
rect 374154 436294 374210 436350
rect 374278 436294 374334 436350
rect 374402 436294 374458 436350
rect 374526 436294 374582 436350
rect 374154 436170 374210 436226
rect 374278 436170 374334 436226
rect 374402 436170 374458 436226
rect 374526 436170 374582 436226
rect 374154 436046 374210 436102
rect 374278 436046 374334 436102
rect 374402 436046 374458 436102
rect 374526 436046 374582 436102
rect 374154 435922 374210 435978
rect 374278 435922 374334 435978
rect 374402 435922 374458 435978
rect 374526 435922 374582 435978
rect 374154 418294 374210 418350
rect 374278 418294 374334 418350
rect 374402 418294 374458 418350
rect 374526 418294 374582 418350
rect 374154 418170 374210 418226
rect 374278 418170 374334 418226
rect 374402 418170 374458 418226
rect 374526 418170 374582 418226
rect 374154 418046 374210 418102
rect 374278 418046 374334 418102
rect 374402 418046 374458 418102
rect 374526 418046 374582 418102
rect 374154 417922 374210 417978
rect 374278 417922 374334 417978
rect 374402 417922 374458 417978
rect 374526 417922 374582 417978
rect 374154 400294 374210 400350
rect 374278 400294 374334 400350
rect 374402 400294 374458 400350
rect 374526 400294 374582 400350
rect 374154 400170 374210 400226
rect 374278 400170 374334 400226
rect 374402 400170 374458 400226
rect 374526 400170 374582 400226
rect 374154 400046 374210 400102
rect 374278 400046 374334 400102
rect 374402 400046 374458 400102
rect 374526 400046 374582 400102
rect 374154 399922 374210 399978
rect 374278 399922 374334 399978
rect 374402 399922 374458 399978
rect 374526 399922 374582 399978
rect 374154 382294 374210 382350
rect 374278 382294 374334 382350
rect 374402 382294 374458 382350
rect 374526 382294 374582 382350
rect 374154 382170 374210 382226
rect 374278 382170 374334 382226
rect 374402 382170 374458 382226
rect 374526 382170 374582 382226
rect 374154 382046 374210 382102
rect 374278 382046 374334 382102
rect 374402 382046 374458 382102
rect 374526 382046 374582 382102
rect 374154 381922 374210 381978
rect 374278 381922 374334 381978
rect 374402 381922 374458 381978
rect 374526 381922 374582 381978
rect 374154 364294 374210 364350
rect 374278 364294 374334 364350
rect 374402 364294 374458 364350
rect 374526 364294 374582 364350
rect 374154 364170 374210 364226
rect 374278 364170 374334 364226
rect 374402 364170 374458 364226
rect 374526 364170 374582 364226
rect 374154 364046 374210 364102
rect 374278 364046 374334 364102
rect 374402 364046 374458 364102
rect 374526 364046 374582 364102
rect 374154 363922 374210 363978
rect 374278 363922 374334 363978
rect 374402 363922 374458 363978
rect 374526 363922 374582 363978
rect 374154 346294 374210 346350
rect 374278 346294 374334 346350
rect 374402 346294 374458 346350
rect 374526 346294 374582 346350
rect 374154 346170 374210 346226
rect 374278 346170 374334 346226
rect 374402 346170 374458 346226
rect 374526 346170 374582 346226
rect 374154 346046 374210 346102
rect 374278 346046 374334 346102
rect 374402 346046 374458 346102
rect 374526 346046 374582 346102
rect 374154 345922 374210 345978
rect 374278 345922 374334 345978
rect 374402 345922 374458 345978
rect 374526 345922 374582 345978
rect 374154 328294 374210 328350
rect 374278 328294 374334 328350
rect 374402 328294 374458 328350
rect 374526 328294 374582 328350
rect 374154 328170 374210 328226
rect 374278 328170 374334 328226
rect 374402 328170 374458 328226
rect 374526 328170 374582 328226
rect 374154 328046 374210 328102
rect 374278 328046 374334 328102
rect 374402 328046 374458 328102
rect 374526 328046 374582 328102
rect 374154 327922 374210 327978
rect 374278 327922 374334 327978
rect 374402 327922 374458 327978
rect 374526 327922 374582 327978
rect 374154 310294 374210 310350
rect 374278 310294 374334 310350
rect 374402 310294 374458 310350
rect 374526 310294 374582 310350
rect 374154 310170 374210 310226
rect 374278 310170 374334 310226
rect 374402 310170 374458 310226
rect 374526 310170 374582 310226
rect 374154 310046 374210 310102
rect 374278 310046 374334 310102
rect 374402 310046 374458 310102
rect 374526 310046 374582 310102
rect 374154 309922 374210 309978
rect 374278 309922 374334 309978
rect 374402 309922 374458 309978
rect 374526 309922 374582 309978
rect 374154 292294 374210 292350
rect 374278 292294 374334 292350
rect 374402 292294 374458 292350
rect 374526 292294 374582 292350
rect 374154 292170 374210 292226
rect 374278 292170 374334 292226
rect 374402 292170 374458 292226
rect 374526 292170 374582 292226
rect 374154 292046 374210 292102
rect 374278 292046 374334 292102
rect 374402 292046 374458 292102
rect 374526 292046 374582 292102
rect 374154 291922 374210 291978
rect 374278 291922 374334 291978
rect 374402 291922 374458 291978
rect 374526 291922 374582 291978
rect 374154 274294 374210 274350
rect 374278 274294 374334 274350
rect 374402 274294 374458 274350
rect 374526 274294 374582 274350
rect 374154 274170 374210 274226
rect 374278 274170 374334 274226
rect 374402 274170 374458 274226
rect 374526 274170 374582 274226
rect 374154 274046 374210 274102
rect 374278 274046 374334 274102
rect 374402 274046 374458 274102
rect 374526 274046 374582 274102
rect 374154 273922 374210 273978
rect 374278 273922 374334 273978
rect 374402 273922 374458 273978
rect 374526 273922 374582 273978
rect 374154 256294 374210 256350
rect 374278 256294 374334 256350
rect 374402 256294 374458 256350
rect 374526 256294 374582 256350
rect 374154 256170 374210 256226
rect 374278 256170 374334 256226
rect 374402 256170 374458 256226
rect 374526 256170 374582 256226
rect 374154 256046 374210 256102
rect 374278 256046 374334 256102
rect 374402 256046 374458 256102
rect 374526 256046 374582 256102
rect 374154 255922 374210 255978
rect 374278 255922 374334 255978
rect 374402 255922 374458 255978
rect 374526 255922 374582 255978
rect 374154 238294 374210 238350
rect 374278 238294 374334 238350
rect 374402 238294 374458 238350
rect 374526 238294 374582 238350
rect 374154 238170 374210 238226
rect 374278 238170 374334 238226
rect 374402 238170 374458 238226
rect 374526 238170 374582 238226
rect 374154 238046 374210 238102
rect 374278 238046 374334 238102
rect 374402 238046 374458 238102
rect 374526 238046 374582 238102
rect 374154 237922 374210 237978
rect 374278 237922 374334 237978
rect 374402 237922 374458 237978
rect 374526 237922 374582 237978
rect 374154 220294 374210 220350
rect 374278 220294 374334 220350
rect 374402 220294 374458 220350
rect 374526 220294 374582 220350
rect 374154 220170 374210 220226
rect 374278 220170 374334 220226
rect 374402 220170 374458 220226
rect 374526 220170 374582 220226
rect 374154 220046 374210 220102
rect 374278 220046 374334 220102
rect 374402 220046 374458 220102
rect 374526 220046 374582 220102
rect 374154 219922 374210 219978
rect 374278 219922 374334 219978
rect 374402 219922 374458 219978
rect 374526 219922 374582 219978
rect 374154 202294 374210 202350
rect 374278 202294 374334 202350
rect 374402 202294 374458 202350
rect 374526 202294 374582 202350
rect 374154 202170 374210 202226
rect 374278 202170 374334 202226
rect 374402 202170 374458 202226
rect 374526 202170 374582 202226
rect 374154 202046 374210 202102
rect 374278 202046 374334 202102
rect 374402 202046 374458 202102
rect 374526 202046 374582 202102
rect 374154 201922 374210 201978
rect 374278 201922 374334 201978
rect 374402 201922 374458 201978
rect 374526 201922 374582 201978
rect 374154 184294 374210 184350
rect 374278 184294 374334 184350
rect 374402 184294 374458 184350
rect 374526 184294 374582 184350
rect 374154 184170 374210 184226
rect 374278 184170 374334 184226
rect 374402 184170 374458 184226
rect 374526 184170 374582 184226
rect 374154 184046 374210 184102
rect 374278 184046 374334 184102
rect 374402 184046 374458 184102
rect 374526 184046 374582 184102
rect 374154 183922 374210 183978
rect 374278 183922 374334 183978
rect 374402 183922 374458 183978
rect 374526 183922 374582 183978
rect 374154 166294 374210 166350
rect 374278 166294 374334 166350
rect 374402 166294 374458 166350
rect 374526 166294 374582 166350
rect 374154 166170 374210 166226
rect 374278 166170 374334 166226
rect 374402 166170 374458 166226
rect 374526 166170 374582 166226
rect 374154 166046 374210 166102
rect 374278 166046 374334 166102
rect 374402 166046 374458 166102
rect 374526 166046 374582 166102
rect 374154 165922 374210 165978
rect 374278 165922 374334 165978
rect 374402 165922 374458 165978
rect 374526 165922 374582 165978
rect 374154 148294 374210 148350
rect 374278 148294 374334 148350
rect 374402 148294 374458 148350
rect 374526 148294 374582 148350
rect 374154 148170 374210 148226
rect 374278 148170 374334 148226
rect 374402 148170 374458 148226
rect 374526 148170 374582 148226
rect 374154 148046 374210 148102
rect 374278 148046 374334 148102
rect 374402 148046 374458 148102
rect 374526 148046 374582 148102
rect 374154 147922 374210 147978
rect 374278 147922 374334 147978
rect 374402 147922 374458 147978
rect 374526 147922 374582 147978
rect 374154 130294 374210 130350
rect 374278 130294 374334 130350
rect 374402 130294 374458 130350
rect 374526 130294 374582 130350
rect 374154 130170 374210 130226
rect 374278 130170 374334 130226
rect 374402 130170 374458 130226
rect 374526 130170 374582 130226
rect 374154 130046 374210 130102
rect 374278 130046 374334 130102
rect 374402 130046 374458 130102
rect 374526 130046 374582 130102
rect 374154 129922 374210 129978
rect 374278 129922 374334 129978
rect 374402 129922 374458 129978
rect 374526 129922 374582 129978
rect 374154 112294 374210 112350
rect 374278 112294 374334 112350
rect 374402 112294 374458 112350
rect 374526 112294 374582 112350
rect 374154 112170 374210 112226
rect 374278 112170 374334 112226
rect 374402 112170 374458 112226
rect 374526 112170 374582 112226
rect 374154 112046 374210 112102
rect 374278 112046 374334 112102
rect 374402 112046 374458 112102
rect 374526 112046 374582 112102
rect 374154 111922 374210 111978
rect 374278 111922 374334 111978
rect 374402 111922 374458 111978
rect 374526 111922 374582 111978
rect 374154 94294 374210 94350
rect 374278 94294 374334 94350
rect 374402 94294 374458 94350
rect 374526 94294 374582 94350
rect 374154 94170 374210 94226
rect 374278 94170 374334 94226
rect 374402 94170 374458 94226
rect 374526 94170 374582 94226
rect 374154 94046 374210 94102
rect 374278 94046 374334 94102
rect 374402 94046 374458 94102
rect 374526 94046 374582 94102
rect 374154 93922 374210 93978
rect 374278 93922 374334 93978
rect 374402 93922 374458 93978
rect 374526 93922 374582 93978
rect 374154 76294 374210 76350
rect 374278 76294 374334 76350
rect 374402 76294 374458 76350
rect 374526 76294 374582 76350
rect 374154 76170 374210 76226
rect 374278 76170 374334 76226
rect 374402 76170 374458 76226
rect 374526 76170 374582 76226
rect 374154 76046 374210 76102
rect 374278 76046 374334 76102
rect 374402 76046 374458 76102
rect 374526 76046 374582 76102
rect 374154 75922 374210 75978
rect 374278 75922 374334 75978
rect 374402 75922 374458 75978
rect 374526 75922 374582 75978
rect 374154 58294 374210 58350
rect 374278 58294 374334 58350
rect 374402 58294 374458 58350
rect 374526 58294 374582 58350
rect 374154 58170 374210 58226
rect 374278 58170 374334 58226
rect 374402 58170 374458 58226
rect 374526 58170 374582 58226
rect 374154 58046 374210 58102
rect 374278 58046 374334 58102
rect 374402 58046 374458 58102
rect 374526 58046 374582 58102
rect 374154 57922 374210 57978
rect 374278 57922 374334 57978
rect 374402 57922 374458 57978
rect 374526 57922 374582 57978
rect 364588 44162 364644 44218
rect 352828 43982 352884 44038
rect 347154 28294 347210 28350
rect 347278 28294 347334 28350
rect 347402 28294 347458 28350
rect 347526 28294 347582 28350
rect 347154 28170 347210 28226
rect 347278 28170 347334 28226
rect 347402 28170 347458 28226
rect 347526 28170 347582 28226
rect 347154 28046 347210 28102
rect 347278 28046 347334 28102
rect 347402 28046 347458 28102
rect 347526 28046 347582 28102
rect 347154 27922 347210 27978
rect 347278 27922 347334 27978
rect 347402 27922 347458 27978
rect 347526 27922 347582 27978
rect 351148 43802 351204 43858
rect 347154 10294 347210 10350
rect 347278 10294 347334 10350
rect 347402 10294 347458 10350
rect 347526 10294 347582 10350
rect 347154 10170 347210 10226
rect 347278 10170 347334 10226
rect 347402 10170 347458 10226
rect 347526 10170 347582 10226
rect 347154 10046 347210 10102
rect 347278 10046 347334 10102
rect 347402 10046 347458 10102
rect 347526 10046 347582 10102
rect 347154 9922 347210 9978
rect 347278 9922 347334 9978
rect 347402 9922 347458 9978
rect 347526 9922 347582 9978
rect 343434 4046 343490 4102
rect 343558 4046 343614 4102
rect 343682 4046 343738 4102
rect 343806 4046 343862 4102
rect 343434 3922 343490 3978
rect 343558 3922 343614 3978
rect 343682 3922 343738 3978
rect 343806 3922 343862 3978
rect 343434 -216 343490 -160
rect 343558 -216 343614 -160
rect 343682 -216 343738 -160
rect 343806 -216 343862 -160
rect 343434 -340 343490 -284
rect 343558 -340 343614 -284
rect 343682 -340 343738 -284
rect 343806 -340 343862 -284
rect 343434 -464 343490 -408
rect 343558 -464 343614 -408
rect 343682 -464 343738 -408
rect 343806 -464 343862 -408
rect 343434 -588 343490 -532
rect 343558 -588 343614 -532
rect 343682 -588 343738 -532
rect 343806 -588 343862 -532
rect 347788 24002 347844 24058
rect 362908 42182 362964 42238
rect 359548 20222 359604 20278
rect 377874 598116 377930 598172
rect 377998 598116 378054 598172
rect 378122 598116 378178 598172
rect 378246 598116 378302 598172
rect 377874 597992 377930 598048
rect 377998 597992 378054 598048
rect 378122 597992 378178 598048
rect 378246 597992 378302 598048
rect 377874 597868 377930 597924
rect 377998 597868 378054 597924
rect 378122 597868 378178 597924
rect 378246 597868 378302 597924
rect 377874 597744 377930 597800
rect 377998 597744 378054 597800
rect 378122 597744 378178 597800
rect 378246 597744 378302 597800
rect 377874 586294 377930 586350
rect 377998 586294 378054 586350
rect 378122 586294 378178 586350
rect 378246 586294 378302 586350
rect 377874 586170 377930 586226
rect 377998 586170 378054 586226
rect 378122 586170 378178 586226
rect 378246 586170 378302 586226
rect 377874 586046 377930 586102
rect 377998 586046 378054 586102
rect 378122 586046 378178 586102
rect 378246 586046 378302 586102
rect 377874 585922 377930 585978
rect 377998 585922 378054 585978
rect 378122 585922 378178 585978
rect 378246 585922 378302 585978
rect 377874 568294 377930 568350
rect 377998 568294 378054 568350
rect 378122 568294 378178 568350
rect 378246 568294 378302 568350
rect 377874 568170 377930 568226
rect 377998 568170 378054 568226
rect 378122 568170 378178 568226
rect 378246 568170 378302 568226
rect 377874 568046 377930 568102
rect 377998 568046 378054 568102
rect 378122 568046 378178 568102
rect 378246 568046 378302 568102
rect 377874 567922 377930 567978
rect 377998 567922 378054 567978
rect 378122 567922 378178 567978
rect 378246 567922 378302 567978
rect 377874 550294 377930 550350
rect 377998 550294 378054 550350
rect 378122 550294 378178 550350
rect 378246 550294 378302 550350
rect 377874 550170 377930 550226
rect 377998 550170 378054 550226
rect 378122 550170 378178 550226
rect 378246 550170 378302 550226
rect 377874 550046 377930 550102
rect 377998 550046 378054 550102
rect 378122 550046 378178 550102
rect 378246 550046 378302 550102
rect 377874 549922 377930 549978
rect 377998 549922 378054 549978
rect 378122 549922 378178 549978
rect 378246 549922 378302 549978
rect 377874 532294 377930 532350
rect 377998 532294 378054 532350
rect 378122 532294 378178 532350
rect 378246 532294 378302 532350
rect 377874 532170 377930 532226
rect 377998 532170 378054 532226
rect 378122 532170 378178 532226
rect 378246 532170 378302 532226
rect 377874 532046 377930 532102
rect 377998 532046 378054 532102
rect 378122 532046 378178 532102
rect 378246 532046 378302 532102
rect 377874 531922 377930 531978
rect 377998 531922 378054 531978
rect 378122 531922 378178 531978
rect 378246 531922 378302 531978
rect 377874 514294 377930 514350
rect 377998 514294 378054 514350
rect 378122 514294 378178 514350
rect 378246 514294 378302 514350
rect 377874 514170 377930 514226
rect 377998 514170 378054 514226
rect 378122 514170 378178 514226
rect 378246 514170 378302 514226
rect 377874 514046 377930 514102
rect 377998 514046 378054 514102
rect 378122 514046 378178 514102
rect 378246 514046 378302 514102
rect 377874 513922 377930 513978
rect 377998 513922 378054 513978
rect 378122 513922 378178 513978
rect 378246 513922 378302 513978
rect 377874 496294 377930 496350
rect 377998 496294 378054 496350
rect 378122 496294 378178 496350
rect 378246 496294 378302 496350
rect 377874 496170 377930 496226
rect 377998 496170 378054 496226
rect 378122 496170 378178 496226
rect 378246 496170 378302 496226
rect 377874 496046 377930 496102
rect 377998 496046 378054 496102
rect 378122 496046 378178 496102
rect 378246 496046 378302 496102
rect 377874 495922 377930 495978
rect 377998 495922 378054 495978
rect 378122 495922 378178 495978
rect 378246 495922 378302 495978
rect 377874 478294 377930 478350
rect 377998 478294 378054 478350
rect 378122 478294 378178 478350
rect 378246 478294 378302 478350
rect 377874 478170 377930 478226
rect 377998 478170 378054 478226
rect 378122 478170 378178 478226
rect 378246 478170 378302 478226
rect 377874 478046 377930 478102
rect 377998 478046 378054 478102
rect 378122 478046 378178 478102
rect 378246 478046 378302 478102
rect 377874 477922 377930 477978
rect 377998 477922 378054 477978
rect 378122 477922 378178 477978
rect 378246 477922 378302 477978
rect 377874 460294 377930 460350
rect 377998 460294 378054 460350
rect 378122 460294 378178 460350
rect 378246 460294 378302 460350
rect 377874 460170 377930 460226
rect 377998 460170 378054 460226
rect 378122 460170 378178 460226
rect 378246 460170 378302 460226
rect 377874 460046 377930 460102
rect 377998 460046 378054 460102
rect 378122 460046 378178 460102
rect 378246 460046 378302 460102
rect 377874 459922 377930 459978
rect 377998 459922 378054 459978
rect 378122 459922 378178 459978
rect 378246 459922 378302 459978
rect 377874 442294 377930 442350
rect 377998 442294 378054 442350
rect 378122 442294 378178 442350
rect 378246 442294 378302 442350
rect 377874 442170 377930 442226
rect 377998 442170 378054 442226
rect 378122 442170 378178 442226
rect 378246 442170 378302 442226
rect 377874 442046 377930 442102
rect 377998 442046 378054 442102
rect 378122 442046 378178 442102
rect 378246 442046 378302 442102
rect 377874 441922 377930 441978
rect 377998 441922 378054 441978
rect 378122 441922 378178 441978
rect 378246 441922 378302 441978
rect 377874 424294 377930 424350
rect 377998 424294 378054 424350
rect 378122 424294 378178 424350
rect 378246 424294 378302 424350
rect 377874 424170 377930 424226
rect 377998 424170 378054 424226
rect 378122 424170 378178 424226
rect 378246 424170 378302 424226
rect 377874 424046 377930 424102
rect 377998 424046 378054 424102
rect 378122 424046 378178 424102
rect 378246 424046 378302 424102
rect 377874 423922 377930 423978
rect 377998 423922 378054 423978
rect 378122 423922 378178 423978
rect 378246 423922 378302 423978
rect 377874 406294 377930 406350
rect 377998 406294 378054 406350
rect 378122 406294 378178 406350
rect 378246 406294 378302 406350
rect 377874 406170 377930 406226
rect 377998 406170 378054 406226
rect 378122 406170 378178 406226
rect 378246 406170 378302 406226
rect 377874 406046 377930 406102
rect 377998 406046 378054 406102
rect 378122 406046 378178 406102
rect 378246 406046 378302 406102
rect 377874 405922 377930 405978
rect 377998 405922 378054 405978
rect 378122 405922 378178 405978
rect 378246 405922 378302 405978
rect 377874 388294 377930 388350
rect 377998 388294 378054 388350
rect 378122 388294 378178 388350
rect 378246 388294 378302 388350
rect 377874 388170 377930 388226
rect 377998 388170 378054 388226
rect 378122 388170 378178 388226
rect 378246 388170 378302 388226
rect 377874 388046 377930 388102
rect 377998 388046 378054 388102
rect 378122 388046 378178 388102
rect 378246 388046 378302 388102
rect 377874 387922 377930 387978
rect 377998 387922 378054 387978
rect 378122 387922 378178 387978
rect 378246 387922 378302 387978
rect 377874 370294 377930 370350
rect 377998 370294 378054 370350
rect 378122 370294 378178 370350
rect 378246 370294 378302 370350
rect 377874 370170 377930 370226
rect 377998 370170 378054 370226
rect 378122 370170 378178 370226
rect 378246 370170 378302 370226
rect 377874 370046 377930 370102
rect 377998 370046 378054 370102
rect 378122 370046 378178 370102
rect 378246 370046 378302 370102
rect 377874 369922 377930 369978
rect 377998 369922 378054 369978
rect 378122 369922 378178 369978
rect 378246 369922 378302 369978
rect 377874 352294 377930 352350
rect 377998 352294 378054 352350
rect 378122 352294 378178 352350
rect 378246 352294 378302 352350
rect 377874 352170 377930 352226
rect 377998 352170 378054 352226
rect 378122 352170 378178 352226
rect 378246 352170 378302 352226
rect 377874 352046 377930 352102
rect 377998 352046 378054 352102
rect 378122 352046 378178 352102
rect 378246 352046 378302 352102
rect 377874 351922 377930 351978
rect 377998 351922 378054 351978
rect 378122 351922 378178 351978
rect 378246 351922 378302 351978
rect 377874 334294 377930 334350
rect 377998 334294 378054 334350
rect 378122 334294 378178 334350
rect 378246 334294 378302 334350
rect 377874 334170 377930 334226
rect 377998 334170 378054 334226
rect 378122 334170 378178 334226
rect 378246 334170 378302 334226
rect 377874 334046 377930 334102
rect 377998 334046 378054 334102
rect 378122 334046 378178 334102
rect 378246 334046 378302 334102
rect 377874 333922 377930 333978
rect 377998 333922 378054 333978
rect 378122 333922 378178 333978
rect 378246 333922 378302 333978
rect 377874 316294 377930 316350
rect 377998 316294 378054 316350
rect 378122 316294 378178 316350
rect 378246 316294 378302 316350
rect 377874 316170 377930 316226
rect 377998 316170 378054 316226
rect 378122 316170 378178 316226
rect 378246 316170 378302 316226
rect 377874 316046 377930 316102
rect 377998 316046 378054 316102
rect 378122 316046 378178 316102
rect 378246 316046 378302 316102
rect 377874 315922 377930 315978
rect 377998 315922 378054 315978
rect 378122 315922 378178 315978
rect 378246 315922 378302 315978
rect 377874 298294 377930 298350
rect 377998 298294 378054 298350
rect 378122 298294 378178 298350
rect 378246 298294 378302 298350
rect 377874 298170 377930 298226
rect 377998 298170 378054 298226
rect 378122 298170 378178 298226
rect 378246 298170 378302 298226
rect 377874 298046 377930 298102
rect 377998 298046 378054 298102
rect 378122 298046 378178 298102
rect 378246 298046 378302 298102
rect 377874 297922 377930 297978
rect 377998 297922 378054 297978
rect 378122 297922 378178 297978
rect 378246 297922 378302 297978
rect 377874 280294 377930 280350
rect 377998 280294 378054 280350
rect 378122 280294 378178 280350
rect 378246 280294 378302 280350
rect 377874 280170 377930 280226
rect 377998 280170 378054 280226
rect 378122 280170 378178 280226
rect 378246 280170 378302 280226
rect 377874 280046 377930 280102
rect 377998 280046 378054 280102
rect 378122 280046 378178 280102
rect 378246 280046 378302 280102
rect 377874 279922 377930 279978
rect 377998 279922 378054 279978
rect 378122 279922 378178 279978
rect 378246 279922 378302 279978
rect 377874 262294 377930 262350
rect 377998 262294 378054 262350
rect 378122 262294 378178 262350
rect 378246 262294 378302 262350
rect 377874 262170 377930 262226
rect 377998 262170 378054 262226
rect 378122 262170 378178 262226
rect 378246 262170 378302 262226
rect 377874 262046 377930 262102
rect 377998 262046 378054 262102
rect 378122 262046 378178 262102
rect 378246 262046 378302 262102
rect 377874 261922 377930 261978
rect 377998 261922 378054 261978
rect 378122 261922 378178 261978
rect 378246 261922 378302 261978
rect 377874 244294 377930 244350
rect 377998 244294 378054 244350
rect 378122 244294 378178 244350
rect 378246 244294 378302 244350
rect 377874 244170 377930 244226
rect 377998 244170 378054 244226
rect 378122 244170 378178 244226
rect 378246 244170 378302 244226
rect 377874 244046 377930 244102
rect 377998 244046 378054 244102
rect 378122 244046 378178 244102
rect 378246 244046 378302 244102
rect 377874 243922 377930 243978
rect 377998 243922 378054 243978
rect 378122 243922 378178 243978
rect 378246 243922 378302 243978
rect 377874 226294 377930 226350
rect 377998 226294 378054 226350
rect 378122 226294 378178 226350
rect 378246 226294 378302 226350
rect 377874 226170 377930 226226
rect 377998 226170 378054 226226
rect 378122 226170 378178 226226
rect 378246 226170 378302 226226
rect 377874 226046 377930 226102
rect 377998 226046 378054 226102
rect 378122 226046 378178 226102
rect 378246 226046 378302 226102
rect 377874 225922 377930 225978
rect 377998 225922 378054 225978
rect 378122 225922 378178 225978
rect 378246 225922 378302 225978
rect 377874 208294 377930 208350
rect 377998 208294 378054 208350
rect 378122 208294 378178 208350
rect 378246 208294 378302 208350
rect 377874 208170 377930 208226
rect 377998 208170 378054 208226
rect 378122 208170 378178 208226
rect 378246 208170 378302 208226
rect 377874 208046 377930 208102
rect 377998 208046 378054 208102
rect 378122 208046 378178 208102
rect 378246 208046 378302 208102
rect 377874 207922 377930 207978
rect 377998 207922 378054 207978
rect 378122 207922 378178 207978
rect 378246 207922 378302 207978
rect 377874 190294 377930 190350
rect 377998 190294 378054 190350
rect 378122 190294 378178 190350
rect 378246 190294 378302 190350
rect 377874 190170 377930 190226
rect 377998 190170 378054 190226
rect 378122 190170 378178 190226
rect 378246 190170 378302 190226
rect 377874 190046 377930 190102
rect 377998 190046 378054 190102
rect 378122 190046 378178 190102
rect 378246 190046 378302 190102
rect 377874 189922 377930 189978
rect 377998 189922 378054 189978
rect 378122 189922 378178 189978
rect 378246 189922 378302 189978
rect 377874 172294 377930 172350
rect 377998 172294 378054 172350
rect 378122 172294 378178 172350
rect 378246 172294 378302 172350
rect 377874 172170 377930 172226
rect 377998 172170 378054 172226
rect 378122 172170 378178 172226
rect 378246 172170 378302 172226
rect 377874 172046 377930 172102
rect 377998 172046 378054 172102
rect 378122 172046 378178 172102
rect 378246 172046 378302 172102
rect 377874 171922 377930 171978
rect 377998 171922 378054 171978
rect 378122 171922 378178 171978
rect 378246 171922 378302 171978
rect 377874 154294 377930 154350
rect 377998 154294 378054 154350
rect 378122 154294 378178 154350
rect 378246 154294 378302 154350
rect 377874 154170 377930 154226
rect 377998 154170 378054 154226
rect 378122 154170 378178 154226
rect 378246 154170 378302 154226
rect 377874 154046 377930 154102
rect 377998 154046 378054 154102
rect 378122 154046 378178 154102
rect 378246 154046 378302 154102
rect 377874 153922 377930 153978
rect 377998 153922 378054 153978
rect 378122 153922 378178 153978
rect 378246 153922 378302 153978
rect 377874 136294 377930 136350
rect 377998 136294 378054 136350
rect 378122 136294 378178 136350
rect 378246 136294 378302 136350
rect 377874 136170 377930 136226
rect 377998 136170 378054 136226
rect 378122 136170 378178 136226
rect 378246 136170 378302 136226
rect 377874 136046 377930 136102
rect 377998 136046 378054 136102
rect 378122 136046 378178 136102
rect 378246 136046 378302 136102
rect 377874 135922 377930 135978
rect 377998 135922 378054 135978
rect 378122 135922 378178 135978
rect 378246 135922 378302 135978
rect 377874 118294 377930 118350
rect 377998 118294 378054 118350
rect 378122 118294 378178 118350
rect 378246 118294 378302 118350
rect 377874 118170 377930 118226
rect 377998 118170 378054 118226
rect 378122 118170 378178 118226
rect 378246 118170 378302 118226
rect 377874 118046 377930 118102
rect 377998 118046 378054 118102
rect 378122 118046 378178 118102
rect 378246 118046 378302 118102
rect 377874 117922 377930 117978
rect 377998 117922 378054 117978
rect 378122 117922 378178 117978
rect 378246 117922 378302 117978
rect 377874 100294 377930 100350
rect 377998 100294 378054 100350
rect 378122 100294 378178 100350
rect 378246 100294 378302 100350
rect 377874 100170 377930 100226
rect 377998 100170 378054 100226
rect 378122 100170 378178 100226
rect 378246 100170 378302 100226
rect 377874 100046 377930 100102
rect 377998 100046 378054 100102
rect 378122 100046 378178 100102
rect 378246 100046 378302 100102
rect 377874 99922 377930 99978
rect 377998 99922 378054 99978
rect 378122 99922 378178 99978
rect 378246 99922 378302 99978
rect 377874 82294 377930 82350
rect 377998 82294 378054 82350
rect 378122 82294 378178 82350
rect 378246 82294 378302 82350
rect 377874 82170 377930 82226
rect 377998 82170 378054 82226
rect 378122 82170 378178 82226
rect 378246 82170 378302 82226
rect 377874 82046 377930 82102
rect 377998 82046 378054 82102
rect 378122 82046 378178 82102
rect 378246 82046 378302 82102
rect 377874 81922 377930 81978
rect 377998 81922 378054 81978
rect 378122 81922 378178 81978
rect 378246 81922 378302 81978
rect 404874 597156 404930 597212
rect 404998 597156 405054 597212
rect 405122 597156 405178 597212
rect 405246 597156 405302 597212
rect 404874 597032 404930 597088
rect 404998 597032 405054 597088
rect 405122 597032 405178 597088
rect 405246 597032 405302 597088
rect 404874 596908 404930 596964
rect 404998 596908 405054 596964
rect 405122 596908 405178 596964
rect 405246 596908 405302 596964
rect 404874 596784 404930 596840
rect 404998 596784 405054 596840
rect 405122 596784 405178 596840
rect 405246 596784 405302 596840
rect 404874 580294 404930 580350
rect 404998 580294 405054 580350
rect 405122 580294 405178 580350
rect 405246 580294 405302 580350
rect 404874 580170 404930 580226
rect 404998 580170 405054 580226
rect 405122 580170 405178 580226
rect 405246 580170 405302 580226
rect 404874 580046 404930 580102
rect 404998 580046 405054 580102
rect 405122 580046 405178 580102
rect 405246 580046 405302 580102
rect 404874 579922 404930 579978
rect 404998 579922 405054 579978
rect 405122 579922 405178 579978
rect 405246 579922 405302 579978
rect 404874 562294 404930 562350
rect 404998 562294 405054 562350
rect 405122 562294 405178 562350
rect 405246 562294 405302 562350
rect 404874 562170 404930 562226
rect 404998 562170 405054 562226
rect 405122 562170 405178 562226
rect 405246 562170 405302 562226
rect 404874 562046 404930 562102
rect 404998 562046 405054 562102
rect 405122 562046 405178 562102
rect 405246 562046 405302 562102
rect 404874 561922 404930 561978
rect 404998 561922 405054 561978
rect 405122 561922 405178 561978
rect 405246 561922 405302 561978
rect 404874 544294 404930 544350
rect 404998 544294 405054 544350
rect 405122 544294 405178 544350
rect 405246 544294 405302 544350
rect 404874 544170 404930 544226
rect 404998 544170 405054 544226
rect 405122 544170 405178 544226
rect 405246 544170 405302 544226
rect 404874 544046 404930 544102
rect 404998 544046 405054 544102
rect 405122 544046 405178 544102
rect 405246 544046 405302 544102
rect 404874 543922 404930 543978
rect 404998 543922 405054 543978
rect 405122 543922 405178 543978
rect 405246 543922 405302 543978
rect 404874 526294 404930 526350
rect 404998 526294 405054 526350
rect 405122 526294 405178 526350
rect 405246 526294 405302 526350
rect 404874 526170 404930 526226
rect 404998 526170 405054 526226
rect 405122 526170 405178 526226
rect 405246 526170 405302 526226
rect 404874 526046 404930 526102
rect 404998 526046 405054 526102
rect 405122 526046 405178 526102
rect 405246 526046 405302 526102
rect 404874 525922 404930 525978
rect 404998 525922 405054 525978
rect 405122 525922 405178 525978
rect 405246 525922 405302 525978
rect 404874 508294 404930 508350
rect 404998 508294 405054 508350
rect 405122 508294 405178 508350
rect 405246 508294 405302 508350
rect 404874 508170 404930 508226
rect 404998 508170 405054 508226
rect 405122 508170 405178 508226
rect 405246 508170 405302 508226
rect 404874 508046 404930 508102
rect 404998 508046 405054 508102
rect 405122 508046 405178 508102
rect 405246 508046 405302 508102
rect 404874 507922 404930 507978
rect 404998 507922 405054 507978
rect 405122 507922 405178 507978
rect 405246 507922 405302 507978
rect 404874 490294 404930 490350
rect 404998 490294 405054 490350
rect 405122 490294 405178 490350
rect 405246 490294 405302 490350
rect 404874 490170 404930 490226
rect 404998 490170 405054 490226
rect 405122 490170 405178 490226
rect 405246 490170 405302 490226
rect 404874 490046 404930 490102
rect 404998 490046 405054 490102
rect 405122 490046 405178 490102
rect 405246 490046 405302 490102
rect 404874 489922 404930 489978
rect 404998 489922 405054 489978
rect 405122 489922 405178 489978
rect 405246 489922 405302 489978
rect 404874 472294 404930 472350
rect 404998 472294 405054 472350
rect 405122 472294 405178 472350
rect 405246 472294 405302 472350
rect 404874 472170 404930 472226
rect 404998 472170 405054 472226
rect 405122 472170 405178 472226
rect 405246 472170 405302 472226
rect 404874 472046 404930 472102
rect 404998 472046 405054 472102
rect 405122 472046 405178 472102
rect 405246 472046 405302 472102
rect 404874 471922 404930 471978
rect 404998 471922 405054 471978
rect 405122 471922 405178 471978
rect 405246 471922 405302 471978
rect 404874 454294 404930 454350
rect 404998 454294 405054 454350
rect 405122 454294 405178 454350
rect 405246 454294 405302 454350
rect 404874 454170 404930 454226
rect 404998 454170 405054 454226
rect 405122 454170 405178 454226
rect 405246 454170 405302 454226
rect 404874 454046 404930 454102
rect 404998 454046 405054 454102
rect 405122 454046 405178 454102
rect 405246 454046 405302 454102
rect 404874 453922 404930 453978
rect 404998 453922 405054 453978
rect 405122 453922 405178 453978
rect 405246 453922 405302 453978
rect 404874 436294 404930 436350
rect 404998 436294 405054 436350
rect 405122 436294 405178 436350
rect 405246 436294 405302 436350
rect 404874 436170 404930 436226
rect 404998 436170 405054 436226
rect 405122 436170 405178 436226
rect 405246 436170 405302 436226
rect 404874 436046 404930 436102
rect 404998 436046 405054 436102
rect 405122 436046 405178 436102
rect 405246 436046 405302 436102
rect 404874 435922 404930 435978
rect 404998 435922 405054 435978
rect 405122 435922 405178 435978
rect 405246 435922 405302 435978
rect 404874 418294 404930 418350
rect 404998 418294 405054 418350
rect 405122 418294 405178 418350
rect 405246 418294 405302 418350
rect 404874 418170 404930 418226
rect 404998 418170 405054 418226
rect 405122 418170 405178 418226
rect 405246 418170 405302 418226
rect 404874 418046 404930 418102
rect 404998 418046 405054 418102
rect 405122 418046 405178 418102
rect 405246 418046 405302 418102
rect 404874 417922 404930 417978
rect 404998 417922 405054 417978
rect 405122 417922 405178 417978
rect 405246 417922 405302 417978
rect 404874 400294 404930 400350
rect 404998 400294 405054 400350
rect 405122 400294 405178 400350
rect 405246 400294 405302 400350
rect 404874 400170 404930 400226
rect 404998 400170 405054 400226
rect 405122 400170 405178 400226
rect 405246 400170 405302 400226
rect 404874 400046 404930 400102
rect 404998 400046 405054 400102
rect 405122 400046 405178 400102
rect 405246 400046 405302 400102
rect 404874 399922 404930 399978
rect 404998 399922 405054 399978
rect 405122 399922 405178 399978
rect 405246 399922 405302 399978
rect 404874 382294 404930 382350
rect 404998 382294 405054 382350
rect 405122 382294 405178 382350
rect 405246 382294 405302 382350
rect 404874 382170 404930 382226
rect 404998 382170 405054 382226
rect 405122 382170 405178 382226
rect 405246 382170 405302 382226
rect 404874 382046 404930 382102
rect 404998 382046 405054 382102
rect 405122 382046 405178 382102
rect 405246 382046 405302 382102
rect 404874 381922 404930 381978
rect 404998 381922 405054 381978
rect 405122 381922 405178 381978
rect 405246 381922 405302 381978
rect 404874 364294 404930 364350
rect 404998 364294 405054 364350
rect 405122 364294 405178 364350
rect 405246 364294 405302 364350
rect 404874 364170 404930 364226
rect 404998 364170 405054 364226
rect 405122 364170 405178 364226
rect 405246 364170 405302 364226
rect 404874 364046 404930 364102
rect 404998 364046 405054 364102
rect 405122 364046 405178 364102
rect 405246 364046 405302 364102
rect 404874 363922 404930 363978
rect 404998 363922 405054 363978
rect 405122 363922 405178 363978
rect 405246 363922 405302 363978
rect 404874 346294 404930 346350
rect 404998 346294 405054 346350
rect 405122 346294 405178 346350
rect 405246 346294 405302 346350
rect 404874 346170 404930 346226
rect 404998 346170 405054 346226
rect 405122 346170 405178 346226
rect 405246 346170 405302 346226
rect 404874 346046 404930 346102
rect 404998 346046 405054 346102
rect 405122 346046 405178 346102
rect 405246 346046 405302 346102
rect 404874 345922 404930 345978
rect 404998 345922 405054 345978
rect 405122 345922 405178 345978
rect 405246 345922 405302 345978
rect 404874 328294 404930 328350
rect 404998 328294 405054 328350
rect 405122 328294 405178 328350
rect 405246 328294 405302 328350
rect 404874 328170 404930 328226
rect 404998 328170 405054 328226
rect 405122 328170 405178 328226
rect 405246 328170 405302 328226
rect 404874 328046 404930 328102
rect 404998 328046 405054 328102
rect 405122 328046 405178 328102
rect 405246 328046 405302 328102
rect 404874 327922 404930 327978
rect 404998 327922 405054 327978
rect 405122 327922 405178 327978
rect 405246 327922 405302 327978
rect 404874 310294 404930 310350
rect 404998 310294 405054 310350
rect 405122 310294 405178 310350
rect 405246 310294 405302 310350
rect 404874 310170 404930 310226
rect 404998 310170 405054 310226
rect 405122 310170 405178 310226
rect 405246 310170 405302 310226
rect 404874 310046 404930 310102
rect 404998 310046 405054 310102
rect 405122 310046 405178 310102
rect 405246 310046 405302 310102
rect 404874 309922 404930 309978
rect 404998 309922 405054 309978
rect 405122 309922 405178 309978
rect 405246 309922 405302 309978
rect 404874 292294 404930 292350
rect 404998 292294 405054 292350
rect 405122 292294 405178 292350
rect 405246 292294 405302 292350
rect 404874 292170 404930 292226
rect 404998 292170 405054 292226
rect 405122 292170 405178 292226
rect 405246 292170 405302 292226
rect 404874 292046 404930 292102
rect 404998 292046 405054 292102
rect 405122 292046 405178 292102
rect 405246 292046 405302 292102
rect 404874 291922 404930 291978
rect 404998 291922 405054 291978
rect 405122 291922 405178 291978
rect 405246 291922 405302 291978
rect 404874 274294 404930 274350
rect 404998 274294 405054 274350
rect 405122 274294 405178 274350
rect 405246 274294 405302 274350
rect 404874 274170 404930 274226
rect 404998 274170 405054 274226
rect 405122 274170 405178 274226
rect 405246 274170 405302 274226
rect 404874 274046 404930 274102
rect 404998 274046 405054 274102
rect 405122 274046 405178 274102
rect 405246 274046 405302 274102
rect 404874 273922 404930 273978
rect 404998 273922 405054 273978
rect 405122 273922 405178 273978
rect 405246 273922 405302 273978
rect 404874 256294 404930 256350
rect 404998 256294 405054 256350
rect 405122 256294 405178 256350
rect 405246 256294 405302 256350
rect 404874 256170 404930 256226
rect 404998 256170 405054 256226
rect 405122 256170 405178 256226
rect 405246 256170 405302 256226
rect 404874 256046 404930 256102
rect 404998 256046 405054 256102
rect 405122 256046 405178 256102
rect 405246 256046 405302 256102
rect 404874 255922 404930 255978
rect 404998 255922 405054 255978
rect 405122 255922 405178 255978
rect 405246 255922 405302 255978
rect 404874 238294 404930 238350
rect 404998 238294 405054 238350
rect 405122 238294 405178 238350
rect 405246 238294 405302 238350
rect 404874 238170 404930 238226
rect 404998 238170 405054 238226
rect 405122 238170 405178 238226
rect 405246 238170 405302 238226
rect 404874 238046 404930 238102
rect 404998 238046 405054 238102
rect 405122 238046 405178 238102
rect 405246 238046 405302 238102
rect 404874 237922 404930 237978
rect 404998 237922 405054 237978
rect 405122 237922 405178 237978
rect 405246 237922 405302 237978
rect 404874 220294 404930 220350
rect 404998 220294 405054 220350
rect 405122 220294 405178 220350
rect 405246 220294 405302 220350
rect 404874 220170 404930 220226
rect 404998 220170 405054 220226
rect 405122 220170 405178 220226
rect 405246 220170 405302 220226
rect 404874 220046 404930 220102
rect 404998 220046 405054 220102
rect 405122 220046 405178 220102
rect 405246 220046 405302 220102
rect 404874 219922 404930 219978
rect 404998 219922 405054 219978
rect 405122 219922 405178 219978
rect 405246 219922 405302 219978
rect 404874 202294 404930 202350
rect 404998 202294 405054 202350
rect 405122 202294 405178 202350
rect 405246 202294 405302 202350
rect 404874 202170 404930 202226
rect 404998 202170 405054 202226
rect 405122 202170 405178 202226
rect 405246 202170 405302 202226
rect 404874 202046 404930 202102
rect 404998 202046 405054 202102
rect 405122 202046 405178 202102
rect 405246 202046 405302 202102
rect 404874 201922 404930 201978
rect 404998 201922 405054 201978
rect 405122 201922 405178 201978
rect 405246 201922 405302 201978
rect 404874 184294 404930 184350
rect 404998 184294 405054 184350
rect 405122 184294 405178 184350
rect 405246 184294 405302 184350
rect 404874 184170 404930 184226
rect 404998 184170 405054 184226
rect 405122 184170 405178 184226
rect 405246 184170 405302 184226
rect 404874 184046 404930 184102
rect 404998 184046 405054 184102
rect 405122 184046 405178 184102
rect 405246 184046 405302 184102
rect 404874 183922 404930 183978
rect 404998 183922 405054 183978
rect 405122 183922 405178 183978
rect 405246 183922 405302 183978
rect 404874 166294 404930 166350
rect 404998 166294 405054 166350
rect 405122 166294 405178 166350
rect 405246 166294 405302 166350
rect 404874 166170 404930 166226
rect 404998 166170 405054 166226
rect 405122 166170 405178 166226
rect 405246 166170 405302 166226
rect 404874 166046 404930 166102
rect 404998 166046 405054 166102
rect 405122 166046 405178 166102
rect 405246 166046 405302 166102
rect 404874 165922 404930 165978
rect 404998 165922 405054 165978
rect 405122 165922 405178 165978
rect 405246 165922 405302 165978
rect 404874 148294 404930 148350
rect 404998 148294 405054 148350
rect 405122 148294 405178 148350
rect 405246 148294 405302 148350
rect 404874 148170 404930 148226
rect 404998 148170 405054 148226
rect 405122 148170 405178 148226
rect 405246 148170 405302 148226
rect 404874 148046 404930 148102
rect 404998 148046 405054 148102
rect 405122 148046 405178 148102
rect 405246 148046 405302 148102
rect 404874 147922 404930 147978
rect 404998 147922 405054 147978
rect 405122 147922 405178 147978
rect 405246 147922 405302 147978
rect 404874 130294 404930 130350
rect 404998 130294 405054 130350
rect 405122 130294 405178 130350
rect 405246 130294 405302 130350
rect 404874 130170 404930 130226
rect 404998 130170 405054 130226
rect 405122 130170 405178 130226
rect 405246 130170 405302 130226
rect 404874 130046 404930 130102
rect 404998 130046 405054 130102
rect 405122 130046 405178 130102
rect 405246 130046 405302 130102
rect 404874 129922 404930 129978
rect 404998 129922 405054 129978
rect 405122 129922 405178 129978
rect 405246 129922 405302 129978
rect 404874 112294 404930 112350
rect 404998 112294 405054 112350
rect 405122 112294 405178 112350
rect 405246 112294 405302 112350
rect 404874 112170 404930 112226
rect 404998 112170 405054 112226
rect 405122 112170 405178 112226
rect 405246 112170 405302 112226
rect 404874 112046 404930 112102
rect 404998 112046 405054 112102
rect 405122 112046 405178 112102
rect 405246 112046 405302 112102
rect 404874 111922 404930 111978
rect 404998 111922 405054 111978
rect 405122 111922 405178 111978
rect 405246 111922 405302 111978
rect 404874 94294 404930 94350
rect 404998 94294 405054 94350
rect 405122 94294 405178 94350
rect 405246 94294 405302 94350
rect 404874 94170 404930 94226
rect 404998 94170 405054 94226
rect 405122 94170 405178 94226
rect 405246 94170 405302 94226
rect 404874 94046 404930 94102
rect 404998 94046 405054 94102
rect 405122 94046 405178 94102
rect 405246 94046 405302 94102
rect 404874 93922 404930 93978
rect 404998 93922 405054 93978
rect 405122 93922 405178 93978
rect 405246 93922 405302 93978
rect 404874 76294 404930 76350
rect 404998 76294 405054 76350
rect 405122 76294 405178 76350
rect 405246 76294 405302 76350
rect 404874 76170 404930 76226
rect 404998 76170 405054 76226
rect 405122 76170 405178 76226
rect 405246 76170 405302 76226
rect 404874 76046 404930 76102
rect 404998 76046 405054 76102
rect 405122 76046 405178 76102
rect 405246 76046 405302 76102
rect 404874 75922 404930 75978
rect 404998 75922 405054 75978
rect 405122 75922 405178 75978
rect 405246 75922 405302 75978
rect 377874 64294 377930 64350
rect 377998 64294 378054 64350
rect 378122 64294 378178 64350
rect 378246 64294 378302 64350
rect 377874 64170 377930 64226
rect 377998 64170 378054 64226
rect 378122 64170 378178 64226
rect 378246 64170 378302 64226
rect 377874 64046 377930 64102
rect 377998 64046 378054 64102
rect 378122 64046 378178 64102
rect 378246 64046 378302 64102
rect 377874 63922 377930 63978
rect 377998 63922 378054 63978
rect 378122 63922 378178 63978
rect 378246 63922 378302 63978
rect 374154 40294 374210 40350
rect 374278 40294 374334 40350
rect 374402 40294 374458 40350
rect 374526 40294 374582 40350
rect 374154 40170 374210 40226
rect 374278 40170 374334 40226
rect 374402 40170 374458 40226
rect 374526 40170 374582 40226
rect 374154 40046 374210 40102
rect 374278 40046 374334 40102
rect 374402 40046 374458 40102
rect 374526 40046 374582 40102
rect 374154 39922 374210 39978
rect 374278 39922 374334 39978
rect 374402 39922 374458 39978
rect 374526 39922 374582 39978
rect 371308 25622 371364 25678
rect 376348 55862 376404 55918
rect 374154 22294 374210 22350
rect 374278 22294 374334 22350
rect 374402 22294 374458 22350
rect 374526 22294 374582 22350
rect 374154 22170 374210 22226
rect 374278 22170 374334 22226
rect 374402 22170 374458 22226
rect 374526 22170 374582 22226
rect 374154 22046 374210 22102
rect 374278 22046 374334 22102
rect 374402 22046 374458 22102
rect 374526 22046 374582 22102
rect 374154 21922 374210 21978
rect 374278 21922 374334 21978
rect 374402 21922 374458 21978
rect 374526 21922 374582 21978
rect 374780 37142 374836 37198
rect 374154 4294 374210 4350
rect 374278 4294 374334 4350
rect 374402 4294 374458 4350
rect 374526 4294 374582 4350
rect 374154 4170 374210 4226
rect 374278 4170 374334 4226
rect 374402 4170 374458 4226
rect 374526 4170 374582 4226
rect 347154 -1176 347210 -1120
rect 347278 -1176 347334 -1120
rect 347402 -1176 347458 -1120
rect 347526 -1176 347582 -1120
rect 347154 -1300 347210 -1244
rect 347278 -1300 347334 -1244
rect 347402 -1300 347458 -1244
rect 347526 -1300 347582 -1244
rect 347154 -1424 347210 -1368
rect 347278 -1424 347334 -1368
rect 347402 -1424 347458 -1368
rect 347526 -1424 347582 -1368
rect 347154 -1548 347210 -1492
rect 347278 -1548 347334 -1492
rect 347402 -1548 347458 -1492
rect 347526 -1548 347582 -1492
rect 377874 46294 377930 46350
rect 377998 46294 378054 46350
rect 378122 46294 378178 46350
rect 378246 46294 378302 46350
rect 377874 46170 377930 46226
rect 377998 46170 378054 46226
rect 378122 46170 378178 46226
rect 378246 46170 378302 46226
rect 377874 46046 377930 46102
rect 377998 46046 378054 46102
rect 378122 46046 378178 46102
rect 378246 46046 378302 46102
rect 377874 45922 377930 45978
rect 377998 45922 378054 45978
rect 378122 45922 378178 45978
rect 378246 45922 378302 45978
rect 383068 72602 383124 72658
rect 377874 28294 377930 28350
rect 377998 28294 378054 28350
rect 378122 28294 378178 28350
rect 378246 28294 378302 28350
rect 377874 28170 377930 28226
rect 377998 28170 378054 28226
rect 378122 28170 378178 28226
rect 378246 28170 378302 28226
rect 377874 28046 377930 28102
rect 377998 28046 378054 28102
rect 378122 28046 378178 28102
rect 378246 28046 378302 28102
rect 377874 27922 377930 27978
rect 377998 27922 378054 27978
rect 378122 27922 378178 27978
rect 378246 27922 378302 27978
rect 377874 10294 377930 10350
rect 377998 10294 378054 10350
rect 378122 10294 378178 10350
rect 378246 10294 378302 10350
rect 377874 10170 377930 10226
rect 377998 10170 378054 10226
rect 378122 10170 378178 10226
rect 378246 10170 378302 10226
rect 377874 10046 377930 10102
rect 377998 10046 378054 10102
rect 378122 10046 378178 10102
rect 378246 10046 378302 10102
rect 377874 9922 377930 9978
rect 377998 9922 378054 9978
rect 378122 9922 378178 9978
rect 378246 9922 378302 9978
rect 374154 4046 374210 4102
rect 374278 4046 374334 4102
rect 374402 4046 374458 4102
rect 374526 4046 374582 4102
rect 374154 3922 374210 3978
rect 374278 3922 374334 3978
rect 374402 3922 374458 3978
rect 374526 3922 374582 3978
rect 374154 -216 374210 -160
rect 374278 -216 374334 -160
rect 374402 -216 374458 -160
rect 374526 -216 374582 -160
rect 374154 -340 374210 -284
rect 374278 -340 374334 -284
rect 374402 -340 374458 -284
rect 374526 -340 374582 -284
rect 374154 -464 374210 -408
rect 374278 -464 374334 -408
rect 374402 -464 374458 -408
rect 374526 -464 374582 -408
rect 374154 -588 374210 -532
rect 374278 -588 374334 -532
rect 374402 -588 374458 -532
rect 374526 -588 374582 -532
rect 379708 34082 379764 34138
rect 396508 60902 396564 60958
rect 386428 36962 386484 37018
rect 388108 23822 388164 23878
rect 391468 23642 391524 23698
rect 393148 12302 393204 12358
rect 394828 12122 394884 12178
rect 408594 598116 408650 598172
rect 408718 598116 408774 598172
rect 408842 598116 408898 598172
rect 408966 598116 409022 598172
rect 408594 597992 408650 598048
rect 408718 597992 408774 598048
rect 408842 597992 408898 598048
rect 408966 597992 409022 598048
rect 408594 597868 408650 597924
rect 408718 597868 408774 597924
rect 408842 597868 408898 597924
rect 408966 597868 409022 597924
rect 408594 597744 408650 597800
rect 408718 597744 408774 597800
rect 408842 597744 408898 597800
rect 408966 597744 409022 597800
rect 408594 586294 408650 586350
rect 408718 586294 408774 586350
rect 408842 586294 408898 586350
rect 408966 586294 409022 586350
rect 408594 586170 408650 586226
rect 408718 586170 408774 586226
rect 408842 586170 408898 586226
rect 408966 586170 409022 586226
rect 408594 586046 408650 586102
rect 408718 586046 408774 586102
rect 408842 586046 408898 586102
rect 408966 586046 409022 586102
rect 408594 585922 408650 585978
rect 408718 585922 408774 585978
rect 408842 585922 408898 585978
rect 408966 585922 409022 585978
rect 408594 568294 408650 568350
rect 408718 568294 408774 568350
rect 408842 568294 408898 568350
rect 408966 568294 409022 568350
rect 408594 568170 408650 568226
rect 408718 568170 408774 568226
rect 408842 568170 408898 568226
rect 408966 568170 409022 568226
rect 408594 568046 408650 568102
rect 408718 568046 408774 568102
rect 408842 568046 408898 568102
rect 408966 568046 409022 568102
rect 408594 567922 408650 567978
rect 408718 567922 408774 567978
rect 408842 567922 408898 567978
rect 408966 567922 409022 567978
rect 408594 550294 408650 550350
rect 408718 550294 408774 550350
rect 408842 550294 408898 550350
rect 408966 550294 409022 550350
rect 408594 550170 408650 550226
rect 408718 550170 408774 550226
rect 408842 550170 408898 550226
rect 408966 550170 409022 550226
rect 408594 550046 408650 550102
rect 408718 550046 408774 550102
rect 408842 550046 408898 550102
rect 408966 550046 409022 550102
rect 408594 549922 408650 549978
rect 408718 549922 408774 549978
rect 408842 549922 408898 549978
rect 408966 549922 409022 549978
rect 408594 532294 408650 532350
rect 408718 532294 408774 532350
rect 408842 532294 408898 532350
rect 408966 532294 409022 532350
rect 408594 532170 408650 532226
rect 408718 532170 408774 532226
rect 408842 532170 408898 532226
rect 408966 532170 409022 532226
rect 408594 532046 408650 532102
rect 408718 532046 408774 532102
rect 408842 532046 408898 532102
rect 408966 532046 409022 532102
rect 408594 531922 408650 531978
rect 408718 531922 408774 531978
rect 408842 531922 408898 531978
rect 408966 531922 409022 531978
rect 408594 514294 408650 514350
rect 408718 514294 408774 514350
rect 408842 514294 408898 514350
rect 408966 514294 409022 514350
rect 408594 514170 408650 514226
rect 408718 514170 408774 514226
rect 408842 514170 408898 514226
rect 408966 514170 409022 514226
rect 408594 514046 408650 514102
rect 408718 514046 408774 514102
rect 408842 514046 408898 514102
rect 408966 514046 409022 514102
rect 408594 513922 408650 513978
rect 408718 513922 408774 513978
rect 408842 513922 408898 513978
rect 408966 513922 409022 513978
rect 408594 496294 408650 496350
rect 408718 496294 408774 496350
rect 408842 496294 408898 496350
rect 408966 496294 409022 496350
rect 408594 496170 408650 496226
rect 408718 496170 408774 496226
rect 408842 496170 408898 496226
rect 408966 496170 409022 496226
rect 408594 496046 408650 496102
rect 408718 496046 408774 496102
rect 408842 496046 408898 496102
rect 408966 496046 409022 496102
rect 408594 495922 408650 495978
rect 408718 495922 408774 495978
rect 408842 495922 408898 495978
rect 408966 495922 409022 495978
rect 408594 478294 408650 478350
rect 408718 478294 408774 478350
rect 408842 478294 408898 478350
rect 408966 478294 409022 478350
rect 408594 478170 408650 478226
rect 408718 478170 408774 478226
rect 408842 478170 408898 478226
rect 408966 478170 409022 478226
rect 408594 478046 408650 478102
rect 408718 478046 408774 478102
rect 408842 478046 408898 478102
rect 408966 478046 409022 478102
rect 408594 477922 408650 477978
rect 408718 477922 408774 477978
rect 408842 477922 408898 477978
rect 408966 477922 409022 477978
rect 408594 460294 408650 460350
rect 408718 460294 408774 460350
rect 408842 460294 408898 460350
rect 408966 460294 409022 460350
rect 408594 460170 408650 460226
rect 408718 460170 408774 460226
rect 408842 460170 408898 460226
rect 408966 460170 409022 460226
rect 408594 460046 408650 460102
rect 408718 460046 408774 460102
rect 408842 460046 408898 460102
rect 408966 460046 409022 460102
rect 408594 459922 408650 459978
rect 408718 459922 408774 459978
rect 408842 459922 408898 459978
rect 408966 459922 409022 459978
rect 408594 442294 408650 442350
rect 408718 442294 408774 442350
rect 408842 442294 408898 442350
rect 408966 442294 409022 442350
rect 408594 442170 408650 442226
rect 408718 442170 408774 442226
rect 408842 442170 408898 442226
rect 408966 442170 409022 442226
rect 408594 442046 408650 442102
rect 408718 442046 408774 442102
rect 408842 442046 408898 442102
rect 408966 442046 409022 442102
rect 408594 441922 408650 441978
rect 408718 441922 408774 441978
rect 408842 441922 408898 441978
rect 408966 441922 409022 441978
rect 408594 424294 408650 424350
rect 408718 424294 408774 424350
rect 408842 424294 408898 424350
rect 408966 424294 409022 424350
rect 408594 424170 408650 424226
rect 408718 424170 408774 424226
rect 408842 424170 408898 424226
rect 408966 424170 409022 424226
rect 408594 424046 408650 424102
rect 408718 424046 408774 424102
rect 408842 424046 408898 424102
rect 408966 424046 409022 424102
rect 408594 423922 408650 423978
rect 408718 423922 408774 423978
rect 408842 423922 408898 423978
rect 408966 423922 409022 423978
rect 408594 406294 408650 406350
rect 408718 406294 408774 406350
rect 408842 406294 408898 406350
rect 408966 406294 409022 406350
rect 408594 406170 408650 406226
rect 408718 406170 408774 406226
rect 408842 406170 408898 406226
rect 408966 406170 409022 406226
rect 408594 406046 408650 406102
rect 408718 406046 408774 406102
rect 408842 406046 408898 406102
rect 408966 406046 409022 406102
rect 408594 405922 408650 405978
rect 408718 405922 408774 405978
rect 408842 405922 408898 405978
rect 408966 405922 409022 405978
rect 408594 388294 408650 388350
rect 408718 388294 408774 388350
rect 408842 388294 408898 388350
rect 408966 388294 409022 388350
rect 408594 388170 408650 388226
rect 408718 388170 408774 388226
rect 408842 388170 408898 388226
rect 408966 388170 409022 388226
rect 408594 388046 408650 388102
rect 408718 388046 408774 388102
rect 408842 388046 408898 388102
rect 408966 388046 409022 388102
rect 408594 387922 408650 387978
rect 408718 387922 408774 387978
rect 408842 387922 408898 387978
rect 408966 387922 409022 387978
rect 408594 370294 408650 370350
rect 408718 370294 408774 370350
rect 408842 370294 408898 370350
rect 408966 370294 409022 370350
rect 408594 370170 408650 370226
rect 408718 370170 408774 370226
rect 408842 370170 408898 370226
rect 408966 370170 409022 370226
rect 408594 370046 408650 370102
rect 408718 370046 408774 370102
rect 408842 370046 408898 370102
rect 408966 370046 409022 370102
rect 408594 369922 408650 369978
rect 408718 369922 408774 369978
rect 408842 369922 408898 369978
rect 408966 369922 409022 369978
rect 408594 352294 408650 352350
rect 408718 352294 408774 352350
rect 408842 352294 408898 352350
rect 408966 352294 409022 352350
rect 408594 352170 408650 352226
rect 408718 352170 408774 352226
rect 408842 352170 408898 352226
rect 408966 352170 409022 352226
rect 408594 352046 408650 352102
rect 408718 352046 408774 352102
rect 408842 352046 408898 352102
rect 408966 352046 409022 352102
rect 408594 351922 408650 351978
rect 408718 351922 408774 351978
rect 408842 351922 408898 351978
rect 408966 351922 409022 351978
rect 408594 334294 408650 334350
rect 408718 334294 408774 334350
rect 408842 334294 408898 334350
rect 408966 334294 409022 334350
rect 408594 334170 408650 334226
rect 408718 334170 408774 334226
rect 408842 334170 408898 334226
rect 408966 334170 409022 334226
rect 408594 334046 408650 334102
rect 408718 334046 408774 334102
rect 408842 334046 408898 334102
rect 408966 334046 409022 334102
rect 408594 333922 408650 333978
rect 408718 333922 408774 333978
rect 408842 333922 408898 333978
rect 408966 333922 409022 333978
rect 408594 316294 408650 316350
rect 408718 316294 408774 316350
rect 408842 316294 408898 316350
rect 408966 316294 409022 316350
rect 408594 316170 408650 316226
rect 408718 316170 408774 316226
rect 408842 316170 408898 316226
rect 408966 316170 409022 316226
rect 408594 316046 408650 316102
rect 408718 316046 408774 316102
rect 408842 316046 408898 316102
rect 408966 316046 409022 316102
rect 408594 315922 408650 315978
rect 408718 315922 408774 315978
rect 408842 315922 408898 315978
rect 408966 315922 409022 315978
rect 408594 298294 408650 298350
rect 408718 298294 408774 298350
rect 408842 298294 408898 298350
rect 408966 298294 409022 298350
rect 408594 298170 408650 298226
rect 408718 298170 408774 298226
rect 408842 298170 408898 298226
rect 408966 298170 409022 298226
rect 408594 298046 408650 298102
rect 408718 298046 408774 298102
rect 408842 298046 408898 298102
rect 408966 298046 409022 298102
rect 408594 297922 408650 297978
rect 408718 297922 408774 297978
rect 408842 297922 408898 297978
rect 408966 297922 409022 297978
rect 408594 280294 408650 280350
rect 408718 280294 408774 280350
rect 408842 280294 408898 280350
rect 408966 280294 409022 280350
rect 408594 280170 408650 280226
rect 408718 280170 408774 280226
rect 408842 280170 408898 280226
rect 408966 280170 409022 280226
rect 408594 280046 408650 280102
rect 408718 280046 408774 280102
rect 408842 280046 408898 280102
rect 408966 280046 409022 280102
rect 408594 279922 408650 279978
rect 408718 279922 408774 279978
rect 408842 279922 408898 279978
rect 408966 279922 409022 279978
rect 408594 262294 408650 262350
rect 408718 262294 408774 262350
rect 408842 262294 408898 262350
rect 408966 262294 409022 262350
rect 408594 262170 408650 262226
rect 408718 262170 408774 262226
rect 408842 262170 408898 262226
rect 408966 262170 409022 262226
rect 408594 262046 408650 262102
rect 408718 262046 408774 262102
rect 408842 262046 408898 262102
rect 408966 262046 409022 262102
rect 408594 261922 408650 261978
rect 408718 261922 408774 261978
rect 408842 261922 408898 261978
rect 408966 261922 409022 261978
rect 408594 244294 408650 244350
rect 408718 244294 408774 244350
rect 408842 244294 408898 244350
rect 408966 244294 409022 244350
rect 408594 244170 408650 244226
rect 408718 244170 408774 244226
rect 408842 244170 408898 244226
rect 408966 244170 409022 244226
rect 408594 244046 408650 244102
rect 408718 244046 408774 244102
rect 408842 244046 408898 244102
rect 408966 244046 409022 244102
rect 408594 243922 408650 243978
rect 408718 243922 408774 243978
rect 408842 243922 408898 243978
rect 408966 243922 409022 243978
rect 408594 226294 408650 226350
rect 408718 226294 408774 226350
rect 408842 226294 408898 226350
rect 408966 226294 409022 226350
rect 408594 226170 408650 226226
rect 408718 226170 408774 226226
rect 408842 226170 408898 226226
rect 408966 226170 409022 226226
rect 408594 226046 408650 226102
rect 408718 226046 408774 226102
rect 408842 226046 408898 226102
rect 408966 226046 409022 226102
rect 408594 225922 408650 225978
rect 408718 225922 408774 225978
rect 408842 225922 408898 225978
rect 408966 225922 409022 225978
rect 408594 208294 408650 208350
rect 408718 208294 408774 208350
rect 408842 208294 408898 208350
rect 408966 208294 409022 208350
rect 408594 208170 408650 208226
rect 408718 208170 408774 208226
rect 408842 208170 408898 208226
rect 408966 208170 409022 208226
rect 408594 208046 408650 208102
rect 408718 208046 408774 208102
rect 408842 208046 408898 208102
rect 408966 208046 409022 208102
rect 408594 207922 408650 207978
rect 408718 207922 408774 207978
rect 408842 207922 408898 207978
rect 408966 207922 409022 207978
rect 408594 190294 408650 190350
rect 408718 190294 408774 190350
rect 408842 190294 408898 190350
rect 408966 190294 409022 190350
rect 408594 190170 408650 190226
rect 408718 190170 408774 190226
rect 408842 190170 408898 190226
rect 408966 190170 409022 190226
rect 408594 190046 408650 190102
rect 408718 190046 408774 190102
rect 408842 190046 408898 190102
rect 408966 190046 409022 190102
rect 408594 189922 408650 189978
rect 408718 189922 408774 189978
rect 408842 189922 408898 189978
rect 408966 189922 409022 189978
rect 408594 172294 408650 172350
rect 408718 172294 408774 172350
rect 408842 172294 408898 172350
rect 408966 172294 409022 172350
rect 408594 172170 408650 172226
rect 408718 172170 408774 172226
rect 408842 172170 408898 172226
rect 408966 172170 409022 172226
rect 408594 172046 408650 172102
rect 408718 172046 408774 172102
rect 408842 172046 408898 172102
rect 408966 172046 409022 172102
rect 408594 171922 408650 171978
rect 408718 171922 408774 171978
rect 408842 171922 408898 171978
rect 408966 171922 409022 171978
rect 408594 154294 408650 154350
rect 408718 154294 408774 154350
rect 408842 154294 408898 154350
rect 408966 154294 409022 154350
rect 408594 154170 408650 154226
rect 408718 154170 408774 154226
rect 408842 154170 408898 154226
rect 408966 154170 409022 154226
rect 408594 154046 408650 154102
rect 408718 154046 408774 154102
rect 408842 154046 408898 154102
rect 408966 154046 409022 154102
rect 408594 153922 408650 153978
rect 408718 153922 408774 153978
rect 408842 153922 408898 153978
rect 408966 153922 409022 153978
rect 408594 136294 408650 136350
rect 408718 136294 408774 136350
rect 408842 136294 408898 136350
rect 408966 136294 409022 136350
rect 408594 136170 408650 136226
rect 408718 136170 408774 136226
rect 408842 136170 408898 136226
rect 408966 136170 409022 136226
rect 408594 136046 408650 136102
rect 408718 136046 408774 136102
rect 408842 136046 408898 136102
rect 408966 136046 409022 136102
rect 408594 135922 408650 135978
rect 408718 135922 408774 135978
rect 408842 135922 408898 135978
rect 408966 135922 409022 135978
rect 408594 118294 408650 118350
rect 408718 118294 408774 118350
rect 408842 118294 408898 118350
rect 408966 118294 409022 118350
rect 408594 118170 408650 118226
rect 408718 118170 408774 118226
rect 408842 118170 408898 118226
rect 408966 118170 409022 118226
rect 408594 118046 408650 118102
rect 408718 118046 408774 118102
rect 408842 118046 408898 118102
rect 408966 118046 409022 118102
rect 408594 117922 408650 117978
rect 408718 117922 408774 117978
rect 408842 117922 408898 117978
rect 408966 117922 409022 117978
rect 408594 100294 408650 100350
rect 408718 100294 408774 100350
rect 408842 100294 408898 100350
rect 408966 100294 409022 100350
rect 408594 100170 408650 100226
rect 408718 100170 408774 100226
rect 408842 100170 408898 100226
rect 408966 100170 409022 100226
rect 408594 100046 408650 100102
rect 408718 100046 408774 100102
rect 408842 100046 408898 100102
rect 408966 100046 409022 100102
rect 408594 99922 408650 99978
rect 408718 99922 408774 99978
rect 408842 99922 408898 99978
rect 408966 99922 409022 99978
rect 408594 82294 408650 82350
rect 408718 82294 408774 82350
rect 408842 82294 408898 82350
rect 408966 82294 409022 82350
rect 408594 82170 408650 82226
rect 408718 82170 408774 82226
rect 408842 82170 408898 82226
rect 408966 82170 409022 82226
rect 408594 82046 408650 82102
rect 408718 82046 408774 82102
rect 408842 82046 408898 82102
rect 408966 82046 409022 82102
rect 408594 81922 408650 81978
rect 408718 81922 408774 81978
rect 408842 81922 408898 81978
rect 408966 81922 409022 81978
rect 404874 58294 404930 58350
rect 404998 58294 405054 58350
rect 405122 58294 405178 58350
rect 405246 58294 405302 58350
rect 404874 58170 404930 58226
rect 404998 58170 405054 58226
rect 405122 58170 405178 58226
rect 405246 58170 405302 58226
rect 404874 58046 404930 58102
rect 404998 58046 405054 58102
rect 405122 58046 405178 58102
rect 405246 58046 405302 58102
rect 404874 57922 404930 57978
rect 404998 57922 405054 57978
rect 405122 57922 405178 57978
rect 405246 57922 405302 57978
rect 404874 40294 404930 40350
rect 404998 40294 405054 40350
rect 405122 40294 405178 40350
rect 405246 40294 405302 40350
rect 404874 40170 404930 40226
rect 404998 40170 405054 40226
rect 405122 40170 405178 40226
rect 405246 40170 405302 40226
rect 404874 40046 404930 40102
rect 404998 40046 405054 40102
rect 405122 40046 405178 40102
rect 405246 40046 405302 40102
rect 404874 39922 404930 39978
rect 404998 39922 405054 39978
rect 405122 39922 405178 39978
rect 405246 39922 405302 39978
rect 403228 33722 403284 33778
rect 404874 22294 404930 22350
rect 404998 22294 405054 22350
rect 405122 22294 405178 22350
rect 405246 22294 405302 22350
rect 404874 22170 404930 22226
rect 404998 22170 405054 22226
rect 405122 22170 405178 22226
rect 405246 22170 405302 22226
rect 404874 22046 404930 22102
rect 404998 22046 405054 22102
rect 405122 22046 405178 22102
rect 405246 22046 405302 22102
rect 404874 21922 404930 21978
rect 404998 21922 405054 21978
rect 405122 21922 405178 21978
rect 405246 21922 405302 21978
rect 404874 4294 404930 4350
rect 404998 4294 405054 4350
rect 405122 4294 405178 4350
rect 405246 4294 405302 4350
rect 404874 4170 404930 4226
rect 404998 4170 405054 4226
rect 405122 4170 405178 4226
rect 405246 4170 405302 4226
rect 377874 -1176 377930 -1120
rect 377998 -1176 378054 -1120
rect 378122 -1176 378178 -1120
rect 378246 -1176 378302 -1120
rect 377874 -1300 377930 -1244
rect 377998 -1300 378054 -1244
rect 378122 -1300 378178 -1244
rect 378246 -1300 378302 -1244
rect 377874 -1424 377930 -1368
rect 377998 -1424 378054 -1368
rect 378122 -1424 378178 -1368
rect 378246 -1424 378302 -1368
rect 377874 -1548 377930 -1492
rect 377998 -1548 378054 -1492
rect 378122 -1548 378178 -1492
rect 378246 -1548 378302 -1492
rect 406588 65762 406644 65818
rect 435594 597156 435650 597212
rect 435718 597156 435774 597212
rect 435842 597156 435898 597212
rect 435966 597156 436022 597212
rect 435594 597032 435650 597088
rect 435718 597032 435774 597088
rect 435842 597032 435898 597088
rect 435966 597032 436022 597088
rect 435594 596908 435650 596964
rect 435718 596908 435774 596964
rect 435842 596908 435898 596964
rect 435966 596908 436022 596964
rect 435594 596784 435650 596840
rect 435718 596784 435774 596840
rect 435842 596784 435898 596840
rect 435966 596784 436022 596840
rect 435594 580294 435650 580350
rect 435718 580294 435774 580350
rect 435842 580294 435898 580350
rect 435966 580294 436022 580350
rect 435594 580170 435650 580226
rect 435718 580170 435774 580226
rect 435842 580170 435898 580226
rect 435966 580170 436022 580226
rect 435594 580046 435650 580102
rect 435718 580046 435774 580102
rect 435842 580046 435898 580102
rect 435966 580046 436022 580102
rect 435594 579922 435650 579978
rect 435718 579922 435774 579978
rect 435842 579922 435898 579978
rect 435966 579922 436022 579978
rect 435594 562294 435650 562350
rect 435718 562294 435774 562350
rect 435842 562294 435898 562350
rect 435966 562294 436022 562350
rect 435594 562170 435650 562226
rect 435718 562170 435774 562226
rect 435842 562170 435898 562226
rect 435966 562170 436022 562226
rect 435594 562046 435650 562102
rect 435718 562046 435774 562102
rect 435842 562046 435898 562102
rect 435966 562046 436022 562102
rect 435594 561922 435650 561978
rect 435718 561922 435774 561978
rect 435842 561922 435898 561978
rect 435966 561922 436022 561978
rect 435594 544294 435650 544350
rect 435718 544294 435774 544350
rect 435842 544294 435898 544350
rect 435966 544294 436022 544350
rect 435594 544170 435650 544226
rect 435718 544170 435774 544226
rect 435842 544170 435898 544226
rect 435966 544170 436022 544226
rect 435594 544046 435650 544102
rect 435718 544046 435774 544102
rect 435842 544046 435898 544102
rect 435966 544046 436022 544102
rect 435594 543922 435650 543978
rect 435718 543922 435774 543978
rect 435842 543922 435898 543978
rect 435966 543922 436022 543978
rect 435594 526294 435650 526350
rect 435718 526294 435774 526350
rect 435842 526294 435898 526350
rect 435966 526294 436022 526350
rect 435594 526170 435650 526226
rect 435718 526170 435774 526226
rect 435842 526170 435898 526226
rect 435966 526170 436022 526226
rect 435594 526046 435650 526102
rect 435718 526046 435774 526102
rect 435842 526046 435898 526102
rect 435966 526046 436022 526102
rect 435594 525922 435650 525978
rect 435718 525922 435774 525978
rect 435842 525922 435898 525978
rect 435966 525922 436022 525978
rect 435594 508294 435650 508350
rect 435718 508294 435774 508350
rect 435842 508294 435898 508350
rect 435966 508294 436022 508350
rect 435594 508170 435650 508226
rect 435718 508170 435774 508226
rect 435842 508170 435898 508226
rect 435966 508170 436022 508226
rect 435594 508046 435650 508102
rect 435718 508046 435774 508102
rect 435842 508046 435898 508102
rect 435966 508046 436022 508102
rect 435594 507922 435650 507978
rect 435718 507922 435774 507978
rect 435842 507922 435898 507978
rect 435966 507922 436022 507978
rect 435594 490294 435650 490350
rect 435718 490294 435774 490350
rect 435842 490294 435898 490350
rect 435966 490294 436022 490350
rect 435594 490170 435650 490226
rect 435718 490170 435774 490226
rect 435842 490170 435898 490226
rect 435966 490170 436022 490226
rect 435594 490046 435650 490102
rect 435718 490046 435774 490102
rect 435842 490046 435898 490102
rect 435966 490046 436022 490102
rect 435594 489922 435650 489978
rect 435718 489922 435774 489978
rect 435842 489922 435898 489978
rect 435966 489922 436022 489978
rect 435594 472294 435650 472350
rect 435718 472294 435774 472350
rect 435842 472294 435898 472350
rect 435966 472294 436022 472350
rect 435594 472170 435650 472226
rect 435718 472170 435774 472226
rect 435842 472170 435898 472226
rect 435966 472170 436022 472226
rect 435594 472046 435650 472102
rect 435718 472046 435774 472102
rect 435842 472046 435898 472102
rect 435966 472046 436022 472102
rect 435594 471922 435650 471978
rect 435718 471922 435774 471978
rect 435842 471922 435898 471978
rect 435966 471922 436022 471978
rect 435594 454294 435650 454350
rect 435718 454294 435774 454350
rect 435842 454294 435898 454350
rect 435966 454294 436022 454350
rect 435594 454170 435650 454226
rect 435718 454170 435774 454226
rect 435842 454170 435898 454226
rect 435966 454170 436022 454226
rect 435594 454046 435650 454102
rect 435718 454046 435774 454102
rect 435842 454046 435898 454102
rect 435966 454046 436022 454102
rect 435594 453922 435650 453978
rect 435718 453922 435774 453978
rect 435842 453922 435898 453978
rect 435966 453922 436022 453978
rect 435594 436294 435650 436350
rect 435718 436294 435774 436350
rect 435842 436294 435898 436350
rect 435966 436294 436022 436350
rect 435594 436170 435650 436226
rect 435718 436170 435774 436226
rect 435842 436170 435898 436226
rect 435966 436170 436022 436226
rect 435594 436046 435650 436102
rect 435718 436046 435774 436102
rect 435842 436046 435898 436102
rect 435966 436046 436022 436102
rect 435594 435922 435650 435978
rect 435718 435922 435774 435978
rect 435842 435922 435898 435978
rect 435966 435922 436022 435978
rect 435594 418294 435650 418350
rect 435718 418294 435774 418350
rect 435842 418294 435898 418350
rect 435966 418294 436022 418350
rect 435594 418170 435650 418226
rect 435718 418170 435774 418226
rect 435842 418170 435898 418226
rect 435966 418170 436022 418226
rect 435594 418046 435650 418102
rect 435718 418046 435774 418102
rect 435842 418046 435898 418102
rect 435966 418046 436022 418102
rect 435594 417922 435650 417978
rect 435718 417922 435774 417978
rect 435842 417922 435898 417978
rect 435966 417922 436022 417978
rect 435594 400294 435650 400350
rect 435718 400294 435774 400350
rect 435842 400294 435898 400350
rect 435966 400294 436022 400350
rect 435594 400170 435650 400226
rect 435718 400170 435774 400226
rect 435842 400170 435898 400226
rect 435966 400170 436022 400226
rect 435594 400046 435650 400102
rect 435718 400046 435774 400102
rect 435842 400046 435898 400102
rect 435966 400046 436022 400102
rect 435594 399922 435650 399978
rect 435718 399922 435774 399978
rect 435842 399922 435898 399978
rect 435966 399922 436022 399978
rect 435594 382294 435650 382350
rect 435718 382294 435774 382350
rect 435842 382294 435898 382350
rect 435966 382294 436022 382350
rect 435594 382170 435650 382226
rect 435718 382170 435774 382226
rect 435842 382170 435898 382226
rect 435966 382170 436022 382226
rect 435594 382046 435650 382102
rect 435718 382046 435774 382102
rect 435842 382046 435898 382102
rect 435966 382046 436022 382102
rect 435594 381922 435650 381978
rect 435718 381922 435774 381978
rect 435842 381922 435898 381978
rect 435966 381922 436022 381978
rect 435594 364294 435650 364350
rect 435718 364294 435774 364350
rect 435842 364294 435898 364350
rect 435966 364294 436022 364350
rect 435594 364170 435650 364226
rect 435718 364170 435774 364226
rect 435842 364170 435898 364226
rect 435966 364170 436022 364226
rect 435594 364046 435650 364102
rect 435718 364046 435774 364102
rect 435842 364046 435898 364102
rect 435966 364046 436022 364102
rect 435594 363922 435650 363978
rect 435718 363922 435774 363978
rect 435842 363922 435898 363978
rect 435966 363922 436022 363978
rect 435594 346294 435650 346350
rect 435718 346294 435774 346350
rect 435842 346294 435898 346350
rect 435966 346294 436022 346350
rect 435594 346170 435650 346226
rect 435718 346170 435774 346226
rect 435842 346170 435898 346226
rect 435966 346170 436022 346226
rect 435594 346046 435650 346102
rect 435718 346046 435774 346102
rect 435842 346046 435898 346102
rect 435966 346046 436022 346102
rect 435594 345922 435650 345978
rect 435718 345922 435774 345978
rect 435842 345922 435898 345978
rect 435966 345922 436022 345978
rect 435594 328294 435650 328350
rect 435718 328294 435774 328350
rect 435842 328294 435898 328350
rect 435966 328294 436022 328350
rect 435594 328170 435650 328226
rect 435718 328170 435774 328226
rect 435842 328170 435898 328226
rect 435966 328170 436022 328226
rect 435594 328046 435650 328102
rect 435718 328046 435774 328102
rect 435842 328046 435898 328102
rect 435966 328046 436022 328102
rect 435594 327922 435650 327978
rect 435718 327922 435774 327978
rect 435842 327922 435898 327978
rect 435966 327922 436022 327978
rect 435594 310294 435650 310350
rect 435718 310294 435774 310350
rect 435842 310294 435898 310350
rect 435966 310294 436022 310350
rect 435594 310170 435650 310226
rect 435718 310170 435774 310226
rect 435842 310170 435898 310226
rect 435966 310170 436022 310226
rect 435594 310046 435650 310102
rect 435718 310046 435774 310102
rect 435842 310046 435898 310102
rect 435966 310046 436022 310102
rect 435594 309922 435650 309978
rect 435718 309922 435774 309978
rect 435842 309922 435898 309978
rect 435966 309922 436022 309978
rect 435594 292294 435650 292350
rect 435718 292294 435774 292350
rect 435842 292294 435898 292350
rect 435966 292294 436022 292350
rect 435594 292170 435650 292226
rect 435718 292170 435774 292226
rect 435842 292170 435898 292226
rect 435966 292170 436022 292226
rect 435594 292046 435650 292102
rect 435718 292046 435774 292102
rect 435842 292046 435898 292102
rect 435966 292046 436022 292102
rect 435594 291922 435650 291978
rect 435718 291922 435774 291978
rect 435842 291922 435898 291978
rect 435966 291922 436022 291978
rect 435594 274294 435650 274350
rect 435718 274294 435774 274350
rect 435842 274294 435898 274350
rect 435966 274294 436022 274350
rect 435594 274170 435650 274226
rect 435718 274170 435774 274226
rect 435842 274170 435898 274226
rect 435966 274170 436022 274226
rect 435594 274046 435650 274102
rect 435718 274046 435774 274102
rect 435842 274046 435898 274102
rect 435966 274046 436022 274102
rect 435594 273922 435650 273978
rect 435718 273922 435774 273978
rect 435842 273922 435898 273978
rect 435966 273922 436022 273978
rect 435594 256294 435650 256350
rect 435718 256294 435774 256350
rect 435842 256294 435898 256350
rect 435966 256294 436022 256350
rect 435594 256170 435650 256226
rect 435718 256170 435774 256226
rect 435842 256170 435898 256226
rect 435966 256170 436022 256226
rect 435594 256046 435650 256102
rect 435718 256046 435774 256102
rect 435842 256046 435898 256102
rect 435966 256046 436022 256102
rect 435594 255922 435650 255978
rect 435718 255922 435774 255978
rect 435842 255922 435898 255978
rect 435966 255922 436022 255978
rect 435594 238294 435650 238350
rect 435718 238294 435774 238350
rect 435842 238294 435898 238350
rect 435966 238294 436022 238350
rect 435594 238170 435650 238226
rect 435718 238170 435774 238226
rect 435842 238170 435898 238226
rect 435966 238170 436022 238226
rect 435594 238046 435650 238102
rect 435718 238046 435774 238102
rect 435842 238046 435898 238102
rect 435966 238046 436022 238102
rect 435594 237922 435650 237978
rect 435718 237922 435774 237978
rect 435842 237922 435898 237978
rect 435966 237922 436022 237978
rect 435594 220294 435650 220350
rect 435718 220294 435774 220350
rect 435842 220294 435898 220350
rect 435966 220294 436022 220350
rect 435594 220170 435650 220226
rect 435718 220170 435774 220226
rect 435842 220170 435898 220226
rect 435966 220170 436022 220226
rect 435594 220046 435650 220102
rect 435718 220046 435774 220102
rect 435842 220046 435898 220102
rect 435966 220046 436022 220102
rect 435594 219922 435650 219978
rect 435718 219922 435774 219978
rect 435842 219922 435898 219978
rect 435966 219922 436022 219978
rect 435594 202294 435650 202350
rect 435718 202294 435774 202350
rect 435842 202294 435898 202350
rect 435966 202294 436022 202350
rect 435594 202170 435650 202226
rect 435718 202170 435774 202226
rect 435842 202170 435898 202226
rect 435966 202170 436022 202226
rect 435594 202046 435650 202102
rect 435718 202046 435774 202102
rect 435842 202046 435898 202102
rect 435966 202046 436022 202102
rect 435594 201922 435650 201978
rect 435718 201922 435774 201978
rect 435842 201922 435898 201978
rect 435966 201922 436022 201978
rect 435594 184294 435650 184350
rect 435718 184294 435774 184350
rect 435842 184294 435898 184350
rect 435966 184294 436022 184350
rect 435594 184170 435650 184226
rect 435718 184170 435774 184226
rect 435842 184170 435898 184226
rect 435966 184170 436022 184226
rect 435594 184046 435650 184102
rect 435718 184046 435774 184102
rect 435842 184046 435898 184102
rect 435966 184046 436022 184102
rect 435594 183922 435650 183978
rect 435718 183922 435774 183978
rect 435842 183922 435898 183978
rect 435966 183922 436022 183978
rect 435594 166294 435650 166350
rect 435718 166294 435774 166350
rect 435842 166294 435898 166350
rect 435966 166294 436022 166350
rect 435594 166170 435650 166226
rect 435718 166170 435774 166226
rect 435842 166170 435898 166226
rect 435966 166170 436022 166226
rect 435594 166046 435650 166102
rect 435718 166046 435774 166102
rect 435842 166046 435898 166102
rect 435966 166046 436022 166102
rect 435594 165922 435650 165978
rect 435718 165922 435774 165978
rect 435842 165922 435898 165978
rect 435966 165922 436022 165978
rect 435594 148294 435650 148350
rect 435718 148294 435774 148350
rect 435842 148294 435898 148350
rect 435966 148294 436022 148350
rect 435594 148170 435650 148226
rect 435718 148170 435774 148226
rect 435842 148170 435898 148226
rect 435966 148170 436022 148226
rect 435594 148046 435650 148102
rect 435718 148046 435774 148102
rect 435842 148046 435898 148102
rect 435966 148046 436022 148102
rect 435594 147922 435650 147978
rect 435718 147922 435774 147978
rect 435842 147922 435898 147978
rect 435966 147922 436022 147978
rect 435594 130294 435650 130350
rect 435718 130294 435774 130350
rect 435842 130294 435898 130350
rect 435966 130294 436022 130350
rect 435594 130170 435650 130226
rect 435718 130170 435774 130226
rect 435842 130170 435898 130226
rect 435966 130170 436022 130226
rect 435594 130046 435650 130102
rect 435718 130046 435774 130102
rect 435842 130046 435898 130102
rect 435966 130046 436022 130102
rect 435594 129922 435650 129978
rect 435718 129922 435774 129978
rect 435842 129922 435898 129978
rect 435966 129922 436022 129978
rect 435594 112294 435650 112350
rect 435718 112294 435774 112350
rect 435842 112294 435898 112350
rect 435966 112294 436022 112350
rect 435594 112170 435650 112226
rect 435718 112170 435774 112226
rect 435842 112170 435898 112226
rect 435966 112170 436022 112226
rect 435594 112046 435650 112102
rect 435718 112046 435774 112102
rect 435842 112046 435898 112102
rect 435966 112046 436022 112102
rect 435594 111922 435650 111978
rect 435718 111922 435774 111978
rect 435842 111922 435898 111978
rect 435966 111922 436022 111978
rect 435594 94294 435650 94350
rect 435718 94294 435774 94350
rect 435842 94294 435898 94350
rect 435966 94294 436022 94350
rect 435594 94170 435650 94226
rect 435718 94170 435774 94226
rect 435842 94170 435898 94226
rect 435966 94170 436022 94226
rect 435594 94046 435650 94102
rect 435718 94046 435774 94102
rect 435842 94046 435898 94102
rect 435966 94046 436022 94102
rect 435594 93922 435650 93978
rect 435718 93922 435774 93978
rect 435842 93922 435898 93978
rect 435966 93922 436022 93978
rect 435594 76294 435650 76350
rect 435718 76294 435774 76350
rect 435842 76294 435898 76350
rect 435966 76294 436022 76350
rect 435594 76170 435650 76226
rect 435718 76170 435774 76226
rect 435842 76170 435898 76226
rect 435966 76170 436022 76226
rect 435594 76046 435650 76102
rect 435718 76046 435774 76102
rect 435842 76046 435898 76102
rect 435966 76046 436022 76102
rect 435594 75922 435650 75978
rect 435718 75922 435774 75978
rect 435842 75922 435898 75978
rect 435966 75922 436022 75978
rect 435148 72422 435204 72478
rect 408594 64294 408650 64350
rect 408718 64294 408774 64350
rect 408842 64294 408898 64350
rect 408966 64294 409022 64350
rect 408594 64170 408650 64226
rect 408718 64170 408774 64226
rect 408842 64170 408898 64226
rect 408966 64170 409022 64226
rect 408594 64046 408650 64102
rect 408718 64046 408774 64102
rect 408842 64046 408898 64102
rect 408966 64046 409022 64102
rect 408594 63922 408650 63978
rect 408718 63922 408774 63978
rect 408842 63922 408898 63978
rect 408966 63922 409022 63978
rect 408594 46294 408650 46350
rect 408718 46294 408774 46350
rect 408842 46294 408898 46350
rect 408966 46294 409022 46350
rect 408594 46170 408650 46226
rect 408718 46170 408774 46226
rect 408842 46170 408898 46226
rect 408966 46170 409022 46226
rect 408594 46046 408650 46102
rect 408718 46046 408774 46102
rect 408842 46046 408898 46102
rect 408966 46046 409022 46102
rect 408594 45922 408650 45978
rect 408718 45922 408774 45978
rect 408842 45922 408898 45978
rect 408966 45922 409022 45978
rect 431788 67382 431844 67438
rect 408594 28294 408650 28350
rect 408718 28294 408774 28350
rect 408842 28294 408898 28350
rect 408966 28294 409022 28350
rect 408594 28170 408650 28226
rect 408718 28170 408774 28226
rect 408842 28170 408898 28226
rect 408966 28170 409022 28226
rect 408594 28046 408650 28102
rect 408718 28046 408774 28102
rect 408842 28046 408898 28102
rect 408966 28046 409022 28102
rect 408594 27922 408650 27978
rect 408718 27922 408774 27978
rect 408842 27922 408898 27978
rect 408966 27922 409022 27978
rect 416668 42002 416724 42058
rect 425068 35522 425124 35578
rect 420028 33902 420084 33958
rect 408594 10294 408650 10350
rect 408718 10294 408774 10350
rect 408842 10294 408898 10350
rect 408966 10294 409022 10350
rect 408594 10170 408650 10226
rect 408718 10170 408774 10226
rect 408842 10170 408898 10226
rect 408966 10170 409022 10226
rect 408594 10046 408650 10102
rect 408718 10046 408774 10102
rect 408842 10046 408898 10102
rect 408966 10046 409022 10102
rect 408594 9922 408650 9978
rect 408718 9922 408774 9978
rect 408842 9922 408898 9978
rect 408966 9922 409022 9978
rect 404874 4046 404930 4102
rect 404998 4046 405054 4102
rect 405122 4046 405178 4102
rect 405246 4046 405302 4102
rect 404874 3922 404930 3978
rect 404998 3922 405054 3978
rect 405122 3922 405178 3978
rect 405246 3922 405302 3978
rect 404874 -216 404930 -160
rect 404998 -216 405054 -160
rect 405122 -216 405178 -160
rect 405246 -216 405302 -160
rect 404874 -340 404930 -284
rect 404998 -340 405054 -284
rect 405122 -340 405178 -284
rect 405246 -340 405302 -284
rect 404874 -464 404930 -408
rect 404998 -464 405054 -408
rect 405122 -464 405178 -408
rect 405246 -464 405302 -408
rect 404874 -588 404930 -532
rect 404998 -588 405054 -532
rect 405122 -588 405178 -532
rect 405246 -588 405302 -532
rect 409948 16982 410004 17038
rect 409276 5822 409332 5878
rect 414988 5282 415044 5338
rect 422604 8702 422660 8758
rect 428428 28862 428484 28918
rect 435594 58294 435650 58350
rect 435718 58294 435774 58350
rect 435842 58294 435898 58350
rect 435966 58294 436022 58350
rect 435594 58170 435650 58226
rect 435718 58170 435774 58226
rect 435842 58170 435898 58226
rect 435966 58170 436022 58226
rect 435594 58046 435650 58102
rect 435718 58046 435774 58102
rect 435842 58046 435898 58102
rect 435966 58046 436022 58102
rect 435594 57922 435650 57978
rect 435718 57922 435774 57978
rect 435842 57922 435898 57978
rect 435966 57922 436022 57978
rect 439314 598116 439370 598172
rect 439438 598116 439494 598172
rect 439562 598116 439618 598172
rect 439686 598116 439742 598172
rect 439314 597992 439370 598048
rect 439438 597992 439494 598048
rect 439562 597992 439618 598048
rect 439686 597992 439742 598048
rect 439314 597868 439370 597924
rect 439438 597868 439494 597924
rect 439562 597868 439618 597924
rect 439686 597868 439742 597924
rect 439314 597744 439370 597800
rect 439438 597744 439494 597800
rect 439562 597744 439618 597800
rect 439686 597744 439742 597800
rect 439314 586294 439370 586350
rect 439438 586294 439494 586350
rect 439562 586294 439618 586350
rect 439686 586294 439742 586350
rect 439314 586170 439370 586226
rect 439438 586170 439494 586226
rect 439562 586170 439618 586226
rect 439686 586170 439742 586226
rect 439314 586046 439370 586102
rect 439438 586046 439494 586102
rect 439562 586046 439618 586102
rect 439686 586046 439742 586102
rect 439314 585922 439370 585978
rect 439438 585922 439494 585978
rect 439562 585922 439618 585978
rect 439686 585922 439742 585978
rect 439314 568294 439370 568350
rect 439438 568294 439494 568350
rect 439562 568294 439618 568350
rect 439686 568294 439742 568350
rect 439314 568170 439370 568226
rect 439438 568170 439494 568226
rect 439562 568170 439618 568226
rect 439686 568170 439742 568226
rect 439314 568046 439370 568102
rect 439438 568046 439494 568102
rect 439562 568046 439618 568102
rect 439686 568046 439742 568102
rect 439314 567922 439370 567978
rect 439438 567922 439494 567978
rect 439562 567922 439618 567978
rect 439686 567922 439742 567978
rect 439314 550294 439370 550350
rect 439438 550294 439494 550350
rect 439562 550294 439618 550350
rect 439686 550294 439742 550350
rect 439314 550170 439370 550226
rect 439438 550170 439494 550226
rect 439562 550170 439618 550226
rect 439686 550170 439742 550226
rect 439314 550046 439370 550102
rect 439438 550046 439494 550102
rect 439562 550046 439618 550102
rect 439686 550046 439742 550102
rect 439314 549922 439370 549978
rect 439438 549922 439494 549978
rect 439562 549922 439618 549978
rect 439686 549922 439742 549978
rect 439314 532294 439370 532350
rect 439438 532294 439494 532350
rect 439562 532294 439618 532350
rect 439686 532294 439742 532350
rect 439314 532170 439370 532226
rect 439438 532170 439494 532226
rect 439562 532170 439618 532226
rect 439686 532170 439742 532226
rect 439314 532046 439370 532102
rect 439438 532046 439494 532102
rect 439562 532046 439618 532102
rect 439686 532046 439742 532102
rect 439314 531922 439370 531978
rect 439438 531922 439494 531978
rect 439562 531922 439618 531978
rect 439686 531922 439742 531978
rect 439314 514294 439370 514350
rect 439438 514294 439494 514350
rect 439562 514294 439618 514350
rect 439686 514294 439742 514350
rect 439314 514170 439370 514226
rect 439438 514170 439494 514226
rect 439562 514170 439618 514226
rect 439686 514170 439742 514226
rect 439314 514046 439370 514102
rect 439438 514046 439494 514102
rect 439562 514046 439618 514102
rect 439686 514046 439742 514102
rect 439314 513922 439370 513978
rect 439438 513922 439494 513978
rect 439562 513922 439618 513978
rect 439686 513922 439742 513978
rect 439314 496294 439370 496350
rect 439438 496294 439494 496350
rect 439562 496294 439618 496350
rect 439686 496294 439742 496350
rect 439314 496170 439370 496226
rect 439438 496170 439494 496226
rect 439562 496170 439618 496226
rect 439686 496170 439742 496226
rect 439314 496046 439370 496102
rect 439438 496046 439494 496102
rect 439562 496046 439618 496102
rect 439686 496046 439742 496102
rect 439314 495922 439370 495978
rect 439438 495922 439494 495978
rect 439562 495922 439618 495978
rect 439686 495922 439742 495978
rect 439314 478294 439370 478350
rect 439438 478294 439494 478350
rect 439562 478294 439618 478350
rect 439686 478294 439742 478350
rect 439314 478170 439370 478226
rect 439438 478170 439494 478226
rect 439562 478170 439618 478226
rect 439686 478170 439742 478226
rect 439314 478046 439370 478102
rect 439438 478046 439494 478102
rect 439562 478046 439618 478102
rect 439686 478046 439742 478102
rect 439314 477922 439370 477978
rect 439438 477922 439494 477978
rect 439562 477922 439618 477978
rect 439686 477922 439742 477978
rect 439314 460294 439370 460350
rect 439438 460294 439494 460350
rect 439562 460294 439618 460350
rect 439686 460294 439742 460350
rect 439314 460170 439370 460226
rect 439438 460170 439494 460226
rect 439562 460170 439618 460226
rect 439686 460170 439742 460226
rect 439314 460046 439370 460102
rect 439438 460046 439494 460102
rect 439562 460046 439618 460102
rect 439686 460046 439742 460102
rect 439314 459922 439370 459978
rect 439438 459922 439494 459978
rect 439562 459922 439618 459978
rect 439686 459922 439742 459978
rect 439314 442294 439370 442350
rect 439438 442294 439494 442350
rect 439562 442294 439618 442350
rect 439686 442294 439742 442350
rect 439314 442170 439370 442226
rect 439438 442170 439494 442226
rect 439562 442170 439618 442226
rect 439686 442170 439742 442226
rect 439314 442046 439370 442102
rect 439438 442046 439494 442102
rect 439562 442046 439618 442102
rect 439686 442046 439742 442102
rect 439314 441922 439370 441978
rect 439438 441922 439494 441978
rect 439562 441922 439618 441978
rect 439686 441922 439742 441978
rect 439314 424294 439370 424350
rect 439438 424294 439494 424350
rect 439562 424294 439618 424350
rect 439686 424294 439742 424350
rect 439314 424170 439370 424226
rect 439438 424170 439494 424226
rect 439562 424170 439618 424226
rect 439686 424170 439742 424226
rect 439314 424046 439370 424102
rect 439438 424046 439494 424102
rect 439562 424046 439618 424102
rect 439686 424046 439742 424102
rect 439314 423922 439370 423978
rect 439438 423922 439494 423978
rect 439562 423922 439618 423978
rect 439686 423922 439742 423978
rect 439314 406294 439370 406350
rect 439438 406294 439494 406350
rect 439562 406294 439618 406350
rect 439686 406294 439742 406350
rect 439314 406170 439370 406226
rect 439438 406170 439494 406226
rect 439562 406170 439618 406226
rect 439686 406170 439742 406226
rect 439314 406046 439370 406102
rect 439438 406046 439494 406102
rect 439562 406046 439618 406102
rect 439686 406046 439742 406102
rect 439314 405922 439370 405978
rect 439438 405922 439494 405978
rect 439562 405922 439618 405978
rect 439686 405922 439742 405978
rect 439314 388294 439370 388350
rect 439438 388294 439494 388350
rect 439562 388294 439618 388350
rect 439686 388294 439742 388350
rect 439314 388170 439370 388226
rect 439438 388170 439494 388226
rect 439562 388170 439618 388226
rect 439686 388170 439742 388226
rect 439314 388046 439370 388102
rect 439438 388046 439494 388102
rect 439562 388046 439618 388102
rect 439686 388046 439742 388102
rect 439314 387922 439370 387978
rect 439438 387922 439494 387978
rect 439562 387922 439618 387978
rect 439686 387922 439742 387978
rect 439314 370294 439370 370350
rect 439438 370294 439494 370350
rect 439562 370294 439618 370350
rect 439686 370294 439742 370350
rect 439314 370170 439370 370226
rect 439438 370170 439494 370226
rect 439562 370170 439618 370226
rect 439686 370170 439742 370226
rect 439314 370046 439370 370102
rect 439438 370046 439494 370102
rect 439562 370046 439618 370102
rect 439686 370046 439742 370102
rect 439314 369922 439370 369978
rect 439438 369922 439494 369978
rect 439562 369922 439618 369978
rect 439686 369922 439742 369978
rect 439314 352294 439370 352350
rect 439438 352294 439494 352350
rect 439562 352294 439618 352350
rect 439686 352294 439742 352350
rect 439314 352170 439370 352226
rect 439438 352170 439494 352226
rect 439562 352170 439618 352226
rect 439686 352170 439742 352226
rect 439314 352046 439370 352102
rect 439438 352046 439494 352102
rect 439562 352046 439618 352102
rect 439686 352046 439742 352102
rect 439314 351922 439370 351978
rect 439438 351922 439494 351978
rect 439562 351922 439618 351978
rect 439686 351922 439742 351978
rect 439314 334294 439370 334350
rect 439438 334294 439494 334350
rect 439562 334294 439618 334350
rect 439686 334294 439742 334350
rect 439314 334170 439370 334226
rect 439438 334170 439494 334226
rect 439562 334170 439618 334226
rect 439686 334170 439742 334226
rect 439314 334046 439370 334102
rect 439438 334046 439494 334102
rect 439562 334046 439618 334102
rect 439686 334046 439742 334102
rect 439314 333922 439370 333978
rect 439438 333922 439494 333978
rect 439562 333922 439618 333978
rect 439686 333922 439742 333978
rect 439314 316294 439370 316350
rect 439438 316294 439494 316350
rect 439562 316294 439618 316350
rect 439686 316294 439742 316350
rect 439314 316170 439370 316226
rect 439438 316170 439494 316226
rect 439562 316170 439618 316226
rect 439686 316170 439742 316226
rect 439314 316046 439370 316102
rect 439438 316046 439494 316102
rect 439562 316046 439618 316102
rect 439686 316046 439742 316102
rect 439314 315922 439370 315978
rect 439438 315922 439494 315978
rect 439562 315922 439618 315978
rect 439686 315922 439742 315978
rect 439314 298294 439370 298350
rect 439438 298294 439494 298350
rect 439562 298294 439618 298350
rect 439686 298294 439742 298350
rect 439314 298170 439370 298226
rect 439438 298170 439494 298226
rect 439562 298170 439618 298226
rect 439686 298170 439742 298226
rect 439314 298046 439370 298102
rect 439438 298046 439494 298102
rect 439562 298046 439618 298102
rect 439686 298046 439742 298102
rect 439314 297922 439370 297978
rect 439438 297922 439494 297978
rect 439562 297922 439618 297978
rect 439686 297922 439742 297978
rect 439314 280294 439370 280350
rect 439438 280294 439494 280350
rect 439562 280294 439618 280350
rect 439686 280294 439742 280350
rect 439314 280170 439370 280226
rect 439438 280170 439494 280226
rect 439562 280170 439618 280226
rect 439686 280170 439742 280226
rect 439314 280046 439370 280102
rect 439438 280046 439494 280102
rect 439562 280046 439618 280102
rect 439686 280046 439742 280102
rect 439314 279922 439370 279978
rect 439438 279922 439494 279978
rect 439562 279922 439618 279978
rect 439686 279922 439742 279978
rect 439314 262294 439370 262350
rect 439438 262294 439494 262350
rect 439562 262294 439618 262350
rect 439686 262294 439742 262350
rect 439314 262170 439370 262226
rect 439438 262170 439494 262226
rect 439562 262170 439618 262226
rect 439686 262170 439742 262226
rect 439314 262046 439370 262102
rect 439438 262046 439494 262102
rect 439562 262046 439618 262102
rect 439686 262046 439742 262102
rect 439314 261922 439370 261978
rect 439438 261922 439494 261978
rect 439562 261922 439618 261978
rect 439686 261922 439742 261978
rect 439314 244294 439370 244350
rect 439438 244294 439494 244350
rect 439562 244294 439618 244350
rect 439686 244294 439742 244350
rect 439314 244170 439370 244226
rect 439438 244170 439494 244226
rect 439562 244170 439618 244226
rect 439686 244170 439742 244226
rect 439314 244046 439370 244102
rect 439438 244046 439494 244102
rect 439562 244046 439618 244102
rect 439686 244046 439742 244102
rect 439314 243922 439370 243978
rect 439438 243922 439494 243978
rect 439562 243922 439618 243978
rect 439686 243922 439742 243978
rect 439314 226294 439370 226350
rect 439438 226294 439494 226350
rect 439562 226294 439618 226350
rect 439686 226294 439742 226350
rect 439314 226170 439370 226226
rect 439438 226170 439494 226226
rect 439562 226170 439618 226226
rect 439686 226170 439742 226226
rect 439314 226046 439370 226102
rect 439438 226046 439494 226102
rect 439562 226046 439618 226102
rect 439686 226046 439742 226102
rect 439314 225922 439370 225978
rect 439438 225922 439494 225978
rect 439562 225922 439618 225978
rect 439686 225922 439742 225978
rect 439314 208294 439370 208350
rect 439438 208294 439494 208350
rect 439562 208294 439618 208350
rect 439686 208294 439742 208350
rect 439314 208170 439370 208226
rect 439438 208170 439494 208226
rect 439562 208170 439618 208226
rect 439686 208170 439742 208226
rect 439314 208046 439370 208102
rect 439438 208046 439494 208102
rect 439562 208046 439618 208102
rect 439686 208046 439742 208102
rect 439314 207922 439370 207978
rect 439438 207922 439494 207978
rect 439562 207922 439618 207978
rect 439686 207922 439742 207978
rect 439314 190294 439370 190350
rect 439438 190294 439494 190350
rect 439562 190294 439618 190350
rect 439686 190294 439742 190350
rect 439314 190170 439370 190226
rect 439438 190170 439494 190226
rect 439562 190170 439618 190226
rect 439686 190170 439742 190226
rect 439314 190046 439370 190102
rect 439438 190046 439494 190102
rect 439562 190046 439618 190102
rect 439686 190046 439742 190102
rect 439314 189922 439370 189978
rect 439438 189922 439494 189978
rect 439562 189922 439618 189978
rect 439686 189922 439742 189978
rect 439314 172294 439370 172350
rect 439438 172294 439494 172350
rect 439562 172294 439618 172350
rect 439686 172294 439742 172350
rect 439314 172170 439370 172226
rect 439438 172170 439494 172226
rect 439562 172170 439618 172226
rect 439686 172170 439742 172226
rect 439314 172046 439370 172102
rect 439438 172046 439494 172102
rect 439562 172046 439618 172102
rect 439686 172046 439742 172102
rect 439314 171922 439370 171978
rect 439438 171922 439494 171978
rect 439562 171922 439618 171978
rect 439686 171922 439742 171978
rect 439314 154294 439370 154350
rect 439438 154294 439494 154350
rect 439562 154294 439618 154350
rect 439686 154294 439742 154350
rect 439314 154170 439370 154226
rect 439438 154170 439494 154226
rect 439562 154170 439618 154226
rect 439686 154170 439742 154226
rect 439314 154046 439370 154102
rect 439438 154046 439494 154102
rect 439562 154046 439618 154102
rect 439686 154046 439742 154102
rect 439314 153922 439370 153978
rect 439438 153922 439494 153978
rect 439562 153922 439618 153978
rect 439686 153922 439742 153978
rect 439314 136294 439370 136350
rect 439438 136294 439494 136350
rect 439562 136294 439618 136350
rect 439686 136294 439742 136350
rect 439314 136170 439370 136226
rect 439438 136170 439494 136226
rect 439562 136170 439618 136226
rect 439686 136170 439742 136226
rect 439314 136046 439370 136102
rect 439438 136046 439494 136102
rect 439562 136046 439618 136102
rect 439686 136046 439742 136102
rect 439314 135922 439370 135978
rect 439438 135922 439494 135978
rect 439562 135922 439618 135978
rect 439686 135922 439742 135978
rect 439314 118294 439370 118350
rect 439438 118294 439494 118350
rect 439562 118294 439618 118350
rect 439686 118294 439742 118350
rect 439314 118170 439370 118226
rect 439438 118170 439494 118226
rect 439562 118170 439618 118226
rect 439686 118170 439742 118226
rect 439314 118046 439370 118102
rect 439438 118046 439494 118102
rect 439562 118046 439618 118102
rect 439686 118046 439742 118102
rect 439314 117922 439370 117978
rect 439438 117922 439494 117978
rect 439562 117922 439618 117978
rect 439686 117922 439742 117978
rect 439314 100294 439370 100350
rect 439438 100294 439494 100350
rect 439562 100294 439618 100350
rect 439686 100294 439742 100350
rect 439314 100170 439370 100226
rect 439438 100170 439494 100226
rect 439562 100170 439618 100226
rect 439686 100170 439742 100226
rect 439314 100046 439370 100102
rect 439438 100046 439494 100102
rect 439562 100046 439618 100102
rect 439686 100046 439742 100102
rect 439314 99922 439370 99978
rect 439438 99922 439494 99978
rect 439562 99922 439618 99978
rect 439686 99922 439742 99978
rect 439314 82294 439370 82350
rect 439438 82294 439494 82350
rect 439562 82294 439618 82350
rect 439686 82294 439742 82350
rect 439314 82170 439370 82226
rect 439438 82170 439494 82226
rect 439562 82170 439618 82226
rect 439686 82170 439742 82226
rect 439314 82046 439370 82102
rect 439438 82046 439494 82102
rect 439562 82046 439618 82102
rect 439686 82046 439742 82102
rect 439314 81922 439370 81978
rect 439438 81922 439494 81978
rect 439562 81922 439618 81978
rect 439686 81922 439742 81978
rect 466314 597156 466370 597212
rect 466438 597156 466494 597212
rect 466562 597156 466618 597212
rect 466686 597156 466742 597212
rect 466314 597032 466370 597088
rect 466438 597032 466494 597088
rect 466562 597032 466618 597088
rect 466686 597032 466742 597088
rect 466314 596908 466370 596964
rect 466438 596908 466494 596964
rect 466562 596908 466618 596964
rect 466686 596908 466742 596964
rect 466314 596784 466370 596840
rect 466438 596784 466494 596840
rect 466562 596784 466618 596840
rect 466686 596784 466742 596840
rect 466314 580294 466370 580350
rect 466438 580294 466494 580350
rect 466562 580294 466618 580350
rect 466686 580294 466742 580350
rect 466314 580170 466370 580226
rect 466438 580170 466494 580226
rect 466562 580170 466618 580226
rect 466686 580170 466742 580226
rect 466314 580046 466370 580102
rect 466438 580046 466494 580102
rect 466562 580046 466618 580102
rect 466686 580046 466742 580102
rect 466314 579922 466370 579978
rect 466438 579922 466494 579978
rect 466562 579922 466618 579978
rect 466686 579922 466742 579978
rect 466314 562294 466370 562350
rect 466438 562294 466494 562350
rect 466562 562294 466618 562350
rect 466686 562294 466742 562350
rect 466314 562170 466370 562226
rect 466438 562170 466494 562226
rect 466562 562170 466618 562226
rect 466686 562170 466742 562226
rect 466314 562046 466370 562102
rect 466438 562046 466494 562102
rect 466562 562046 466618 562102
rect 466686 562046 466742 562102
rect 466314 561922 466370 561978
rect 466438 561922 466494 561978
rect 466562 561922 466618 561978
rect 466686 561922 466742 561978
rect 466314 544294 466370 544350
rect 466438 544294 466494 544350
rect 466562 544294 466618 544350
rect 466686 544294 466742 544350
rect 466314 544170 466370 544226
rect 466438 544170 466494 544226
rect 466562 544170 466618 544226
rect 466686 544170 466742 544226
rect 466314 544046 466370 544102
rect 466438 544046 466494 544102
rect 466562 544046 466618 544102
rect 466686 544046 466742 544102
rect 466314 543922 466370 543978
rect 466438 543922 466494 543978
rect 466562 543922 466618 543978
rect 466686 543922 466742 543978
rect 466314 526294 466370 526350
rect 466438 526294 466494 526350
rect 466562 526294 466618 526350
rect 466686 526294 466742 526350
rect 466314 526170 466370 526226
rect 466438 526170 466494 526226
rect 466562 526170 466618 526226
rect 466686 526170 466742 526226
rect 466314 526046 466370 526102
rect 466438 526046 466494 526102
rect 466562 526046 466618 526102
rect 466686 526046 466742 526102
rect 466314 525922 466370 525978
rect 466438 525922 466494 525978
rect 466562 525922 466618 525978
rect 466686 525922 466742 525978
rect 466314 508294 466370 508350
rect 466438 508294 466494 508350
rect 466562 508294 466618 508350
rect 466686 508294 466742 508350
rect 466314 508170 466370 508226
rect 466438 508170 466494 508226
rect 466562 508170 466618 508226
rect 466686 508170 466742 508226
rect 466314 508046 466370 508102
rect 466438 508046 466494 508102
rect 466562 508046 466618 508102
rect 466686 508046 466742 508102
rect 466314 507922 466370 507978
rect 466438 507922 466494 507978
rect 466562 507922 466618 507978
rect 466686 507922 466742 507978
rect 466314 490294 466370 490350
rect 466438 490294 466494 490350
rect 466562 490294 466618 490350
rect 466686 490294 466742 490350
rect 466314 490170 466370 490226
rect 466438 490170 466494 490226
rect 466562 490170 466618 490226
rect 466686 490170 466742 490226
rect 466314 490046 466370 490102
rect 466438 490046 466494 490102
rect 466562 490046 466618 490102
rect 466686 490046 466742 490102
rect 466314 489922 466370 489978
rect 466438 489922 466494 489978
rect 466562 489922 466618 489978
rect 466686 489922 466742 489978
rect 466314 472294 466370 472350
rect 466438 472294 466494 472350
rect 466562 472294 466618 472350
rect 466686 472294 466742 472350
rect 466314 472170 466370 472226
rect 466438 472170 466494 472226
rect 466562 472170 466618 472226
rect 466686 472170 466742 472226
rect 466314 472046 466370 472102
rect 466438 472046 466494 472102
rect 466562 472046 466618 472102
rect 466686 472046 466742 472102
rect 466314 471922 466370 471978
rect 466438 471922 466494 471978
rect 466562 471922 466618 471978
rect 466686 471922 466742 471978
rect 466314 454294 466370 454350
rect 466438 454294 466494 454350
rect 466562 454294 466618 454350
rect 466686 454294 466742 454350
rect 466314 454170 466370 454226
rect 466438 454170 466494 454226
rect 466562 454170 466618 454226
rect 466686 454170 466742 454226
rect 466314 454046 466370 454102
rect 466438 454046 466494 454102
rect 466562 454046 466618 454102
rect 466686 454046 466742 454102
rect 466314 453922 466370 453978
rect 466438 453922 466494 453978
rect 466562 453922 466618 453978
rect 466686 453922 466742 453978
rect 466314 436294 466370 436350
rect 466438 436294 466494 436350
rect 466562 436294 466618 436350
rect 466686 436294 466742 436350
rect 466314 436170 466370 436226
rect 466438 436170 466494 436226
rect 466562 436170 466618 436226
rect 466686 436170 466742 436226
rect 466314 436046 466370 436102
rect 466438 436046 466494 436102
rect 466562 436046 466618 436102
rect 466686 436046 466742 436102
rect 466314 435922 466370 435978
rect 466438 435922 466494 435978
rect 466562 435922 466618 435978
rect 466686 435922 466742 435978
rect 466314 418294 466370 418350
rect 466438 418294 466494 418350
rect 466562 418294 466618 418350
rect 466686 418294 466742 418350
rect 466314 418170 466370 418226
rect 466438 418170 466494 418226
rect 466562 418170 466618 418226
rect 466686 418170 466742 418226
rect 466314 418046 466370 418102
rect 466438 418046 466494 418102
rect 466562 418046 466618 418102
rect 466686 418046 466742 418102
rect 466314 417922 466370 417978
rect 466438 417922 466494 417978
rect 466562 417922 466618 417978
rect 466686 417922 466742 417978
rect 466314 400294 466370 400350
rect 466438 400294 466494 400350
rect 466562 400294 466618 400350
rect 466686 400294 466742 400350
rect 466314 400170 466370 400226
rect 466438 400170 466494 400226
rect 466562 400170 466618 400226
rect 466686 400170 466742 400226
rect 466314 400046 466370 400102
rect 466438 400046 466494 400102
rect 466562 400046 466618 400102
rect 466686 400046 466742 400102
rect 466314 399922 466370 399978
rect 466438 399922 466494 399978
rect 466562 399922 466618 399978
rect 466686 399922 466742 399978
rect 466314 382294 466370 382350
rect 466438 382294 466494 382350
rect 466562 382294 466618 382350
rect 466686 382294 466742 382350
rect 466314 382170 466370 382226
rect 466438 382170 466494 382226
rect 466562 382170 466618 382226
rect 466686 382170 466742 382226
rect 466314 382046 466370 382102
rect 466438 382046 466494 382102
rect 466562 382046 466618 382102
rect 466686 382046 466742 382102
rect 466314 381922 466370 381978
rect 466438 381922 466494 381978
rect 466562 381922 466618 381978
rect 466686 381922 466742 381978
rect 466314 364294 466370 364350
rect 466438 364294 466494 364350
rect 466562 364294 466618 364350
rect 466686 364294 466742 364350
rect 466314 364170 466370 364226
rect 466438 364170 466494 364226
rect 466562 364170 466618 364226
rect 466686 364170 466742 364226
rect 466314 364046 466370 364102
rect 466438 364046 466494 364102
rect 466562 364046 466618 364102
rect 466686 364046 466742 364102
rect 466314 363922 466370 363978
rect 466438 363922 466494 363978
rect 466562 363922 466618 363978
rect 466686 363922 466742 363978
rect 466314 346294 466370 346350
rect 466438 346294 466494 346350
rect 466562 346294 466618 346350
rect 466686 346294 466742 346350
rect 466314 346170 466370 346226
rect 466438 346170 466494 346226
rect 466562 346170 466618 346226
rect 466686 346170 466742 346226
rect 466314 346046 466370 346102
rect 466438 346046 466494 346102
rect 466562 346046 466618 346102
rect 466686 346046 466742 346102
rect 466314 345922 466370 345978
rect 466438 345922 466494 345978
rect 466562 345922 466618 345978
rect 466686 345922 466742 345978
rect 466314 328294 466370 328350
rect 466438 328294 466494 328350
rect 466562 328294 466618 328350
rect 466686 328294 466742 328350
rect 466314 328170 466370 328226
rect 466438 328170 466494 328226
rect 466562 328170 466618 328226
rect 466686 328170 466742 328226
rect 466314 328046 466370 328102
rect 466438 328046 466494 328102
rect 466562 328046 466618 328102
rect 466686 328046 466742 328102
rect 466314 327922 466370 327978
rect 466438 327922 466494 327978
rect 466562 327922 466618 327978
rect 466686 327922 466742 327978
rect 466314 310294 466370 310350
rect 466438 310294 466494 310350
rect 466562 310294 466618 310350
rect 466686 310294 466742 310350
rect 466314 310170 466370 310226
rect 466438 310170 466494 310226
rect 466562 310170 466618 310226
rect 466686 310170 466742 310226
rect 466314 310046 466370 310102
rect 466438 310046 466494 310102
rect 466562 310046 466618 310102
rect 466686 310046 466742 310102
rect 466314 309922 466370 309978
rect 466438 309922 466494 309978
rect 466562 309922 466618 309978
rect 466686 309922 466742 309978
rect 466314 292294 466370 292350
rect 466438 292294 466494 292350
rect 466562 292294 466618 292350
rect 466686 292294 466742 292350
rect 466314 292170 466370 292226
rect 466438 292170 466494 292226
rect 466562 292170 466618 292226
rect 466686 292170 466742 292226
rect 466314 292046 466370 292102
rect 466438 292046 466494 292102
rect 466562 292046 466618 292102
rect 466686 292046 466742 292102
rect 466314 291922 466370 291978
rect 466438 291922 466494 291978
rect 466562 291922 466618 291978
rect 466686 291922 466742 291978
rect 466314 274294 466370 274350
rect 466438 274294 466494 274350
rect 466562 274294 466618 274350
rect 466686 274294 466742 274350
rect 466314 274170 466370 274226
rect 466438 274170 466494 274226
rect 466562 274170 466618 274226
rect 466686 274170 466742 274226
rect 466314 274046 466370 274102
rect 466438 274046 466494 274102
rect 466562 274046 466618 274102
rect 466686 274046 466742 274102
rect 466314 273922 466370 273978
rect 466438 273922 466494 273978
rect 466562 273922 466618 273978
rect 466686 273922 466742 273978
rect 466314 256294 466370 256350
rect 466438 256294 466494 256350
rect 466562 256294 466618 256350
rect 466686 256294 466742 256350
rect 466314 256170 466370 256226
rect 466438 256170 466494 256226
rect 466562 256170 466618 256226
rect 466686 256170 466742 256226
rect 466314 256046 466370 256102
rect 466438 256046 466494 256102
rect 466562 256046 466618 256102
rect 466686 256046 466742 256102
rect 466314 255922 466370 255978
rect 466438 255922 466494 255978
rect 466562 255922 466618 255978
rect 466686 255922 466742 255978
rect 466314 238294 466370 238350
rect 466438 238294 466494 238350
rect 466562 238294 466618 238350
rect 466686 238294 466742 238350
rect 466314 238170 466370 238226
rect 466438 238170 466494 238226
rect 466562 238170 466618 238226
rect 466686 238170 466742 238226
rect 466314 238046 466370 238102
rect 466438 238046 466494 238102
rect 466562 238046 466618 238102
rect 466686 238046 466742 238102
rect 466314 237922 466370 237978
rect 466438 237922 466494 237978
rect 466562 237922 466618 237978
rect 466686 237922 466742 237978
rect 466314 220294 466370 220350
rect 466438 220294 466494 220350
rect 466562 220294 466618 220350
rect 466686 220294 466742 220350
rect 466314 220170 466370 220226
rect 466438 220170 466494 220226
rect 466562 220170 466618 220226
rect 466686 220170 466742 220226
rect 466314 220046 466370 220102
rect 466438 220046 466494 220102
rect 466562 220046 466618 220102
rect 466686 220046 466742 220102
rect 466314 219922 466370 219978
rect 466438 219922 466494 219978
rect 466562 219922 466618 219978
rect 466686 219922 466742 219978
rect 466314 202294 466370 202350
rect 466438 202294 466494 202350
rect 466562 202294 466618 202350
rect 466686 202294 466742 202350
rect 466314 202170 466370 202226
rect 466438 202170 466494 202226
rect 466562 202170 466618 202226
rect 466686 202170 466742 202226
rect 466314 202046 466370 202102
rect 466438 202046 466494 202102
rect 466562 202046 466618 202102
rect 466686 202046 466742 202102
rect 466314 201922 466370 201978
rect 466438 201922 466494 201978
rect 466562 201922 466618 201978
rect 466686 201922 466742 201978
rect 466314 184294 466370 184350
rect 466438 184294 466494 184350
rect 466562 184294 466618 184350
rect 466686 184294 466742 184350
rect 466314 184170 466370 184226
rect 466438 184170 466494 184226
rect 466562 184170 466618 184226
rect 466686 184170 466742 184226
rect 466314 184046 466370 184102
rect 466438 184046 466494 184102
rect 466562 184046 466618 184102
rect 466686 184046 466742 184102
rect 466314 183922 466370 183978
rect 466438 183922 466494 183978
rect 466562 183922 466618 183978
rect 466686 183922 466742 183978
rect 466314 166294 466370 166350
rect 466438 166294 466494 166350
rect 466562 166294 466618 166350
rect 466686 166294 466742 166350
rect 466314 166170 466370 166226
rect 466438 166170 466494 166226
rect 466562 166170 466618 166226
rect 466686 166170 466742 166226
rect 466314 166046 466370 166102
rect 466438 166046 466494 166102
rect 466562 166046 466618 166102
rect 466686 166046 466742 166102
rect 466314 165922 466370 165978
rect 466438 165922 466494 165978
rect 466562 165922 466618 165978
rect 466686 165922 466742 165978
rect 466314 148294 466370 148350
rect 466438 148294 466494 148350
rect 466562 148294 466618 148350
rect 466686 148294 466742 148350
rect 466314 148170 466370 148226
rect 466438 148170 466494 148226
rect 466562 148170 466618 148226
rect 466686 148170 466742 148226
rect 466314 148046 466370 148102
rect 466438 148046 466494 148102
rect 466562 148046 466618 148102
rect 466686 148046 466742 148102
rect 466314 147922 466370 147978
rect 466438 147922 466494 147978
rect 466562 147922 466618 147978
rect 466686 147922 466742 147978
rect 466314 130294 466370 130350
rect 466438 130294 466494 130350
rect 466562 130294 466618 130350
rect 466686 130294 466742 130350
rect 466314 130170 466370 130226
rect 466438 130170 466494 130226
rect 466562 130170 466618 130226
rect 466686 130170 466742 130226
rect 466314 130046 466370 130102
rect 466438 130046 466494 130102
rect 466562 130046 466618 130102
rect 466686 130046 466742 130102
rect 466314 129922 466370 129978
rect 466438 129922 466494 129978
rect 466562 129922 466618 129978
rect 466686 129922 466742 129978
rect 466314 112294 466370 112350
rect 466438 112294 466494 112350
rect 466562 112294 466618 112350
rect 466686 112294 466742 112350
rect 466314 112170 466370 112226
rect 466438 112170 466494 112226
rect 466562 112170 466618 112226
rect 466686 112170 466742 112226
rect 466314 112046 466370 112102
rect 466438 112046 466494 112102
rect 466562 112046 466618 112102
rect 466686 112046 466742 112102
rect 466314 111922 466370 111978
rect 466438 111922 466494 111978
rect 466562 111922 466618 111978
rect 466686 111922 466742 111978
rect 466314 94294 466370 94350
rect 466438 94294 466494 94350
rect 466562 94294 466618 94350
rect 466686 94294 466742 94350
rect 466314 94170 466370 94226
rect 466438 94170 466494 94226
rect 466562 94170 466618 94226
rect 466686 94170 466742 94226
rect 466314 94046 466370 94102
rect 466438 94046 466494 94102
rect 466562 94046 466618 94102
rect 466686 94046 466742 94102
rect 466314 93922 466370 93978
rect 466438 93922 466494 93978
rect 466562 93922 466618 93978
rect 466686 93922 466742 93978
rect 439314 64294 439370 64350
rect 439438 64294 439494 64350
rect 439562 64294 439618 64350
rect 439686 64294 439742 64350
rect 439314 64170 439370 64226
rect 439438 64170 439494 64226
rect 439562 64170 439618 64226
rect 439686 64170 439742 64226
rect 439314 64046 439370 64102
rect 439438 64046 439494 64102
rect 439562 64046 439618 64102
rect 439686 64046 439742 64102
rect 439314 63922 439370 63978
rect 439438 63922 439494 63978
rect 439562 63922 439618 63978
rect 439686 63922 439742 63978
rect 435594 40294 435650 40350
rect 435718 40294 435774 40350
rect 435842 40294 435898 40350
rect 435966 40294 436022 40350
rect 435594 40170 435650 40226
rect 435718 40170 435774 40226
rect 435842 40170 435898 40226
rect 435966 40170 436022 40226
rect 435594 40046 435650 40102
rect 435718 40046 435774 40102
rect 435842 40046 435898 40102
rect 435966 40046 436022 40102
rect 435594 39922 435650 39978
rect 435718 39922 435774 39978
rect 435842 39922 435898 39978
rect 435966 39922 436022 39978
rect 435594 22294 435650 22350
rect 435718 22294 435774 22350
rect 435842 22294 435898 22350
rect 435966 22294 436022 22350
rect 435594 22170 435650 22226
rect 435718 22170 435774 22226
rect 435842 22170 435898 22226
rect 435966 22170 436022 22226
rect 435594 22046 435650 22102
rect 435718 22046 435774 22102
rect 435842 22046 435898 22102
rect 435966 22046 436022 22102
rect 435594 21922 435650 21978
rect 435718 21922 435774 21978
rect 435842 21922 435898 21978
rect 435966 21922 436022 21978
rect 435594 4294 435650 4350
rect 435718 4294 435774 4350
rect 435842 4294 435898 4350
rect 435966 4294 436022 4350
rect 435594 4170 435650 4226
rect 435718 4170 435774 4226
rect 435842 4170 435898 4226
rect 435966 4170 436022 4226
rect 436828 51002 436884 51058
rect 446908 79262 446964 79318
rect 439314 46294 439370 46350
rect 439438 46294 439494 46350
rect 439562 46294 439618 46350
rect 439686 46294 439742 46350
rect 439314 46170 439370 46226
rect 439438 46170 439494 46226
rect 439562 46170 439618 46226
rect 439686 46170 439742 46226
rect 439314 46046 439370 46102
rect 439438 46046 439494 46102
rect 439562 46046 439618 46102
rect 439686 46046 439742 46102
rect 439314 45922 439370 45978
rect 439438 45922 439494 45978
rect 439562 45922 439618 45978
rect 439686 45922 439742 45978
rect 439314 28294 439370 28350
rect 439438 28294 439494 28350
rect 439562 28294 439618 28350
rect 439686 28294 439742 28350
rect 439314 28170 439370 28226
rect 439438 28170 439494 28226
rect 439562 28170 439618 28226
rect 439686 28170 439742 28226
rect 439314 28046 439370 28102
rect 439438 28046 439494 28102
rect 439562 28046 439618 28102
rect 439686 28046 439742 28102
rect 439314 27922 439370 27978
rect 439438 27922 439494 27978
rect 439562 27922 439618 27978
rect 439686 27922 439742 27978
rect 438508 11942 438564 11998
rect 439314 10294 439370 10350
rect 439438 10294 439494 10350
rect 439562 10294 439618 10350
rect 439686 10294 439742 10350
rect 439314 10170 439370 10226
rect 439438 10170 439494 10226
rect 439562 10170 439618 10226
rect 439686 10170 439742 10226
rect 439314 10046 439370 10102
rect 439438 10046 439494 10102
rect 439562 10046 439618 10102
rect 439686 10046 439742 10102
rect 439314 9922 439370 9978
rect 439438 9922 439494 9978
rect 439562 9922 439618 9978
rect 439686 9922 439742 9978
rect 435594 4046 435650 4102
rect 435718 4046 435774 4102
rect 435842 4046 435898 4102
rect 435966 4046 436022 4102
rect 435594 3922 435650 3978
rect 435718 3922 435774 3978
rect 435842 3922 435898 3978
rect 435966 3922 436022 3978
rect 408594 -1176 408650 -1120
rect 408718 -1176 408774 -1120
rect 408842 -1176 408898 -1120
rect 408966 -1176 409022 -1120
rect 408594 -1300 408650 -1244
rect 408718 -1300 408774 -1244
rect 408842 -1300 408898 -1244
rect 408966 -1300 409022 -1244
rect 408594 -1424 408650 -1368
rect 408718 -1424 408774 -1368
rect 408842 -1424 408898 -1368
rect 408966 -1424 409022 -1368
rect 408594 -1548 408650 -1492
rect 408718 -1548 408774 -1492
rect 408842 -1548 408898 -1492
rect 408966 -1548 409022 -1492
rect 435594 -216 435650 -160
rect 435718 -216 435774 -160
rect 435842 -216 435898 -160
rect 435966 -216 436022 -160
rect 435594 -340 435650 -284
rect 435718 -340 435774 -284
rect 435842 -340 435898 -284
rect 435966 -340 436022 -284
rect 435594 -464 435650 -408
rect 435718 -464 435774 -408
rect 435842 -464 435898 -408
rect 435966 -464 436022 -408
rect 435594 -588 435650 -532
rect 435718 -588 435774 -532
rect 435842 -588 435898 -532
rect 435966 -588 436022 -532
rect 443548 49022 443604 49078
rect 466314 76294 466370 76350
rect 466438 76294 466494 76350
rect 466562 76294 466618 76350
rect 466686 76294 466742 76350
rect 466314 76170 466370 76226
rect 466438 76170 466494 76226
rect 466562 76170 466618 76226
rect 466686 76170 466742 76226
rect 466314 76046 466370 76102
rect 466438 76046 466494 76102
rect 466562 76046 466618 76102
rect 466686 76046 466742 76102
rect 466314 75922 466370 75978
rect 466438 75922 466494 75978
rect 466562 75922 466618 75978
rect 466686 75922 466742 75978
rect 451948 74042 452004 74098
rect 448588 47402 448644 47458
rect 450268 22562 450324 22618
rect 458668 59282 458724 59338
rect 453628 54422 453684 54478
rect 470034 598116 470090 598172
rect 470158 598116 470214 598172
rect 470282 598116 470338 598172
rect 470406 598116 470462 598172
rect 470034 597992 470090 598048
rect 470158 597992 470214 598048
rect 470282 597992 470338 598048
rect 470406 597992 470462 598048
rect 470034 597868 470090 597924
rect 470158 597868 470214 597924
rect 470282 597868 470338 597924
rect 470406 597868 470462 597924
rect 470034 597744 470090 597800
rect 470158 597744 470214 597800
rect 470282 597744 470338 597800
rect 470406 597744 470462 597800
rect 470034 586294 470090 586350
rect 470158 586294 470214 586350
rect 470282 586294 470338 586350
rect 470406 586294 470462 586350
rect 470034 586170 470090 586226
rect 470158 586170 470214 586226
rect 470282 586170 470338 586226
rect 470406 586170 470462 586226
rect 470034 586046 470090 586102
rect 470158 586046 470214 586102
rect 470282 586046 470338 586102
rect 470406 586046 470462 586102
rect 470034 585922 470090 585978
rect 470158 585922 470214 585978
rect 470282 585922 470338 585978
rect 470406 585922 470462 585978
rect 470034 568294 470090 568350
rect 470158 568294 470214 568350
rect 470282 568294 470338 568350
rect 470406 568294 470462 568350
rect 470034 568170 470090 568226
rect 470158 568170 470214 568226
rect 470282 568170 470338 568226
rect 470406 568170 470462 568226
rect 470034 568046 470090 568102
rect 470158 568046 470214 568102
rect 470282 568046 470338 568102
rect 470406 568046 470462 568102
rect 470034 567922 470090 567978
rect 470158 567922 470214 567978
rect 470282 567922 470338 567978
rect 470406 567922 470462 567978
rect 470034 550294 470090 550350
rect 470158 550294 470214 550350
rect 470282 550294 470338 550350
rect 470406 550294 470462 550350
rect 470034 550170 470090 550226
rect 470158 550170 470214 550226
rect 470282 550170 470338 550226
rect 470406 550170 470462 550226
rect 470034 550046 470090 550102
rect 470158 550046 470214 550102
rect 470282 550046 470338 550102
rect 470406 550046 470462 550102
rect 470034 549922 470090 549978
rect 470158 549922 470214 549978
rect 470282 549922 470338 549978
rect 470406 549922 470462 549978
rect 470034 532294 470090 532350
rect 470158 532294 470214 532350
rect 470282 532294 470338 532350
rect 470406 532294 470462 532350
rect 470034 532170 470090 532226
rect 470158 532170 470214 532226
rect 470282 532170 470338 532226
rect 470406 532170 470462 532226
rect 470034 532046 470090 532102
rect 470158 532046 470214 532102
rect 470282 532046 470338 532102
rect 470406 532046 470462 532102
rect 470034 531922 470090 531978
rect 470158 531922 470214 531978
rect 470282 531922 470338 531978
rect 470406 531922 470462 531978
rect 470034 514294 470090 514350
rect 470158 514294 470214 514350
rect 470282 514294 470338 514350
rect 470406 514294 470462 514350
rect 470034 514170 470090 514226
rect 470158 514170 470214 514226
rect 470282 514170 470338 514226
rect 470406 514170 470462 514226
rect 470034 514046 470090 514102
rect 470158 514046 470214 514102
rect 470282 514046 470338 514102
rect 470406 514046 470462 514102
rect 470034 513922 470090 513978
rect 470158 513922 470214 513978
rect 470282 513922 470338 513978
rect 470406 513922 470462 513978
rect 470034 496294 470090 496350
rect 470158 496294 470214 496350
rect 470282 496294 470338 496350
rect 470406 496294 470462 496350
rect 470034 496170 470090 496226
rect 470158 496170 470214 496226
rect 470282 496170 470338 496226
rect 470406 496170 470462 496226
rect 470034 496046 470090 496102
rect 470158 496046 470214 496102
rect 470282 496046 470338 496102
rect 470406 496046 470462 496102
rect 470034 495922 470090 495978
rect 470158 495922 470214 495978
rect 470282 495922 470338 495978
rect 470406 495922 470462 495978
rect 470034 478294 470090 478350
rect 470158 478294 470214 478350
rect 470282 478294 470338 478350
rect 470406 478294 470462 478350
rect 470034 478170 470090 478226
rect 470158 478170 470214 478226
rect 470282 478170 470338 478226
rect 470406 478170 470462 478226
rect 470034 478046 470090 478102
rect 470158 478046 470214 478102
rect 470282 478046 470338 478102
rect 470406 478046 470462 478102
rect 470034 477922 470090 477978
rect 470158 477922 470214 477978
rect 470282 477922 470338 477978
rect 470406 477922 470462 477978
rect 470034 460294 470090 460350
rect 470158 460294 470214 460350
rect 470282 460294 470338 460350
rect 470406 460294 470462 460350
rect 470034 460170 470090 460226
rect 470158 460170 470214 460226
rect 470282 460170 470338 460226
rect 470406 460170 470462 460226
rect 470034 460046 470090 460102
rect 470158 460046 470214 460102
rect 470282 460046 470338 460102
rect 470406 460046 470462 460102
rect 470034 459922 470090 459978
rect 470158 459922 470214 459978
rect 470282 459922 470338 459978
rect 470406 459922 470462 459978
rect 470034 442294 470090 442350
rect 470158 442294 470214 442350
rect 470282 442294 470338 442350
rect 470406 442294 470462 442350
rect 470034 442170 470090 442226
rect 470158 442170 470214 442226
rect 470282 442170 470338 442226
rect 470406 442170 470462 442226
rect 470034 442046 470090 442102
rect 470158 442046 470214 442102
rect 470282 442046 470338 442102
rect 470406 442046 470462 442102
rect 470034 441922 470090 441978
rect 470158 441922 470214 441978
rect 470282 441922 470338 441978
rect 470406 441922 470462 441978
rect 470034 424294 470090 424350
rect 470158 424294 470214 424350
rect 470282 424294 470338 424350
rect 470406 424294 470462 424350
rect 470034 424170 470090 424226
rect 470158 424170 470214 424226
rect 470282 424170 470338 424226
rect 470406 424170 470462 424226
rect 470034 424046 470090 424102
rect 470158 424046 470214 424102
rect 470282 424046 470338 424102
rect 470406 424046 470462 424102
rect 470034 423922 470090 423978
rect 470158 423922 470214 423978
rect 470282 423922 470338 423978
rect 470406 423922 470462 423978
rect 470034 406294 470090 406350
rect 470158 406294 470214 406350
rect 470282 406294 470338 406350
rect 470406 406294 470462 406350
rect 470034 406170 470090 406226
rect 470158 406170 470214 406226
rect 470282 406170 470338 406226
rect 470406 406170 470462 406226
rect 470034 406046 470090 406102
rect 470158 406046 470214 406102
rect 470282 406046 470338 406102
rect 470406 406046 470462 406102
rect 470034 405922 470090 405978
rect 470158 405922 470214 405978
rect 470282 405922 470338 405978
rect 470406 405922 470462 405978
rect 470034 388294 470090 388350
rect 470158 388294 470214 388350
rect 470282 388294 470338 388350
rect 470406 388294 470462 388350
rect 470034 388170 470090 388226
rect 470158 388170 470214 388226
rect 470282 388170 470338 388226
rect 470406 388170 470462 388226
rect 470034 388046 470090 388102
rect 470158 388046 470214 388102
rect 470282 388046 470338 388102
rect 470406 388046 470462 388102
rect 470034 387922 470090 387978
rect 470158 387922 470214 387978
rect 470282 387922 470338 387978
rect 470406 387922 470462 387978
rect 470034 370294 470090 370350
rect 470158 370294 470214 370350
rect 470282 370294 470338 370350
rect 470406 370294 470462 370350
rect 470034 370170 470090 370226
rect 470158 370170 470214 370226
rect 470282 370170 470338 370226
rect 470406 370170 470462 370226
rect 470034 370046 470090 370102
rect 470158 370046 470214 370102
rect 470282 370046 470338 370102
rect 470406 370046 470462 370102
rect 470034 369922 470090 369978
rect 470158 369922 470214 369978
rect 470282 369922 470338 369978
rect 470406 369922 470462 369978
rect 470034 352294 470090 352350
rect 470158 352294 470214 352350
rect 470282 352294 470338 352350
rect 470406 352294 470462 352350
rect 470034 352170 470090 352226
rect 470158 352170 470214 352226
rect 470282 352170 470338 352226
rect 470406 352170 470462 352226
rect 470034 352046 470090 352102
rect 470158 352046 470214 352102
rect 470282 352046 470338 352102
rect 470406 352046 470462 352102
rect 470034 351922 470090 351978
rect 470158 351922 470214 351978
rect 470282 351922 470338 351978
rect 470406 351922 470462 351978
rect 470034 334294 470090 334350
rect 470158 334294 470214 334350
rect 470282 334294 470338 334350
rect 470406 334294 470462 334350
rect 470034 334170 470090 334226
rect 470158 334170 470214 334226
rect 470282 334170 470338 334226
rect 470406 334170 470462 334226
rect 470034 334046 470090 334102
rect 470158 334046 470214 334102
rect 470282 334046 470338 334102
rect 470406 334046 470462 334102
rect 470034 333922 470090 333978
rect 470158 333922 470214 333978
rect 470282 333922 470338 333978
rect 470406 333922 470462 333978
rect 470034 316294 470090 316350
rect 470158 316294 470214 316350
rect 470282 316294 470338 316350
rect 470406 316294 470462 316350
rect 470034 316170 470090 316226
rect 470158 316170 470214 316226
rect 470282 316170 470338 316226
rect 470406 316170 470462 316226
rect 470034 316046 470090 316102
rect 470158 316046 470214 316102
rect 470282 316046 470338 316102
rect 470406 316046 470462 316102
rect 470034 315922 470090 315978
rect 470158 315922 470214 315978
rect 470282 315922 470338 315978
rect 470406 315922 470462 315978
rect 470034 298294 470090 298350
rect 470158 298294 470214 298350
rect 470282 298294 470338 298350
rect 470406 298294 470462 298350
rect 470034 298170 470090 298226
rect 470158 298170 470214 298226
rect 470282 298170 470338 298226
rect 470406 298170 470462 298226
rect 470034 298046 470090 298102
rect 470158 298046 470214 298102
rect 470282 298046 470338 298102
rect 470406 298046 470462 298102
rect 470034 297922 470090 297978
rect 470158 297922 470214 297978
rect 470282 297922 470338 297978
rect 470406 297922 470462 297978
rect 470034 280294 470090 280350
rect 470158 280294 470214 280350
rect 470282 280294 470338 280350
rect 470406 280294 470462 280350
rect 470034 280170 470090 280226
rect 470158 280170 470214 280226
rect 470282 280170 470338 280226
rect 470406 280170 470462 280226
rect 470034 280046 470090 280102
rect 470158 280046 470214 280102
rect 470282 280046 470338 280102
rect 470406 280046 470462 280102
rect 470034 279922 470090 279978
rect 470158 279922 470214 279978
rect 470282 279922 470338 279978
rect 470406 279922 470462 279978
rect 470034 262294 470090 262350
rect 470158 262294 470214 262350
rect 470282 262294 470338 262350
rect 470406 262294 470462 262350
rect 470034 262170 470090 262226
rect 470158 262170 470214 262226
rect 470282 262170 470338 262226
rect 470406 262170 470462 262226
rect 470034 262046 470090 262102
rect 470158 262046 470214 262102
rect 470282 262046 470338 262102
rect 470406 262046 470462 262102
rect 470034 261922 470090 261978
rect 470158 261922 470214 261978
rect 470282 261922 470338 261978
rect 470406 261922 470462 261978
rect 470034 244294 470090 244350
rect 470158 244294 470214 244350
rect 470282 244294 470338 244350
rect 470406 244294 470462 244350
rect 470034 244170 470090 244226
rect 470158 244170 470214 244226
rect 470282 244170 470338 244226
rect 470406 244170 470462 244226
rect 470034 244046 470090 244102
rect 470158 244046 470214 244102
rect 470282 244046 470338 244102
rect 470406 244046 470462 244102
rect 470034 243922 470090 243978
rect 470158 243922 470214 243978
rect 470282 243922 470338 243978
rect 470406 243922 470462 243978
rect 470034 226294 470090 226350
rect 470158 226294 470214 226350
rect 470282 226294 470338 226350
rect 470406 226294 470462 226350
rect 470034 226170 470090 226226
rect 470158 226170 470214 226226
rect 470282 226170 470338 226226
rect 470406 226170 470462 226226
rect 470034 226046 470090 226102
rect 470158 226046 470214 226102
rect 470282 226046 470338 226102
rect 470406 226046 470462 226102
rect 470034 225922 470090 225978
rect 470158 225922 470214 225978
rect 470282 225922 470338 225978
rect 470406 225922 470462 225978
rect 470034 208294 470090 208350
rect 470158 208294 470214 208350
rect 470282 208294 470338 208350
rect 470406 208294 470462 208350
rect 470034 208170 470090 208226
rect 470158 208170 470214 208226
rect 470282 208170 470338 208226
rect 470406 208170 470462 208226
rect 470034 208046 470090 208102
rect 470158 208046 470214 208102
rect 470282 208046 470338 208102
rect 470406 208046 470462 208102
rect 470034 207922 470090 207978
rect 470158 207922 470214 207978
rect 470282 207922 470338 207978
rect 470406 207922 470462 207978
rect 470034 190294 470090 190350
rect 470158 190294 470214 190350
rect 470282 190294 470338 190350
rect 470406 190294 470462 190350
rect 470034 190170 470090 190226
rect 470158 190170 470214 190226
rect 470282 190170 470338 190226
rect 470406 190170 470462 190226
rect 470034 190046 470090 190102
rect 470158 190046 470214 190102
rect 470282 190046 470338 190102
rect 470406 190046 470462 190102
rect 470034 189922 470090 189978
rect 470158 189922 470214 189978
rect 470282 189922 470338 189978
rect 470406 189922 470462 189978
rect 470034 172294 470090 172350
rect 470158 172294 470214 172350
rect 470282 172294 470338 172350
rect 470406 172294 470462 172350
rect 470034 172170 470090 172226
rect 470158 172170 470214 172226
rect 470282 172170 470338 172226
rect 470406 172170 470462 172226
rect 470034 172046 470090 172102
rect 470158 172046 470214 172102
rect 470282 172046 470338 172102
rect 470406 172046 470462 172102
rect 470034 171922 470090 171978
rect 470158 171922 470214 171978
rect 470282 171922 470338 171978
rect 470406 171922 470462 171978
rect 470034 154294 470090 154350
rect 470158 154294 470214 154350
rect 470282 154294 470338 154350
rect 470406 154294 470462 154350
rect 470034 154170 470090 154226
rect 470158 154170 470214 154226
rect 470282 154170 470338 154226
rect 470406 154170 470462 154226
rect 470034 154046 470090 154102
rect 470158 154046 470214 154102
rect 470282 154046 470338 154102
rect 470406 154046 470462 154102
rect 470034 153922 470090 153978
rect 470158 153922 470214 153978
rect 470282 153922 470338 153978
rect 470406 153922 470462 153978
rect 470034 136294 470090 136350
rect 470158 136294 470214 136350
rect 470282 136294 470338 136350
rect 470406 136294 470462 136350
rect 470034 136170 470090 136226
rect 470158 136170 470214 136226
rect 470282 136170 470338 136226
rect 470406 136170 470462 136226
rect 470034 136046 470090 136102
rect 470158 136046 470214 136102
rect 470282 136046 470338 136102
rect 470406 136046 470462 136102
rect 470034 135922 470090 135978
rect 470158 135922 470214 135978
rect 470282 135922 470338 135978
rect 470406 135922 470462 135978
rect 470034 118294 470090 118350
rect 470158 118294 470214 118350
rect 470282 118294 470338 118350
rect 470406 118294 470462 118350
rect 470034 118170 470090 118226
rect 470158 118170 470214 118226
rect 470282 118170 470338 118226
rect 470406 118170 470462 118226
rect 470034 118046 470090 118102
rect 470158 118046 470214 118102
rect 470282 118046 470338 118102
rect 470406 118046 470462 118102
rect 470034 117922 470090 117978
rect 470158 117922 470214 117978
rect 470282 117922 470338 117978
rect 470406 117922 470462 117978
rect 470034 100294 470090 100350
rect 470158 100294 470214 100350
rect 470282 100294 470338 100350
rect 470406 100294 470462 100350
rect 470034 100170 470090 100226
rect 470158 100170 470214 100226
rect 470282 100170 470338 100226
rect 470406 100170 470462 100226
rect 470034 100046 470090 100102
rect 470158 100046 470214 100102
rect 470282 100046 470338 100102
rect 470406 100046 470462 100102
rect 470034 99922 470090 99978
rect 470158 99922 470214 99978
rect 470282 99922 470338 99978
rect 470406 99922 470462 99978
rect 497034 597156 497090 597212
rect 497158 597156 497214 597212
rect 497282 597156 497338 597212
rect 497406 597156 497462 597212
rect 497034 597032 497090 597088
rect 497158 597032 497214 597088
rect 497282 597032 497338 597088
rect 497406 597032 497462 597088
rect 497034 596908 497090 596964
rect 497158 596908 497214 596964
rect 497282 596908 497338 596964
rect 497406 596908 497462 596964
rect 497034 596784 497090 596840
rect 497158 596784 497214 596840
rect 497282 596784 497338 596840
rect 497406 596784 497462 596840
rect 497034 580294 497090 580350
rect 497158 580294 497214 580350
rect 497282 580294 497338 580350
rect 497406 580294 497462 580350
rect 497034 580170 497090 580226
rect 497158 580170 497214 580226
rect 497282 580170 497338 580226
rect 497406 580170 497462 580226
rect 497034 580046 497090 580102
rect 497158 580046 497214 580102
rect 497282 580046 497338 580102
rect 497406 580046 497462 580102
rect 497034 579922 497090 579978
rect 497158 579922 497214 579978
rect 497282 579922 497338 579978
rect 497406 579922 497462 579978
rect 497034 562294 497090 562350
rect 497158 562294 497214 562350
rect 497282 562294 497338 562350
rect 497406 562294 497462 562350
rect 497034 562170 497090 562226
rect 497158 562170 497214 562226
rect 497282 562170 497338 562226
rect 497406 562170 497462 562226
rect 497034 562046 497090 562102
rect 497158 562046 497214 562102
rect 497282 562046 497338 562102
rect 497406 562046 497462 562102
rect 497034 561922 497090 561978
rect 497158 561922 497214 561978
rect 497282 561922 497338 561978
rect 497406 561922 497462 561978
rect 497034 544294 497090 544350
rect 497158 544294 497214 544350
rect 497282 544294 497338 544350
rect 497406 544294 497462 544350
rect 497034 544170 497090 544226
rect 497158 544170 497214 544226
rect 497282 544170 497338 544226
rect 497406 544170 497462 544226
rect 497034 544046 497090 544102
rect 497158 544046 497214 544102
rect 497282 544046 497338 544102
rect 497406 544046 497462 544102
rect 497034 543922 497090 543978
rect 497158 543922 497214 543978
rect 497282 543922 497338 543978
rect 497406 543922 497462 543978
rect 497034 526294 497090 526350
rect 497158 526294 497214 526350
rect 497282 526294 497338 526350
rect 497406 526294 497462 526350
rect 497034 526170 497090 526226
rect 497158 526170 497214 526226
rect 497282 526170 497338 526226
rect 497406 526170 497462 526226
rect 497034 526046 497090 526102
rect 497158 526046 497214 526102
rect 497282 526046 497338 526102
rect 497406 526046 497462 526102
rect 497034 525922 497090 525978
rect 497158 525922 497214 525978
rect 497282 525922 497338 525978
rect 497406 525922 497462 525978
rect 497034 508294 497090 508350
rect 497158 508294 497214 508350
rect 497282 508294 497338 508350
rect 497406 508294 497462 508350
rect 497034 508170 497090 508226
rect 497158 508170 497214 508226
rect 497282 508170 497338 508226
rect 497406 508170 497462 508226
rect 497034 508046 497090 508102
rect 497158 508046 497214 508102
rect 497282 508046 497338 508102
rect 497406 508046 497462 508102
rect 497034 507922 497090 507978
rect 497158 507922 497214 507978
rect 497282 507922 497338 507978
rect 497406 507922 497462 507978
rect 497034 490294 497090 490350
rect 497158 490294 497214 490350
rect 497282 490294 497338 490350
rect 497406 490294 497462 490350
rect 497034 490170 497090 490226
rect 497158 490170 497214 490226
rect 497282 490170 497338 490226
rect 497406 490170 497462 490226
rect 497034 490046 497090 490102
rect 497158 490046 497214 490102
rect 497282 490046 497338 490102
rect 497406 490046 497462 490102
rect 497034 489922 497090 489978
rect 497158 489922 497214 489978
rect 497282 489922 497338 489978
rect 497406 489922 497462 489978
rect 497034 472294 497090 472350
rect 497158 472294 497214 472350
rect 497282 472294 497338 472350
rect 497406 472294 497462 472350
rect 497034 472170 497090 472226
rect 497158 472170 497214 472226
rect 497282 472170 497338 472226
rect 497406 472170 497462 472226
rect 497034 472046 497090 472102
rect 497158 472046 497214 472102
rect 497282 472046 497338 472102
rect 497406 472046 497462 472102
rect 497034 471922 497090 471978
rect 497158 471922 497214 471978
rect 497282 471922 497338 471978
rect 497406 471922 497462 471978
rect 497034 454294 497090 454350
rect 497158 454294 497214 454350
rect 497282 454294 497338 454350
rect 497406 454294 497462 454350
rect 497034 454170 497090 454226
rect 497158 454170 497214 454226
rect 497282 454170 497338 454226
rect 497406 454170 497462 454226
rect 497034 454046 497090 454102
rect 497158 454046 497214 454102
rect 497282 454046 497338 454102
rect 497406 454046 497462 454102
rect 497034 453922 497090 453978
rect 497158 453922 497214 453978
rect 497282 453922 497338 453978
rect 497406 453922 497462 453978
rect 497034 436294 497090 436350
rect 497158 436294 497214 436350
rect 497282 436294 497338 436350
rect 497406 436294 497462 436350
rect 497034 436170 497090 436226
rect 497158 436170 497214 436226
rect 497282 436170 497338 436226
rect 497406 436170 497462 436226
rect 497034 436046 497090 436102
rect 497158 436046 497214 436102
rect 497282 436046 497338 436102
rect 497406 436046 497462 436102
rect 497034 435922 497090 435978
rect 497158 435922 497214 435978
rect 497282 435922 497338 435978
rect 497406 435922 497462 435978
rect 497034 418294 497090 418350
rect 497158 418294 497214 418350
rect 497282 418294 497338 418350
rect 497406 418294 497462 418350
rect 497034 418170 497090 418226
rect 497158 418170 497214 418226
rect 497282 418170 497338 418226
rect 497406 418170 497462 418226
rect 497034 418046 497090 418102
rect 497158 418046 497214 418102
rect 497282 418046 497338 418102
rect 497406 418046 497462 418102
rect 497034 417922 497090 417978
rect 497158 417922 497214 417978
rect 497282 417922 497338 417978
rect 497406 417922 497462 417978
rect 497034 400294 497090 400350
rect 497158 400294 497214 400350
rect 497282 400294 497338 400350
rect 497406 400294 497462 400350
rect 497034 400170 497090 400226
rect 497158 400170 497214 400226
rect 497282 400170 497338 400226
rect 497406 400170 497462 400226
rect 497034 400046 497090 400102
rect 497158 400046 497214 400102
rect 497282 400046 497338 400102
rect 497406 400046 497462 400102
rect 497034 399922 497090 399978
rect 497158 399922 497214 399978
rect 497282 399922 497338 399978
rect 497406 399922 497462 399978
rect 497034 382294 497090 382350
rect 497158 382294 497214 382350
rect 497282 382294 497338 382350
rect 497406 382294 497462 382350
rect 497034 382170 497090 382226
rect 497158 382170 497214 382226
rect 497282 382170 497338 382226
rect 497406 382170 497462 382226
rect 497034 382046 497090 382102
rect 497158 382046 497214 382102
rect 497282 382046 497338 382102
rect 497406 382046 497462 382102
rect 497034 381922 497090 381978
rect 497158 381922 497214 381978
rect 497282 381922 497338 381978
rect 497406 381922 497462 381978
rect 497034 364294 497090 364350
rect 497158 364294 497214 364350
rect 497282 364294 497338 364350
rect 497406 364294 497462 364350
rect 497034 364170 497090 364226
rect 497158 364170 497214 364226
rect 497282 364170 497338 364226
rect 497406 364170 497462 364226
rect 497034 364046 497090 364102
rect 497158 364046 497214 364102
rect 497282 364046 497338 364102
rect 497406 364046 497462 364102
rect 497034 363922 497090 363978
rect 497158 363922 497214 363978
rect 497282 363922 497338 363978
rect 497406 363922 497462 363978
rect 497034 346294 497090 346350
rect 497158 346294 497214 346350
rect 497282 346294 497338 346350
rect 497406 346294 497462 346350
rect 497034 346170 497090 346226
rect 497158 346170 497214 346226
rect 497282 346170 497338 346226
rect 497406 346170 497462 346226
rect 497034 346046 497090 346102
rect 497158 346046 497214 346102
rect 497282 346046 497338 346102
rect 497406 346046 497462 346102
rect 497034 345922 497090 345978
rect 497158 345922 497214 345978
rect 497282 345922 497338 345978
rect 497406 345922 497462 345978
rect 497034 328294 497090 328350
rect 497158 328294 497214 328350
rect 497282 328294 497338 328350
rect 497406 328294 497462 328350
rect 497034 328170 497090 328226
rect 497158 328170 497214 328226
rect 497282 328170 497338 328226
rect 497406 328170 497462 328226
rect 497034 328046 497090 328102
rect 497158 328046 497214 328102
rect 497282 328046 497338 328102
rect 497406 328046 497462 328102
rect 497034 327922 497090 327978
rect 497158 327922 497214 327978
rect 497282 327922 497338 327978
rect 497406 327922 497462 327978
rect 497034 310294 497090 310350
rect 497158 310294 497214 310350
rect 497282 310294 497338 310350
rect 497406 310294 497462 310350
rect 497034 310170 497090 310226
rect 497158 310170 497214 310226
rect 497282 310170 497338 310226
rect 497406 310170 497462 310226
rect 497034 310046 497090 310102
rect 497158 310046 497214 310102
rect 497282 310046 497338 310102
rect 497406 310046 497462 310102
rect 497034 309922 497090 309978
rect 497158 309922 497214 309978
rect 497282 309922 497338 309978
rect 497406 309922 497462 309978
rect 497034 292294 497090 292350
rect 497158 292294 497214 292350
rect 497282 292294 497338 292350
rect 497406 292294 497462 292350
rect 497034 292170 497090 292226
rect 497158 292170 497214 292226
rect 497282 292170 497338 292226
rect 497406 292170 497462 292226
rect 497034 292046 497090 292102
rect 497158 292046 497214 292102
rect 497282 292046 497338 292102
rect 497406 292046 497462 292102
rect 497034 291922 497090 291978
rect 497158 291922 497214 291978
rect 497282 291922 497338 291978
rect 497406 291922 497462 291978
rect 497034 274294 497090 274350
rect 497158 274294 497214 274350
rect 497282 274294 497338 274350
rect 497406 274294 497462 274350
rect 497034 274170 497090 274226
rect 497158 274170 497214 274226
rect 497282 274170 497338 274226
rect 497406 274170 497462 274226
rect 497034 274046 497090 274102
rect 497158 274046 497214 274102
rect 497282 274046 497338 274102
rect 497406 274046 497462 274102
rect 497034 273922 497090 273978
rect 497158 273922 497214 273978
rect 497282 273922 497338 273978
rect 497406 273922 497462 273978
rect 497034 256294 497090 256350
rect 497158 256294 497214 256350
rect 497282 256294 497338 256350
rect 497406 256294 497462 256350
rect 497034 256170 497090 256226
rect 497158 256170 497214 256226
rect 497282 256170 497338 256226
rect 497406 256170 497462 256226
rect 497034 256046 497090 256102
rect 497158 256046 497214 256102
rect 497282 256046 497338 256102
rect 497406 256046 497462 256102
rect 497034 255922 497090 255978
rect 497158 255922 497214 255978
rect 497282 255922 497338 255978
rect 497406 255922 497462 255978
rect 497034 238294 497090 238350
rect 497158 238294 497214 238350
rect 497282 238294 497338 238350
rect 497406 238294 497462 238350
rect 497034 238170 497090 238226
rect 497158 238170 497214 238226
rect 497282 238170 497338 238226
rect 497406 238170 497462 238226
rect 497034 238046 497090 238102
rect 497158 238046 497214 238102
rect 497282 238046 497338 238102
rect 497406 238046 497462 238102
rect 497034 237922 497090 237978
rect 497158 237922 497214 237978
rect 497282 237922 497338 237978
rect 497406 237922 497462 237978
rect 497034 220294 497090 220350
rect 497158 220294 497214 220350
rect 497282 220294 497338 220350
rect 497406 220294 497462 220350
rect 497034 220170 497090 220226
rect 497158 220170 497214 220226
rect 497282 220170 497338 220226
rect 497406 220170 497462 220226
rect 497034 220046 497090 220102
rect 497158 220046 497214 220102
rect 497282 220046 497338 220102
rect 497406 220046 497462 220102
rect 497034 219922 497090 219978
rect 497158 219922 497214 219978
rect 497282 219922 497338 219978
rect 497406 219922 497462 219978
rect 497034 202294 497090 202350
rect 497158 202294 497214 202350
rect 497282 202294 497338 202350
rect 497406 202294 497462 202350
rect 497034 202170 497090 202226
rect 497158 202170 497214 202226
rect 497282 202170 497338 202226
rect 497406 202170 497462 202226
rect 497034 202046 497090 202102
rect 497158 202046 497214 202102
rect 497282 202046 497338 202102
rect 497406 202046 497462 202102
rect 497034 201922 497090 201978
rect 497158 201922 497214 201978
rect 497282 201922 497338 201978
rect 497406 201922 497462 201978
rect 497034 184294 497090 184350
rect 497158 184294 497214 184350
rect 497282 184294 497338 184350
rect 497406 184294 497462 184350
rect 497034 184170 497090 184226
rect 497158 184170 497214 184226
rect 497282 184170 497338 184226
rect 497406 184170 497462 184226
rect 497034 184046 497090 184102
rect 497158 184046 497214 184102
rect 497282 184046 497338 184102
rect 497406 184046 497462 184102
rect 497034 183922 497090 183978
rect 497158 183922 497214 183978
rect 497282 183922 497338 183978
rect 497406 183922 497462 183978
rect 497034 166294 497090 166350
rect 497158 166294 497214 166350
rect 497282 166294 497338 166350
rect 497406 166294 497462 166350
rect 497034 166170 497090 166226
rect 497158 166170 497214 166226
rect 497282 166170 497338 166226
rect 497406 166170 497462 166226
rect 497034 166046 497090 166102
rect 497158 166046 497214 166102
rect 497282 166046 497338 166102
rect 497406 166046 497462 166102
rect 497034 165922 497090 165978
rect 497158 165922 497214 165978
rect 497282 165922 497338 165978
rect 497406 165922 497462 165978
rect 497034 148294 497090 148350
rect 497158 148294 497214 148350
rect 497282 148294 497338 148350
rect 497406 148294 497462 148350
rect 497034 148170 497090 148226
rect 497158 148170 497214 148226
rect 497282 148170 497338 148226
rect 497406 148170 497462 148226
rect 497034 148046 497090 148102
rect 497158 148046 497214 148102
rect 497282 148046 497338 148102
rect 497406 148046 497462 148102
rect 497034 147922 497090 147978
rect 497158 147922 497214 147978
rect 497282 147922 497338 147978
rect 497406 147922 497462 147978
rect 497034 130294 497090 130350
rect 497158 130294 497214 130350
rect 497282 130294 497338 130350
rect 497406 130294 497462 130350
rect 497034 130170 497090 130226
rect 497158 130170 497214 130226
rect 497282 130170 497338 130226
rect 497406 130170 497462 130226
rect 497034 130046 497090 130102
rect 497158 130046 497214 130102
rect 497282 130046 497338 130102
rect 497406 130046 497462 130102
rect 497034 129922 497090 129978
rect 497158 129922 497214 129978
rect 497282 129922 497338 129978
rect 497406 129922 497462 129978
rect 497034 112294 497090 112350
rect 497158 112294 497214 112350
rect 497282 112294 497338 112350
rect 497406 112294 497462 112350
rect 497034 112170 497090 112226
rect 497158 112170 497214 112226
rect 497282 112170 497338 112226
rect 497406 112170 497462 112226
rect 497034 112046 497090 112102
rect 497158 112046 497214 112102
rect 497282 112046 497338 112102
rect 497406 112046 497462 112102
rect 497034 111922 497090 111978
rect 497158 111922 497214 111978
rect 497282 111922 497338 111978
rect 497406 111922 497462 111978
rect 470034 82294 470090 82350
rect 470158 82294 470214 82350
rect 470282 82294 470338 82350
rect 470406 82294 470462 82350
rect 470034 82170 470090 82226
rect 470158 82170 470214 82226
rect 470282 82170 470338 82226
rect 470406 82170 470462 82226
rect 470034 82046 470090 82102
rect 470158 82046 470214 82102
rect 470282 82046 470338 82102
rect 470406 82046 470462 82102
rect 470034 81922 470090 81978
rect 470158 81922 470214 81978
rect 470282 81922 470338 81978
rect 470406 81922 470462 81978
rect 466314 58294 466370 58350
rect 466438 58294 466494 58350
rect 466562 58294 466618 58350
rect 466686 58294 466742 58350
rect 466314 58170 466370 58226
rect 466438 58170 466494 58226
rect 466562 58170 466618 58226
rect 466686 58170 466742 58226
rect 466314 58046 466370 58102
rect 466438 58046 466494 58102
rect 466562 58046 466618 58102
rect 466686 58046 466742 58102
rect 466314 57922 466370 57978
rect 466438 57922 466494 57978
rect 466562 57922 466618 57978
rect 466686 57922 466742 57978
rect 465388 52442 465444 52498
rect 460348 25442 460404 25498
rect 456988 8522 457044 8578
rect 462588 5102 462644 5158
rect 466314 40294 466370 40350
rect 466438 40294 466494 40350
rect 466562 40294 466618 40350
rect 466686 40294 466742 40350
rect 466314 40170 466370 40226
rect 466438 40170 466494 40226
rect 466562 40170 466618 40226
rect 466686 40170 466742 40226
rect 466314 40046 466370 40102
rect 466438 40046 466494 40102
rect 466562 40046 466618 40102
rect 466686 40046 466742 40102
rect 466314 39922 466370 39978
rect 466438 39922 466494 39978
rect 466562 39922 466618 39978
rect 466686 39922 466742 39978
rect 466314 22294 466370 22350
rect 466438 22294 466494 22350
rect 466562 22294 466618 22350
rect 466686 22294 466742 22350
rect 466314 22170 466370 22226
rect 466438 22170 466494 22226
rect 466562 22170 466618 22226
rect 466686 22170 466742 22226
rect 466314 22046 466370 22102
rect 466438 22046 466494 22102
rect 466562 22046 466618 22102
rect 466686 22046 466742 22102
rect 466314 21922 466370 21978
rect 466438 21922 466494 21978
rect 466562 21922 466618 21978
rect 466686 21922 466742 21978
rect 468748 72242 468804 72298
rect 466314 4294 466370 4350
rect 466438 4294 466494 4350
rect 466562 4294 466618 4350
rect 466686 4294 466742 4350
rect 466314 4170 466370 4226
rect 466438 4170 466494 4226
rect 466562 4170 466618 4226
rect 466686 4170 466742 4226
rect 466314 4046 466370 4102
rect 466438 4046 466494 4102
rect 466562 4046 466618 4102
rect 466686 4046 466742 4102
rect 466314 3922 466370 3978
rect 466438 3922 466494 3978
rect 466562 3922 466618 3978
rect 466686 3922 466742 3978
rect 439314 -1176 439370 -1120
rect 439438 -1176 439494 -1120
rect 439562 -1176 439618 -1120
rect 439686 -1176 439742 -1120
rect 439314 -1300 439370 -1244
rect 439438 -1300 439494 -1244
rect 439562 -1300 439618 -1244
rect 439686 -1300 439742 -1244
rect 439314 -1424 439370 -1368
rect 439438 -1424 439494 -1368
rect 439562 -1424 439618 -1368
rect 439686 -1424 439742 -1368
rect 439314 -1548 439370 -1492
rect 439438 -1548 439494 -1492
rect 439562 -1548 439618 -1492
rect 439686 -1548 439742 -1492
rect 468300 6902 468356 6958
rect 470034 64294 470090 64350
rect 470158 64294 470214 64350
rect 470282 64294 470338 64350
rect 470406 64294 470462 64350
rect 470034 64170 470090 64226
rect 470158 64170 470214 64226
rect 470282 64170 470338 64226
rect 470406 64170 470462 64226
rect 470034 64046 470090 64102
rect 470158 64046 470214 64102
rect 470282 64046 470338 64102
rect 470406 64046 470462 64102
rect 470034 63922 470090 63978
rect 470158 63922 470214 63978
rect 470282 63922 470338 63978
rect 470406 63922 470462 63978
rect 470034 46294 470090 46350
rect 470158 46294 470214 46350
rect 470282 46294 470338 46350
rect 470406 46294 470462 46350
rect 470034 46170 470090 46226
rect 470158 46170 470214 46226
rect 470282 46170 470338 46226
rect 470406 46170 470462 46226
rect 470034 46046 470090 46102
rect 470158 46046 470214 46102
rect 470282 46046 470338 46102
rect 470406 46046 470462 46102
rect 470034 45922 470090 45978
rect 470158 45922 470214 45978
rect 470282 45922 470338 45978
rect 470406 45922 470462 45978
rect 470034 28294 470090 28350
rect 470158 28294 470214 28350
rect 470282 28294 470338 28350
rect 470406 28294 470462 28350
rect 470034 28170 470090 28226
rect 470158 28170 470214 28226
rect 470282 28170 470338 28226
rect 470406 28170 470462 28226
rect 470034 28046 470090 28102
rect 470158 28046 470214 28102
rect 470282 28046 470338 28102
rect 470406 28046 470462 28102
rect 470034 27922 470090 27978
rect 470158 27922 470214 27978
rect 470282 27922 470338 27978
rect 470406 27922 470462 27978
rect 470034 10294 470090 10350
rect 470158 10294 470214 10350
rect 470282 10294 470338 10350
rect 470406 10294 470462 10350
rect 470034 10170 470090 10226
rect 470158 10170 470214 10226
rect 470282 10170 470338 10226
rect 470406 10170 470462 10226
rect 470034 10046 470090 10102
rect 470158 10046 470214 10102
rect 470282 10046 470338 10102
rect 470406 10046 470462 10102
rect 470034 9922 470090 9978
rect 470158 9922 470214 9978
rect 470282 9922 470338 9978
rect 470406 9922 470462 9978
rect 466314 -216 466370 -160
rect 466438 -216 466494 -160
rect 466562 -216 466618 -160
rect 466686 -216 466742 -160
rect 466314 -340 466370 -284
rect 466438 -340 466494 -284
rect 466562 -340 466618 -284
rect 466686 -340 466742 -284
rect 466314 -464 466370 -408
rect 466438 -464 466494 -408
rect 466562 -464 466618 -408
rect 466686 -464 466742 -408
rect 466314 -588 466370 -532
rect 466438 -588 466494 -532
rect 466562 -588 466618 -532
rect 466686 -588 466742 -532
rect 472108 62342 472164 62398
rect 497034 94294 497090 94350
rect 497158 94294 497214 94350
rect 497282 94294 497338 94350
rect 497406 94294 497462 94350
rect 497034 94170 497090 94226
rect 497158 94170 497214 94226
rect 497282 94170 497338 94226
rect 497406 94170 497462 94226
rect 497034 94046 497090 94102
rect 497158 94046 497214 94102
rect 497282 94046 497338 94102
rect 497406 94046 497462 94102
rect 497034 93922 497090 93978
rect 497158 93922 497214 93978
rect 497282 93922 497338 93978
rect 497406 93922 497462 93978
rect 480508 79082 480564 79138
rect 477148 59102 477204 59158
rect 475468 50822 475524 50878
rect 474012 13562 474068 13618
rect 478828 15362 478884 15418
rect 500754 598116 500810 598172
rect 500878 598116 500934 598172
rect 501002 598116 501058 598172
rect 501126 598116 501182 598172
rect 500754 597992 500810 598048
rect 500878 597992 500934 598048
rect 501002 597992 501058 598048
rect 501126 597992 501182 598048
rect 500754 597868 500810 597924
rect 500878 597868 500934 597924
rect 501002 597868 501058 597924
rect 501126 597868 501182 597924
rect 500754 597744 500810 597800
rect 500878 597744 500934 597800
rect 501002 597744 501058 597800
rect 501126 597744 501182 597800
rect 500754 586294 500810 586350
rect 500878 586294 500934 586350
rect 501002 586294 501058 586350
rect 501126 586294 501182 586350
rect 500754 586170 500810 586226
rect 500878 586170 500934 586226
rect 501002 586170 501058 586226
rect 501126 586170 501182 586226
rect 500754 586046 500810 586102
rect 500878 586046 500934 586102
rect 501002 586046 501058 586102
rect 501126 586046 501182 586102
rect 500754 585922 500810 585978
rect 500878 585922 500934 585978
rect 501002 585922 501058 585978
rect 501126 585922 501182 585978
rect 500754 568294 500810 568350
rect 500878 568294 500934 568350
rect 501002 568294 501058 568350
rect 501126 568294 501182 568350
rect 500754 568170 500810 568226
rect 500878 568170 500934 568226
rect 501002 568170 501058 568226
rect 501126 568170 501182 568226
rect 500754 568046 500810 568102
rect 500878 568046 500934 568102
rect 501002 568046 501058 568102
rect 501126 568046 501182 568102
rect 500754 567922 500810 567978
rect 500878 567922 500934 567978
rect 501002 567922 501058 567978
rect 501126 567922 501182 567978
rect 500754 550294 500810 550350
rect 500878 550294 500934 550350
rect 501002 550294 501058 550350
rect 501126 550294 501182 550350
rect 500754 550170 500810 550226
rect 500878 550170 500934 550226
rect 501002 550170 501058 550226
rect 501126 550170 501182 550226
rect 500754 550046 500810 550102
rect 500878 550046 500934 550102
rect 501002 550046 501058 550102
rect 501126 550046 501182 550102
rect 500754 549922 500810 549978
rect 500878 549922 500934 549978
rect 501002 549922 501058 549978
rect 501126 549922 501182 549978
rect 500754 532294 500810 532350
rect 500878 532294 500934 532350
rect 501002 532294 501058 532350
rect 501126 532294 501182 532350
rect 500754 532170 500810 532226
rect 500878 532170 500934 532226
rect 501002 532170 501058 532226
rect 501126 532170 501182 532226
rect 500754 532046 500810 532102
rect 500878 532046 500934 532102
rect 501002 532046 501058 532102
rect 501126 532046 501182 532102
rect 500754 531922 500810 531978
rect 500878 531922 500934 531978
rect 501002 531922 501058 531978
rect 501126 531922 501182 531978
rect 500754 514294 500810 514350
rect 500878 514294 500934 514350
rect 501002 514294 501058 514350
rect 501126 514294 501182 514350
rect 500754 514170 500810 514226
rect 500878 514170 500934 514226
rect 501002 514170 501058 514226
rect 501126 514170 501182 514226
rect 500754 514046 500810 514102
rect 500878 514046 500934 514102
rect 501002 514046 501058 514102
rect 501126 514046 501182 514102
rect 500754 513922 500810 513978
rect 500878 513922 500934 513978
rect 501002 513922 501058 513978
rect 501126 513922 501182 513978
rect 500754 496294 500810 496350
rect 500878 496294 500934 496350
rect 501002 496294 501058 496350
rect 501126 496294 501182 496350
rect 500754 496170 500810 496226
rect 500878 496170 500934 496226
rect 501002 496170 501058 496226
rect 501126 496170 501182 496226
rect 500754 496046 500810 496102
rect 500878 496046 500934 496102
rect 501002 496046 501058 496102
rect 501126 496046 501182 496102
rect 500754 495922 500810 495978
rect 500878 495922 500934 495978
rect 501002 495922 501058 495978
rect 501126 495922 501182 495978
rect 500754 478294 500810 478350
rect 500878 478294 500934 478350
rect 501002 478294 501058 478350
rect 501126 478294 501182 478350
rect 500754 478170 500810 478226
rect 500878 478170 500934 478226
rect 501002 478170 501058 478226
rect 501126 478170 501182 478226
rect 500754 478046 500810 478102
rect 500878 478046 500934 478102
rect 501002 478046 501058 478102
rect 501126 478046 501182 478102
rect 500754 477922 500810 477978
rect 500878 477922 500934 477978
rect 501002 477922 501058 477978
rect 501126 477922 501182 477978
rect 500754 460294 500810 460350
rect 500878 460294 500934 460350
rect 501002 460294 501058 460350
rect 501126 460294 501182 460350
rect 500754 460170 500810 460226
rect 500878 460170 500934 460226
rect 501002 460170 501058 460226
rect 501126 460170 501182 460226
rect 500754 460046 500810 460102
rect 500878 460046 500934 460102
rect 501002 460046 501058 460102
rect 501126 460046 501182 460102
rect 500754 459922 500810 459978
rect 500878 459922 500934 459978
rect 501002 459922 501058 459978
rect 501126 459922 501182 459978
rect 500754 442294 500810 442350
rect 500878 442294 500934 442350
rect 501002 442294 501058 442350
rect 501126 442294 501182 442350
rect 500754 442170 500810 442226
rect 500878 442170 500934 442226
rect 501002 442170 501058 442226
rect 501126 442170 501182 442226
rect 500754 442046 500810 442102
rect 500878 442046 500934 442102
rect 501002 442046 501058 442102
rect 501126 442046 501182 442102
rect 500754 441922 500810 441978
rect 500878 441922 500934 441978
rect 501002 441922 501058 441978
rect 501126 441922 501182 441978
rect 500754 424294 500810 424350
rect 500878 424294 500934 424350
rect 501002 424294 501058 424350
rect 501126 424294 501182 424350
rect 500754 424170 500810 424226
rect 500878 424170 500934 424226
rect 501002 424170 501058 424226
rect 501126 424170 501182 424226
rect 500754 424046 500810 424102
rect 500878 424046 500934 424102
rect 501002 424046 501058 424102
rect 501126 424046 501182 424102
rect 500754 423922 500810 423978
rect 500878 423922 500934 423978
rect 501002 423922 501058 423978
rect 501126 423922 501182 423978
rect 500754 406294 500810 406350
rect 500878 406294 500934 406350
rect 501002 406294 501058 406350
rect 501126 406294 501182 406350
rect 500754 406170 500810 406226
rect 500878 406170 500934 406226
rect 501002 406170 501058 406226
rect 501126 406170 501182 406226
rect 500754 406046 500810 406102
rect 500878 406046 500934 406102
rect 501002 406046 501058 406102
rect 501126 406046 501182 406102
rect 500754 405922 500810 405978
rect 500878 405922 500934 405978
rect 501002 405922 501058 405978
rect 501126 405922 501182 405978
rect 500754 388294 500810 388350
rect 500878 388294 500934 388350
rect 501002 388294 501058 388350
rect 501126 388294 501182 388350
rect 500754 388170 500810 388226
rect 500878 388170 500934 388226
rect 501002 388170 501058 388226
rect 501126 388170 501182 388226
rect 500754 388046 500810 388102
rect 500878 388046 500934 388102
rect 501002 388046 501058 388102
rect 501126 388046 501182 388102
rect 500754 387922 500810 387978
rect 500878 387922 500934 387978
rect 501002 387922 501058 387978
rect 501126 387922 501182 387978
rect 500754 370294 500810 370350
rect 500878 370294 500934 370350
rect 501002 370294 501058 370350
rect 501126 370294 501182 370350
rect 500754 370170 500810 370226
rect 500878 370170 500934 370226
rect 501002 370170 501058 370226
rect 501126 370170 501182 370226
rect 500754 370046 500810 370102
rect 500878 370046 500934 370102
rect 501002 370046 501058 370102
rect 501126 370046 501182 370102
rect 500754 369922 500810 369978
rect 500878 369922 500934 369978
rect 501002 369922 501058 369978
rect 501126 369922 501182 369978
rect 500754 352294 500810 352350
rect 500878 352294 500934 352350
rect 501002 352294 501058 352350
rect 501126 352294 501182 352350
rect 500754 352170 500810 352226
rect 500878 352170 500934 352226
rect 501002 352170 501058 352226
rect 501126 352170 501182 352226
rect 500754 352046 500810 352102
rect 500878 352046 500934 352102
rect 501002 352046 501058 352102
rect 501126 352046 501182 352102
rect 500754 351922 500810 351978
rect 500878 351922 500934 351978
rect 501002 351922 501058 351978
rect 501126 351922 501182 351978
rect 500754 334294 500810 334350
rect 500878 334294 500934 334350
rect 501002 334294 501058 334350
rect 501126 334294 501182 334350
rect 500754 334170 500810 334226
rect 500878 334170 500934 334226
rect 501002 334170 501058 334226
rect 501126 334170 501182 334226
rect 500754 334046 500810 334102
rect 500878 334046 500934 334102
rect 501002 334046 501058 334102
rect 501126 334046 501182 334102
rect 500754 333922 500810 333978
rect 500878 333922 500934 333978
rect 501002 333922 501058 333978
rect 501126 333922 501182 333978
rect 500754 316294 500810 316350
rect 500878 316294 500934 316350
rect 501002 316294 501058 316350
rect 501126 316294 501182 316350
rect 500754 316170 500810 316226
rect 500878 316170 500934 316226
rect 501002 316170 501058 316226
rect 501126 316170 501182 316226
rect 500754 316046 500810 316102
rect 500878 316046 500934 316102
rect 501002 316046 501058 316102
rect 501126 316046 501182 316102
rect 500754 315922 500810 315978
rect 500878 315922 500934 315978
rect 501002 315922 501058 315978
rect 501126 315922 501182 315978
rect 500754 298294 500810 298350
rect 500878 298294 500934 298350
rect 501002 298294 501058 298350
rect 501126 298294 501182 298350
rect 500754 298170 500810 298226
rect 500878 298170 500934 298226
rect 501002 298170 501058 298226
rect 501126 298170 501182 298226
rect 500754 298046 500810 298102
rect 500878 298046 500934 298102
rect 501002 298046 501058 298102
rect 501126 298046 501182 298102
rect 500754 297922 500810 297978
rect 500878 297922 500934 297978
rect 501002 297922 501058 297978
rect 501126 297922 501182 297978
rect 500754 280294 500810 280350
rect 500878 280294 500934 280350
rect 501002 280294 501058 280350
rect 501126 280294 501182 280350
rect 500754 280170 500810 280226
rect 500878 280170 500934 280226
rect 501002 280170 501058 280226
rect 501126 280170 501182 280226
rect 500754 280046 500810 280102
rect 500878 280046 500934 280102
rect 501002 280046 501058 280102
rect 501126 280046 501182 280102
rect 500754 279922 500810 279978
rect 500878 279922 500934 279978
rect 501002 279922 501058 279978
rect 501126 279922 501182 279978
rect 500754 262294 500810 262350
rect 500878 262294 500934 262350
rect 501002 262294 501058 262350
rect 501126 262294 501182 262350
rect 500754 262170 500810 262226
rect 500878 262170 500934 262226
rect 501002 262170 501058 262226
rect 501126 262170 501182 262226
rect 500754 262046 500810 262102
rect 500878 262046 500934 262102
rect 501002 262046 501058 262102
rect 501126 262046 501182 262102
rect 500754 261922 500810 261978
rect 500878 261922 500934 261978
rect 501002 261922 501058 261978
rect 501126 261922 501182 261978
rect 500754 244294 500810 244350
rect 500878 244294 500934 244350
rect 501002 244294 501058 244350
rect 501126 244294 501182 244350
rect 500754 244170 500810 244226
rect 500878 244170 500934 244226
rect 501002 244170 501058 244226
rect 501126 244170 501182 244226
rect 500754 244046 500810 244102
rect 500878 244046 500934 244102
rect 501002 244046 501058 244102
rect 501126 244046 501182 244102
rect 500754 243922 500810 243978
rect 500878 243922 500934 243978
rect 501002 243922 501058 243978
rect 501126 243922 501182 243978
rect 500754 226294 500810 226350
rect 500878 226294 500934 226350
rect 501002 226294 501058 226350
rect 501126 226294 501182 226350
rect 500754 226170 500810 226226
rect 500878 226170 500934 226226
rect 501002 226170 501058 226226
rect 501126 226170 501182 226226
rect 500754 226046 500810 226102
rect 500878 226046 500934 226102
rect 501002 226046 501058 226102
rect 501126 226046 501182 226102
rect 500754 225922 500810 225978
rect 500878 225922 500934 225978
rect 501002 225922 501058 225978
rect 501126 225922 501182 225978
rect 500754 208294 500810 208350
rect 500878 208294 500934 208350
rect 501002 208294 501058 208350
rect 501126 208294 501182 208350
rect 500754 208170 500810 208226
rect 500878 208170 500934 208226
rect 501002 208170 501058 208226
rect 501126 208170 501182 208226
rect 500754 208046 500810 208102
rect 500878 208046 500934 208102
rect 501002 208046 501058 208102
rect 501126 208046 501182 208102
rect 500754 207922 500810 207978
rect 500878 207922 500934 207978
rect 501002 207922 501058 207978
rect 501126 207922 501182 207978
rect 500754 190294 500810 190350
rect 500878 190294 500934 190350
rect 501002 190294 501058 190350
rect 501126 190294 501182 190350
rect 500754 190170 500810 190226
rect 500878 190170 500934 190226
rect 501002 190170 501058 190226
rect 501126 190170 501182 190226
rect 500754 190046 500810 190102
rect 500878 190046 500934 190102
rect 501002 190046 501058 190102
rect 501126 190046 501182 190102
rect 500754 189922 500810 189978
rect 500878 189922 500934 189978
rect 501002 189922 501058 189978
rect 501126 189922 501182 189978
rect 500754 172294 500810 172350
rect 500878 172294 500934 172350
rect 501002 172294 501058 172350
rect 501126 172294 501182 172350
rect 500754 172170 500810 172226
rect 500878 172170 500934 172226
rect 501002 172170 501058 172226
rect 501126 172170 501182 172226
rect 500754 172046 500810 172102
rect 500878 172046 500934 172102
rect 501002 172046 501058 172102
rect 501126 172046 501182 172102
rect 500754 171922 500810 171978
rect 500878 171922 500934 171978
rect 501002 171922 501058 171978
rect 501126 171922 501182 171978
rect 500754 154294 500810 154350
rect 500878 154294 500934 154350
rect 501002 154294 501058 154350
rect 501126 154294 501182 154350
rect 500754 154170 500810 154226
rect 500878 154170 500934 154226
rect 501002 154170 501058 154226
rect 501126 154170 501182 154226
rect 500754 154046 500810 154102
rect 500878 154046 500934 154102
rect 501002 154046 501058 154102
rect 501126 154046 501182 154102
rect 500754 153922 500810 153978
rect 500878 153922 500934 153978
rect 501002 153922 501058 153978
rect 501126 153922 501182 153978
rect 500754 136294 500810 136350
rect 500878 136294 500934 136350
rect 501002 136294 501058 136350
rect 501126 136294 501182 136350
rect 500754 136170 500810 136226
rect 500878 136170 500934 136226
rect 501002 136170 501058 136226
rect 501126 136170 501182 136226
rect 500754 136046 500810 136102
rect 500878 136046 500934 136102
rect 501002 136046 501058 136102
rect 501126 136046 501182 136102
rect 500754 135922 500810 135978
rect 500878 135922 500934 135978
rect 501002 135922 501058 135978
rect 501126 135922 501182 135978
rect 500754 118294 500810 118350
rect 500878 118294 500934 118350
rect 501002 118294 501058 118350
rect 501126 118294 501182 118350
rect 500754 118170 500810 118226
rect 500878 118170 500934 118226
rect 501002 118170 501058 118226
rect 501126 118170 501182 118226
rect 500754 118046 500810 118102
rect 500878 118046 500934 118102
rect 501002 118046 501058 118102
rect 501126 118046 501182 118102
rect 500754 117922 500810 117978
rect 500878 117922 500934 117978
rect 501002 117922 501058 117978
rect 501126 117922 501182 117978
rect 500754 100294 500810 100350
rect 500878 100294 500934 100350
rect 501002 100294 501058 100350
rect 501126 100294 501182 100350
rect 500754 100170 500810 100226
rect 500878 100170 500934 100226
rect 501002 100170 501058 100226
rect 501126 100170 501182 100226
rect 500754 100046 500810 100102
rect 500878 100046 500934 100102
rect 501002 100046 501058 100102
rect 501126 100046 501182 100102
rect 500754 99922 500810 99978
rect 500878 99922 500934 99978
rect 501002 99922 501058 99978
rect 501126 99922 501182 99978
rect 527754 597156 527810 597212
rect 527878 597156 527934 597212
rect 528002 597156 528058 597212
rect 528126 597156 528182 597212
rect 527754 597032 527810 597088
rect 527878 597032 527934 597088
rect 528002 597032 528058 597088
rect 528126 597032 528182 597088
rect 527754 596908 527810 596964
rect 527878 596908 527934 596964
rect 528002 596908 528058 596964
rect 528126 596908 528182 596964
rect 527754 596784 527810 596840
rect 527878 596784 527934 596840
rect 528002 596784 528058 596840
rect 528126 596784 528182 596840
rect 527754 580294 527810 580350
rect 527878 580294 527934 580350
rect 528002 580294 528058 580350
rect 528126 580294 528182 580350
rect 527754 580170 527810 580226
rect 527878 580170 527934 580226
rect 528002 580170 528058 580226
rect 528126 580170 528182 580226
rect 527754 580046 527810 580102
rect 527878 580046 527934 580102
rect 528002 580046 528058 580102
rect 528126 580046 528182 580102
rect 527754 579922 527810 579978
rect 527878 579922 527934 579978
rect 528002 579922 528058 579978
rect 528126 579922 528182 579978
rect 527754 562294 527810 562350
rect 527878 562294 527934 562350
rect 528002 562294 528058 562350
rect 528126 562294 528182 562350
rect 527754 562170 527810 562226
rect 527878 562170 527934 562226
rect 528002 562170 528058 562226
rect 528126 562170 528182 562226
rect 527754 562046 527810 562102
rect 527878 562046 527934 562102
rect 528002 562046 528058 562102
rect 528126 562046 528182 562102
rect 527754 561922 527810 561978
rect 527878 561922 527934 561978
rect 528002 561922 528058 561978
rect 528126 561922 528182 561978
rect 527754 544294 527810 544350
rect 527878 544294 527934 544350
rect 528002 544294 528058 544350
rect 528126 544294 528182 544350
rect 527754 544170 527810 544226
rect 527878 544170 527934 544226
rect 528002 544170 528058 544226
rect 528126 544170 528182 544226
rect 527754 544046 527810 544102
rect 527878 544046 527934 544102
rect 528002 544046 528058 544102
rect 528126 544046 528182 544102
rect 527754 543922 527810 543978
rect 527878 543922 527934 543978
rect 528002 543922 528058 543978
rect 528126 543922 528182 543978
rect 527754 526294 527810 526350
rect 527878 526294 527934 526350
rect 528002 526294 528058 526350
rect 528126 526294 528182 526350
rect 527754 526170 527810 526226
rect 527878 526170 527934 526226
rect 528002 526170 528058 526226
rect 528126 526170 528182 526226
rect 527754 526046 527810 526102
rect 527878 526046 527934 526102
rect 528002 526046 528058 526102
rect 528126 526046 528182 526102
rect 527754 525922 527810 525978
rect 527878 525922 527934 525978
rect 528002 525922 528058 525978
rect 528126 525922 528182 525978
rect 527754 508294 527810 508350
rect 527878 508294 527934 508350
rect 528002 508294 528058 508350
rect 528126 508294 528182 508350
rect 527754 508170 527810 508226
rect 527878 508170 527934 508226
rect 528002 508170 528058 508226
rect 528126 508170 528182 508226
rect 527754 508046 527810 508102
rect 527878 508046 527934 508102
rect 528002 508046 528058 508102
rect 528126 508046 528182 508102
rect 527754 507922 527810 507978
rect 527878 507922 527934 507978
rect 528002 507922 528058 507978
rect 528126 507922 528182 507978
rect 527754 490294 527810 490350
rect 527878 490294 527934 490350
rect 528002 490294 528058 490350
rect 528126 490294 528182 490350
rect 527754 490170 527810 490226
rect 527878 490170 527934 490226
rect 528002 490170 528058 490226
rect 528126 490170 528182 490226
rect 527754 490046 527810 490102
rect 527878 490046 527934 490102
rect 528002 490046 528058 490102
rect 528126 490046 528182 490102
rect 527754 489922 527810 489978
rect 527878 489922 527934 489978
rect 528002 489922 528058 489978
rect 528126 489922 528182 489978
rect 527754 472294 527810 472350
rect 527878 472294 527934 472350
rect 528002 472294 528058 472350
rect 528126 472294 528182 472350
rect 527754 472170 527810 472226
rect 527878 472170 527934 472226
rect 528002 472170 528058 472226
rect 528126 472170 528182 472226
rect 527754 472046 527810 472102
rect 527878 472046 527934 472102
rect 528002 472046 528058 472102
rect 528126 472046 528182 472102
rect 527754 471922 527810 471978
rect 527878 471922 527934 471978
rect 528002 471922 528058 471978
rect 528126 471922 528182 471978
rect 527754 454294 527810 454350
rect 527878 454294 527934 454350
rect 528002 454294 528058 454350
rect 528126 454294 528182 454350
rect 527754 454170 527810 454226
rect 527878 454170 527934 454226
rect 528002 454170 528058 454226
rect 528126 454170 528182 454226
rect 527754 454046 527810 454102
rect 527878 454046 527934 454102
rect 528002 454046 528058 454102
rect 528126 454046 528182 454102
rect 527754 453922 527810 453978
rect 527878 453922 527934 453978
rect 528002 453922 528058 453978
rect 528126 453922 528182 453978
rect 527754 436294 527810 436350
rect 527878 436294 527934 436350
rect 528002 436294 528058 436350
rect 528126 436294 528182 436350
rect 527754 436170 527810 436226
rect 527878 436170 527934 436226
rect 528002 436170 528058 436226
rect 528126 436170 528182 436226
rect 527754 436046 527810 436102
rect 527878 436046 527934 436102
rect 528002 436046 528058 436102
rect 528126 436046 528182 436102
rect 527754 435922 527810 435978
rect 527878 435922 527934 435978
rect 528002 435922 528058 435978
rect 528126 435922 528182 435978
rect 527754 418294 527810 418350
rect 527878 418294 527934 418350
rect 528002 418294 528058 418350
rect 528126 418294 528182 418350
rect 527754 418170 527810 418226
rect 527878 418170 527934 418226
rect 528002 418170 528058 418226
rect 528126 418170 528182 418226
rect 527754 418046 527810 418102
rect 527878 418046 527934 418102
rect 528002 418046 528058 418102
rect 528126 418046 528182 418102
rect 527754 417922 527810 417978
rect 527878 417922 527934 417978
rect 528002 417922 528058 417978
rect 528126 417922 528182 417978
rect 527754 400294 527810 400350
rect 527878 400294 527934 400350
rect 528002 400294 528058 400350
rect 528126 400294 528182 400350
rect 527754 400170 527810 400226
rect 527878 400170 527934 400226
rect 528002 400170 528058 400226
rect 528126 400170 528182 400226
rect 527754 400046 527810 400102
rect 527878 400046 527934 400102
rect 528002 400046 528058 400102
rect 528126 400046 528182 400102
rect 527754 399922 527810 399978
rect 527878 399922 527934 399978
rect 528002 399922 528058 399978
rect 528126 399922 528182 399978
rect 527754 382294 527810 382350
rect 527878 382294 527934 382350
rect 528002 382294 528058 382350
rect 528126 382294 528182 382350
rect 527754 382170 527810 382226
rect 527878 382170 527934 382226
rect 528002 382170 528058 382226
rect 528126 382170 528182 382226
rect 527754 382046 527810 382102
rect 527878 382046 527934 382102
rect 528002 382046 528058 382102
rect 528126 382046 528182 382102
rect 527754 381922 527810 381978
rect 527878 381922 527934 381978
rect 528002 381922 528058 381978
rect 528126 381922 528182 381978
rect 527754 364294 527810 364350
rect 527878 364294 527934 364350
rect 528002 364294 528058 364350
rect 528126 364294 528182 364350
rect 527754 364170 527810 364226
rect 527878 364170 527934 364226
rect 528002 364170 528058 364226
rect 528126 364170 528182 364226
rect 527754 364046 527810 364102
rect 527878 364046 527934 364102
rect 528002 364046 528058 364102
rect 528126 364046 528182 364102
rect 527754 363922 527810 363978
rect 527878 363922 527934 363978
rect 528002 363922 528058 363978
rect 528126 363922 528182 363978
rect 527754 346294 527810 346350
rect 527878 346294 527934 346350
rect 528002 346294 528058 346350
rect 528126 346294 528182 346350
rect 527754 346170 527810 346226
rect 527878 346170 527934 346226
rect 528002 346170 528058 346226
rect 528126 346170 528182 346226
rect 527754 346046 527810 346102
rect 527878 346046 527934 346102
rect 528002 346046 528058 346102
rect 528126 346046 528182 346102
rect 527754 345922 527810 345978
rect 527878 345922 527934 345978
rect 528002 345922 528058 345978
rect 528126 345922 528182 345978
rect 527754 328294 527810 328350
rect 527878 328294 527934 328350
rect 528002 328294 528058 328350
rect 528126 328294 528182 328350
rect 527754 328170 527810 328226
rect 527878 328170 527934 328226
rect 528002 328170 528058 328226
rect 528126 328170 528182 328226
rect 527754 328046 527810 328102
rect 527878 328046 527934 328102
rect 528002 328046 528058 328102
rect 528126 328046 528182 328102
rect 527754 327922 527810 327978
rect 527878 327922 527934 327978
rect 528002 327922 528058 327978
rect 528126 327922 528182 327978
rect 527754 310294 527810 310350
rect 527878 310294 527934 310350
rect 528002 310294 528058 310350
rect 528126 310294 528182 310350
rect 527754 310170 527810 310226
rect 527878 310170 527934 310226
rect 528002 310170 528058 310226
rect 528126 310170 528182 310226
rect 527754 310046 527810 310102
rect 527878 310046 527934 310102
rect 528002 310046 528058 310102
rect 528126 310046 528182 310102
rect 527754 309922 527810 309978
rect 527878 309922 527934 309978
rect 528002 309922 528058 309978
rect 528126 309922 528182 309978
rect 527754 292294 527810 292350
rect 527878 292294 527934 292350
rect 528002 292294 528058 292350
rect 528126 292294 528182 292350
rect 527754 292170 527810 292226
rect 527878 292170 527934 292226
rect 528002 292170 528058 292226
rect 528126 292170 528182 292226
rect 527754 292046 527810 292102
rect 527878 292046 527934 292102
rect 528002 292046 528058 292102
rect 528126 292046 528182 292102
rect 527754 291922 527810 291978
rect 527878 291922 527934 291978
rect 528002 291922 528058 291978
rect 528126 291922 528182 291978
rect 527754 274294 527810 274350
rect 527878 274294 527934 274350
rect 528002 274294 528058 274350
rect 528126 274294 528182 274350
rect 527754 274170 527810 274226
rect 527878 274170 527934 274226
rect 528002 274170 528058 274226
rect 528126 274170 528182 274226
rect 527754 274046 527810 274102
rect 527878 274046 527934 274102
rect 528002 274046 528058 274102
rect 528126 274046 528182 274102
rect 527754 273922 527810 273978
rect 527878 273922 527934 273978
rect 528002 273922 528058 273978
rect 528126 273922 528182 273978
rect 527754 256294 527810 256350
rect 527878 256294 527934 256350
rect 528002 256294 528058 256350
rect 528126 256294 528182 256350
rect 527754 256170 527810 256226
rect 527878 256170 527934 256226
rect 528002 256170 528058 256226
rect 528126 256170 528182 256226
rect 527754 256046 527810 256102
rect 527878 256046 527934 256102
rect 528002 256046 528058 256102
rect 528126 256046 528182 256102
rect 527754 255922 527810 255978
rect 527878 255922 527934 255978
rect 528002 255922 528058 255978
rect 528126 255922 528182 255978
rect 527754 238294 527810 238350
rect 527878 238294 527934 238350
rect 528002 238294 528058 238350
rect 528126 238294 528182 238350
rect 527754 238170 527810 238226
rect 527878 238170 527934 238226
rect 528002 238170 528058 238226
rect 528126 238170 528182 238226
rect 527754 238046 527810 238102
rect 527878 238046 527934 238102
rect 528002 238046 528058 238102
rect 528126 238046 528182 238102
rect 527754 237922 527810 237978
rect 527878 237922 527934 237978
rect 528002 237922 528058 237978
rect 528126 237922 528182 237978
rect 527754 220294 527810 220350
rect 527878 220294 527934 220350
rect 528002 220294 528058 220350
rect 528126 220294 528182 220350
rect 527754 220170 527810 220226
rect 527878 220170 527934 220226
rect 528002 220170 528058 220226
rect 528126 220170 528182 220226
rect 527754 220046 527810 220102
rect 527878 220046 527934 220102
rect 528002 220046 528058 220102
rect 528126 220046 528182 220102
rect 527754 219922 527810 219978
rect 527878 219922 527934 219978
rect 528002 219922 528058 219978
rect 528126 219922 528182 219978
rect 527754 202294 527810 202350
rect 527878 202294 527934 202350
rect 528002 202294 528058 202350
rect 528126 202294 528182 202350
rect 527754 202170 527810 202226
rect 527878 202170 527934 202226
rect 528002 202170 528058 202226
rect 528126 202170 528182 202226
rect 527754 202046 527810 202102
rect 527878 202046 527934 202102
rect 528002 202046 528058 202102
rect 528126 202046 528182 202102
rect 527754 201922 527810 201978
rect 527878 201922 527934 201978
rect 528002 201922 528058 201978
rect 528126 201922 528182 201978
rect 527754 184294 527810 184350
rect 527878 184294 527934 184350
rect 528002 184294 528058 184350
rect 528126 184294 528182 184350
rect 527754 184170 527810 184226
rect 527878 184170 527934 184226
rect 528002 184170 528058 184226
rect 528126 184170 528182 184226
rect 527754 184046 527810 184102
rect 527878 184046 527934 184102
rect 528002 184046 528058 184102
rect 528126 184046 528182 184102
rect 527754 183922 527810 183978
rect 527878 183922 527934 183978
rect 528002 183922 528058 183978
rect 528126 183922 528182 183978
rect 527754 166294 527810 166350
rect 527878 166294 527934 166350
rect 528002 166294 528058 166350
rect 528126 166294 528182 166350
rect 527754 166170 527810 166226
rect 527878 166170 527934 166226
rect 528002 166170 528058 166226
rect 528126 166170 528182 166226
rect 527754 166046 527810 166102
rect 527878 166046 527934 166102
rect 528002 166046 528058 166102
rect 528126 166046 528182 166102
rect 527754 165922 527810 165978
rect 527878 165922 527934 165978
rect 528002 165922 528058 165978
rect 528126 165922 528182 165978
rect 527754 148294 527810 148350
rect 527878 148294 527934 148350
rect 528002 148294 528058 148350
rect 528126 148294 528182 148350
rect 527754 148170 527810 148226
rect 527878 148170 527934 148226
rect 528002 148170 528058 148226
rect 528126 148170 528182 148226
rect 527754 148046 527810 148102
rect 527878 148046 527934 148102
rect 528002 148046 528058 148102
rect 528126 148046 528182 148102
rect 527754 147922 527810 147978
rect 527878 147922 527934 147978
rect 528002 147922 528058 147978
rect 528126 147922 528182 147978
rect 527754 130294 527810 130350
rect 527878 130294 527934 130350
rect 528002 130294 528058 130350
rect 528126 130294 528182 130350
rect 527754 130170 527810 130226
rect 527878 130170 527934 130226
rect 528002 130170 528058 130226
rect 528126 130170 528182 130226
rect 527754 130046 527810 130102
rect 527878 130046 527934 130102
rect 528002 130046 528058 130102
rect 528126 130046 528182 130102
rect 527754 129922 527810 129978
rect 527878 129922 527934 129978
rect 528002 129922 528058 129978
rect 528126 129922 528182 129978
rect 527754 112294 527810 112350
rect 527878 112294 527934 112350
rect 528002 112294 528058 112350
rect 528126 112294 528182 112350
rect 527754 112170 527810 112226
rect 527878 112170 527934 112226
rect 528002 112170 528058 112226
rect 528126 112170 528182 112226
rect 527754 112046 527810 112102
rect 527878 112046 527934 112102
rect 528002 112046 528058 112102
rect 528126 112046 528182 112102
rect 527754 111922 527810 111978
rect 527878 111922 527934 111978
rect 528002 111922 528058 111978
rect 528126 111922 528182 111978
rect 527754 94294 527810 94350
rect 527878 94294 527934 94350
rect 528002 94294 528058 94350
rect 528126 94294 528182 94350
rect 527754 94170 527810 94226
rect 527878 94170 527934 94226
rect 528002 94170 528058 94226
rect 528126 94170 528182 94226
rect 527754 94046 527810 94102
rect 527878 94046 527934 94102
rect 528002 94046 528058 94102
rect 528126 94046 528182 94102
rect 527754 93922 527810 93978
rect 527878 93922 527934 93978
rect 528002 93922 528058 93978
rect 528126 93922 528182 93978
rect 500754 82294 500810 82350
rect 500878 82294 500934 82350
rect 501002 82294 501058 82350
rect 501126 82294 501182 82350
rect 500754 82170 500810 82226
rect 500878 82170 500934 82226
rect 501002 82170 501058 82226
rect 501126 82170 501182 82226
rect 500754 82046 500810 82102
rect 500878 82046 500934 82102
rect 501002 82046 501058 82102
rect 501126 82046 501182 82102
rect 500754 81922 500810 81978
rect 500878 81922 500934 81978
rect 501002 81922 501058 81978
rect 501126 81922 501182 81978
rect 497034 76294 497090 76350
rect 497158 76294 497214 76350
rect 497282 76294 497338 76350
rect 497406 76294 497462 76350
rect 497034 76170 497090 76226
rect 497158 76170 497214 76226
rect 497282 76170 497338 76226
rect 497406 76170 497462 76226
rect 497034 76046 497090 76102
rect 497158 76046 497214 76102
rect 497282 76046 497338 76102
rect 497406 76046 497462 76102
rect 497034 75922 497090 75978
rect 497158 75922 497214 75978
rect 497282 75922 497338 75978
rect 497406 75922 497462 75978
rect 482188 60722 482244 60778
rect 497034 58294 497090 58350
rect 497158 58294 497214 58350
rect 497282 58294 497338 58350
rect 497406 58294 497462 58350
rect 497034 58170 497090 58226
rect 497158 58170 497214 58226
rect 497282 58170 497338 58226
rect 497406 58170 497462 58226
rect 497034 58046 497090 58102
rect 497158 58046 497214 58102
rect 497282 58046 497338 58102
rect 497406 58046 497462 58102
rect 497034 57922 497090 57978
rect 497158 57922 497214 57978
rect 497282 57922 497338 57978
rect 497406 57922 497462 57978
rect 487228 54242 487284 54298
rect 488908 47222 488964 47278
rect 497034 40294 497090 40350
rect 497158 40294 497214 40350
rect 497282 40294 497338 40350
rect 497406 40294 497462 40350
rect 497034 40170 497090 40226
rect 497158 40170 497214 40226
rect 497282 40170 497338 40226
rect 497406 40170 497462 40226
rect 497034 40046 497090 40102
rect 497158 40046 497214 40102
rect 497282 40046 497338 40102
rect 497406 40046 497462 40102
rect 497034 39922 497090 39978
rect 497158 39922 497214 39978
rect 497282 39922 497338 39978
rect 497406 39922 497462 39978
rect 492268 38762 492324 38818
rect 493948 30302 494004 30358
rect 497034 22294 497090 22350
rect 497158 22294 497214 22350
rect 497282 22294 497338 22350
rect 497406 22294 497462 22350
rect 497034 22170 497090 22226
rect 497158 22170 497214 22226
rect 497282 22170 497338 22226
rect 497406 22170 497462 22226
rect 497034 22046 497090 22102
rect 497158 22046 497214 22102
rect 497282 22046 497338 22102
rect 497406 22046 497462 22102
rect 497034 21922 497090 21978
rect 497158 21922 497214 21978
rect 497282 21922 497338 21978
rect 497406 21922 497462 21978
rect 495628 11762 495684 11818
rect 497034 4294 497090 4350
rect 497158 4294 497214 4350
rect 497282 4294 497338 4350
rect 497406 4294 497462 4350
rect 497034 4170 497090 4226
rect 497158 4170 497214 4226
rect 497282 4170 497338 4226
rect 497406 4170 497462 4226
rect 470034 -1176 470090 -1120
rect 470158 -1176 470214 -1120
rect 470282 -1176 470338 -1120
rect 470406 -1176 470462 -1120
rect 470034 -1300 470090 -1244
rect 470158 -1300 470214 -1244
rect 470282 -1300 470338 -1244
rect 470406 -1300 470462 -1244
rect 470034 -1424 470090 -1368
rect 470158 -1424 470214 -1368
rect 470282 -1424 470338 -1368
rect 470406 -1424 470462 -1368
rect 470034 -1548 470090 -1492
rect 470158 -1548 470214 -1492
rect 470282 -1548 470338 -1492
rect 470406 -1548 470462 -1492
rect 497644 77282 497700 77338
rect 500754 64294 500810 64350
rect 500878 64294 500934 64350
rect 501002 64294 501058 64350
rect 501126 64294 501182 64350
rect 500754 64170 500810 64226
rect 500878 64170 500934 64226
rect 501002 64170 501058 64226
rect 501126 64170 501182 64226
rect 500754 64046 500810 64102
rect 500878 64046 500934 64102
rect 501002 64046 501058 64102
rect 501126 64046 501182 64102
rect 500754 63922 500810 63978
rect 500878 63922 500934 63978
rect 501002 63922 501058 63978
rect 501126 63922 501182 63978
rect 500754 46294 500810 46350
rect 500878 46294 500934 46350
rect 501002 46294 501058 46350
rect 501126 46294 501182 46350
rect 500754 46170 500810 46226
rect 500878 46170 500934 46226
rect 501002 46170 501058 46226
rect 501126 46170 501182 46226
rect 500754 46046 500810 46102
rect 500878 46046 500934 46102
rect 501002 46046 501058 46102
rect 501126 46046 501182 46102
rect 500754 45922 500810 45978
rect 500878 45922 500934 45978
rect 501002 45922 501058 45978
rect 501126 45922 501182 45978
rect 527754 76294 527810 76350
rect 527878 76294 527934 76350
rect 528002 76294 528058 76350
rect 528126 76294 528182 76350
rect 527754 76170 527810 76226
rect 527878 76170 527934 76226
rect 528002 76170 528058 76226
rect 528126 76170 528182 76226
rect 527754 76046 527810 76102
rect 527878 76046 527934 76102
rect 528002 76046 528058 76102
rect 528126 76046 528182 76102
rect 527754 75922 527810 75978
rect 527878 75922 527934 75978
rect 528002 75922 528058 75978
rect 528126 75922 528182 75978
rect 525868 62162 525924 62218
rect 515788 60542 515844 60598
rect 509068 57302 509124 57358
rect 505708 35342 505764 35398
rect 500754 28294 500810 28350
rect 500878 28294 500934 28350
rect 501002 28294 501058 28350
rect 501126 28294 501182 28350
rect 500754 28170 500810 28226
rect 500878 28170 500934 28226
rect 501002 28170 501058 28226
rect 501126 28170 501182 28226
rect 500754 28046 500810 28102
rect 500878 28046 500934 28102
rect 501002 28046 501058 28102
rect 501126 28046 501182 28102
rect 500754 27922 500810 27978
rect 500878 27922 500934 27978
rect 501002 27922 501058 27978
rect 501126 27922 501182 27978
rect 500754 10294 500810 10350
rect 500878 10294 500934 10350
rect 501002 10294 501058 10350
rect 501126 10294 501182 10350
rect 500754 10170 500810 10226
rect 500878 10170 500934 10226
rect 501002 10170 501058 10226
rect 501126 10170 501182 10226
rect 500754 10046 500810 10102
rect 500878 10046 500934 10102
rect 501002 10046 501058 10102
rect 501126 10046 501182 10102
rect 500754 9922 500810 9978
rect 500878 9922 500934 9978
rect 501002 9922 501058 9978
rect 501126 9922 501182 9978
rect 497034 4046 497090 4102
rect 497158 4046 497214 4102
rect 497282 4046 497338 4102
rect 497406 4046 497462 4102
rect 497034 3922 497090 3978
rect 497158 3922 497214 3978
rect 497282 3922 497338 3978
rect 497406 3922 497462 3978
rect 497034 -216 497090 -160
rect 497158 -216 497214 -160
rect 497282 -216 497338 -160
rect 497406 -216 497462 -160
rect 497034 -340 497090 -284
rect 497158 -340 497214 -284
rect 497282 -340 497338 -284
rect 497406 -340 497462 -284
rect 497034 -464 497090 -408
rect 497158 -464 497214 -408
rect 497282 -464 497338 -408
rect 497406 -464 497462 -408
rect 497034 -588 497090 -532
rect 497158 -588 497214 -532
rect 497282 -588 497338 -532
rect 497406 -588 497462 -532
rect 501340 28682 501396 28738
rect 504028 16802 504084 16858
rect 508284 10682 508340 10738
rect 510748 54062 510804 54118
rect 520828 58922 520884 58978
rect 517468 52262 517524 52318
rect 522508 55682 522564 55738
rect 527754 58294 527810 58350
rect 527878 58294 527934 58350
rect 528002 58294 528058 58350
rect 528126 58294 528182 58350
rect 527754 58170 527810 58226
rect 527878 58170 527934 58226
rect 528002 58170 528058 58226
rect 528126 58170 528182 58226
rect 527754 58046 527810 58102
rect 527878 58046 527934 58102
rect 528002 58046 528058 58102
rect 528126 58046 528182 58102
rect 527754 57922 527810 57978
rect 527878 57922 527934 57978
rect 528002 57922 528058 57978
rect 528126 57922 528182 57978
rect 527754 40294 527810 40350
rect 527878 40294 527934 40350
rect 528002 40294 528058 40350
rect 528126 40294 528182 40350
rect 527754 40170 527810 40226
rect 527878 40170 527934 40226
rect 528002 40170 528058 40226
rect 528126 40170 528182 40226
rect 527754 40046 527810 40102
rect 527878 40046 527934 40102
rect 528002 40046 528058 40102
rect 528126 40046 528182 40102
rect 527754 39922 527810 39978
rect 527878 39922 527934 39978
rect 528002 39922 528058 39978
rect 528126 39922 528182 39978
rect 527754 22294 527810 22350
rect 527878 22294 527934 22350
rect 528002 22294 528058 22350
rect 528126 22294 528182 22350
rect 527754 22170 527810 22226
rect 527878 22170 527934 22226
rect 528002 22170 528058 22226
rect 528126 22170 528182 22226
rect 527754 22046 527810 22102
rect 527878 22046 527934 22102
rect 528002 22046 528058 22102
rect 528126 22046 528182 22102
rect 527754 21922 527810 21978
rect 527878 21922 527934 21978
rect 528002 21922 528058 21978
rect 528126 21922 528182 21978
rect 531474 598116 531530 598172
rect 531598 598116 531654 598172
rect 531722 598116 531778 598172
rect 531846 598116 531902 598172
rect 531474 597992 531530 598048
rect 531598 597992 531654 598048
rect 531722 597992 531778 598048
rect 531846 597992 531902 598048
rect 531474 597868 531530 597924
rect 531598 597868 531654 597924
rect 531722 597868 531778 597924
rect 531846 597868 531902 597924
rect 531474 597744 531530 597800
rect 531598 597744 531654 597800
rect 531722 597744 531778 597800
rect 531846 597744 531902 597800
rect 531474 586294 531530 586350
rect 531598 586294 531654 586350
rect 531722 586294 531778 586350
rect 531846 586294 531902 586350
rect 531474 586170 531530 586226
rect 531598 586170 531654 586226
rect 531722 586170 531778 586226
rect 531846 586170 531902 586226
rect 531474 586046 531530 586102
rect 531598 586046 531654 586102
rect 531722 586046 531778 586102
rect 531846 586046 531902 586102
rect 531474 585922 531530 585978
rect 531598 585922 531654 585978
rect 531722 585922 531778 585978
rect 531846 585922 531902 585978
rect 531474 568294 531530 568350
rect 531598 568294 531654 568350
rect 531722 568294 531778 568350
rect 531846 568294 531902 568350
rect 531474 568170 531530 568226
rect 531598 568170 531654 568226
rect 531722 568170 531778 568226
rect 531846 568170 531902 568226
rect 531474 568046 531530 568102
rect 531598 568046 531654 568102
rect 531722 568046 531778 568102
rect 531846 568046 531902 568102
rect 531474 567922 531530 567978
rect 531598 567922 531654 567978
rect 531722 567922 531778 567978
rect 531846 567922 531902 567978
rect 531474 550294 531530 550350
rect 531598 550294 531654 550350
rect 531722 550294 531778 550350
rect 531846 550294 531902 550350
rect 531474 550170 531530 550226
rect 531598 550170 531654 550226
rect 531722 550170 531778 550226
rect 531846 550170 531902 550226
rect 531474 550046 531530 550102
rect 531598 550046 531654 550102
rect 531722 550046 531778 550102
rect 531846 550046 531902 550102
rect 531474 549922 531530 549978
rect 531598 549922 531654 549978
rect 531722 549922 531778 549978
rect 531846 549922 531902 549978
rect 531474 532294 531530 532350
rect 531598 532294 531654 532350
rect 531722 532294 531778 532350
rect 531846 532294 531902 532350
rect 531474 532170 531530 532226
rect 531598 532170 531654 532226
rect 531722 532170 531778 532226
rect 531846 532170 531902 532226
rect 531474 532046 531530 532102
rect 531598 532046 531654 532102
rect 531722 532046 531778 532102
rect 531846 532046 531902 532102
rect 531474 531922 531530 531978
rect 531598 531922 531654 531978
rect 531722 531922 531778 531978
rect 531846 531922 531902 531978
rect 531474 514294 531530 514350
rect 531598 514294 531654 514350
rect 531722 514294 531778 514350
rect 531846 514294 531902 514350
rect 531474 514170 531530 514226
rect 531598 514170 531654 514226
rect 531722 514170 531778 514226
rect 531846 514170 531902 514226
rect 531474 514046 531530 514102
rect 531598 514046 531654 514102
rect 531722 514046 531778 514102
rect 531846 514046 531902 514102
rect 531474 513922 531530 513978
rect 531598 513922 531654 513978
rect 531722 513922 531778 513978
rect 531846 513922 531902 513978
rect 531474 496294 531530 496350
rect 531598 496294 531654 496350
rect 531722 496294 531778 496350
rect 531846 496294 531902 496350
rect 531474 496170 531530 496226
rect 531598 496170 531654 496226
rect 531722 496170 531778 496226
rect 531846 496170 531902 496226
rect 531474 496046 531530 496102
rect 531598 496046 531654 496102
rect 531722 496046 531778 496102
rect 531846 496046 531902 496102
rect 531474 495922 531530 495978
rect 531598 495922 531654 495978
rect 531722 495922 531778 495978
rect 531846 495922 531902 495978
rect 531474 478294 531530 478350
rect 531598 478294 531654 478350
rect 531722 478294 531778 478350
rect 531846 478294 531902 478350
rect 531474 478170 531530 478226
rect 531598 478170 531654 478226
rect 531722 478170 531778 478226
rect 531846 478170 531902 478226
rect 531474 478046 531530 478102
rect 531598 478046 531654 478102
rect 531722 478046 531778 478102
rect 531846 478046 531902 478102
rect 531474 477922 531530 477978
rect 531598 477922 531654 477978
rect 531722 477922 531778 477978
rect 531846 477922 531902 477978
rect 531474 460294 531530 460350
rect 531598 460294 531654 460350
rect 531722 460294 531778 460350
rect 531846 460294 531902 460350
rect 531474 460170 531530 460226
rect 531598 460170 531654 460226
rect 531722 460170 531778 460226
rect 531846 460170 531902 460226
rect 531474 460046 531530 460102
rect 531598 460046 531654 460102
rect 531722 460046 531778 460102
rect 531846 460046 531902 460102
rect 531474 459922 531530 459978
rect 531598 459922 531654 459978
rect 531722 459922 531778 459978
rect 531846 459922 531902 459978
rect 531474 442294 531530 442350
rect 531598 442294 531654 442350
rect 531722 442294 531778 442350
rect 531846 442294 531902 442350
rect 531474 442170 531530 442226
rect 531598 442170 531654 442226
rect 531722 442170 531778 442226
rect 531846 442170 531902 442226
rect 531474 442046 531530 442102
rect 531598 442046 531654 442102
rect 531722 442046 531778 442102
rect 531846 442046 531902 442102
rect 531474 441922 531530 441978
rect 531598 441922 531654 441978
rect 531722 441922 531778 441978
rect 531846 441922 531902 441978
rect 531474 424294 531530 424350
rect 531598 424294 531654 424350
rect 531722 424294 531778 424350
rect 531846 424294 531902 424350
rect 531474 424170 531530 424226
rect 531598 424170 531654 424226
rect 531722 424170 531778 424226
rect 531846 424170 531902 424226
rect 531474 424046 531530 424102
rect 531598 424046 531654 424102
rect 531722 424046 531778 424102
rect 531846 424046 531902 424102
rect 531474 423922 531530 423978
rect 531598 423922 531654 423978
rect 531722 423922 531778 423978
rect 531846 423922 531902 423978
rect 531474 406294 531530 406350
rect 531598 406294 531654 406350
rect 531722 406294 531778 406350
rect 531846 406294 531902 406350
rect 531474 406170 531530 406226
rect 531598 406170 531654 406226
rect 531722 406170 531778 406226
rect 531846 406170 531902 406226
rect 531474 406046 531530 406102
rect 531598 406046 531654 406102
rect 531722 406046 531778 406102
rect 531846 406046 531902 406102
rect 531474 405922 531530 405978
rect 531598 405922 531654 405978
rect 531722 405922 531778 405978
rect 531846 405922 531902 405978
rect 531474 388294 531530 388350
rect 531598 388294 531654 388350
rect 531722 388294 531778 388350
rect 531846 388294 531902 388350
rect 531474 388170 531530 388226
rect 531598 388170 531654 388226
rect 531722 388170 531778 388226
rect 531846 388170 531902 388226
rect 531474 388046 531530 388102
rect 531598 388046 531654 388102
rect 531722 388046 531778 388102
rect 531846 388046 531902 388102
rect 531474 387922 531530 387978
rect 531598 387922 531654 387978
rect 531722 387922 531778 387978
rect 531846 387922 531902 387978
rect 531474 370294 531530 370350
rect 531598 370294 531654 370350
rect 531722 370294 531778 370350
rect 531846 370294 531902 370350
rect 531474 370170 531530 370226
rect 531598 370170 531654 370226
rect 531722 370170 531778 370226
rect 531846 370170 531902 370226
rect 531474 370046 531530 370102
rect 531598 370046 531654 370102
rect 531722 370046 531778 370102
rect 531846 370046 531902 370102
rect 531474 369922 531530 369978
rect 531598 369922 531654 369978
rect 531722 369922 531778 369978
rect 531846 369922 531902 369978
rect 531474 352294 531530 352350
rect 531598 352294 531654 352350
rect 531722 352294 531778 352350
rect 531846 352294 531902 352350
rect 531474 352170 531530 352226
rect 531598 352170 531654 352226
rect 531722 352170 531778 352226
rect 531846 352170 531902 352226
rect 531474 352046 531530 352102
rect 531598 352046 531654 352102
rect 531722 352046 531778 352102
rect 531846 352046 531902 352102
rect 531474 351922 531530 351978
rect 531598 351922 531654 351978
rect 531722 351922 531778 351978
rect 531846 351922 531902 351978
rect 531474 334294 531530 334350
rect 531598 334294 531654 334350
rect 531722 334294 531778 334350
rect 531846 334294 531902 334350
rect 531474 334170 531530 334226
rect 531598 334170 531654 334226
rect 531722 334170 531778 334226
rect 531846 334170 531902 334226
rect 531474 334046 531530 334102
rect 531598 334046 531654 334102
rect 531722 334046 531778 334102
rect 531846 334046 531902 334102
rect 531474 333922 531530 333978
rect 531598 333922 531654 333978
rect 531722 333922 531778 333978
rect 531846 333922 531902 333978
rect 531474 316294 531530 316350
rect 531598 316294 531654 316350
rect 531722 316294 531778 316350
rect 531846 316294 531902 316350
rect 531474 316170 531530 316226
rect 531598 316170 531654 316226
rect 531722 316170 531778 316226
rect 531846 316170 531902 316226
rect 531474 316046 531530 316102
rect 531598 316046 531654 316102
rect 531722 316046 531778 316102
rect 531846 316046 531902 316102
rect 531474 315922 531530 315978
rect 531598 315922 531654 315978
rect 531722 315922 531778 315978
rect 531846 315922 531902 315978
rect 531474 298294 531530 298350
rect 531598 298294 531654 298350
rect 531722 298294 531778 298350
rect 531846 298294 531902 298350
rect 531474 298170 531530 298226
rect 531598 298170 531654 298226
rect 531722 298170 531778 298226
rect 531846 298170 531902 298226
rect 531474 298046 531530 298102
rect 531598 298046 531654 298102
rect 531722 298046 531778 298102
rect 531846 298046 531902 298102
rect 531474 297922 531530 297978
rect 531598 297922 531654 297978
rect 531722 297922 531778 297978
rect 531846 297922 531902 297978
rect 531474 280294 531530 280350
rect 531598 280294 531654 280350
rect 531722 280294 531778 280350
rect 531846 280294 531902 280350
rect 531474 280170 531530 280226
rect 531598 280170 531654 280226
rect 531722 280170 531778 280226
rect 531846 280170 531902 280226
rect 531474 280046 531530 280102
rect 531598 280046 531654 280102
rect 531722 280046 531778 280102
rect 531846 280046 531902 280102
rect 531474 279922 531530 279978
rect 531598 279922 531654 279978
rect 531722 279922 531778 279978
rect 531846 279922 531902 279978
rect 531474 262294 531530 262350
rect 531598 262294 531654 262350
rect 531722 262294 531778 262350
rect 531846 262294 531902 262350
rect 531474 262170 531530 262226
rect 531598 262170 531654 262226
rect 531722 262170 531778 262226
rect 531846 262170 531902 262226
rect 531474 262046 531530 262102
rect 531598 262046 531654 262102
rect 531722 262046 531778 262102
rect 531846 262046 531902 262102
rect 531474 261922 531530 261978
rect 531598 261922 531654 261978
rect 531722 261922 531778 261978
rect 531846 261922 531902 261978
rect 531474 244294 531530 244350
rect 531598 244294 531654 244350
rect 531722 244294 531778 244350
rect 531846 244294 531902 244350
rect 531474 244170 531530 244226
rect 531598 244170 531654 244226
rect 531722 244170 531778 244226
rect 531846 244170 531902 244226
rect 531474 244046 531530 244102
rect 531598 244046 531654 244102
rect 531722 244046 531778 244102
rect 531846 244046 531902 244102
rect 531474 243922 531530 243978
rect 531598 243922 531654 243978
rect 531722 243922 531778 243978
rect 531846 243922 531902 243978
rect 531474 226294 531530 226350
rect 531598 226294 531654 226350
rect 531722 226294 531778 226350
rect 531846 226294 531902 226350
rect 531474 226170 531530 226226
rect 531598 226170 531654 226226
rect 531722 226170 531778 226226
rect 531846 226170 531902 226226
rect 531474 226046 531530 226102
rect 531598 226046 531654 226102
rect 531722 226046 531778 226102
rect 531846 226046 531902 226102
rect 531474 225922 531530 225978
rect 531598 225922 531654 225978
rect 531722 225922 531778 225978
rect 531846 225922 531902 225978
rect 531474 208294 531530 208350
rect 531598 208294 531654 208350
rect 531722 208294 531778 208350
rect 531846 208294 531902 208350
rect 531474 208170 531530 208226
rect 531598 208170 531654 208226
rect 531722 208170 531778 208226
rect 531846 208170 531902 208226
rect 531474 208046 531530 208102
rect 531598 208046 531654 208102
rect 531722 208046 531778 208102
rect 531846 208046 531902 208102
rect 531474 207922 531530 207978
rect 531598 207922 531654 207978
rect 531722 207922 531778 207978
rect 531846 207922 531902 207978
rect 531474 190294 531530 190350
rect 531598 190294 531654 190350
rect 531722 190294 531778 190350
rect 531846 190294 531902 190350
rect 531474 190170 531530 190226
rect 531598 190170 531654 190226
rect 531722 190170 531778 190226
rect 531846 190170 531902 190226
rect 531474 190046 531530 190102
rect 531598 190046 531654 190102
rect 531722 190046 531778 190102
rect 531846 190046 531902 190102
rect 531474 189922 531530 189978
rect 531598 189922 531654 189978
rect 531722 189922 531778 189978
rect 531846 189922 531902 189978
rect 531474 172294 531530 172350
rect 531598 172294 531654 172350
rect 531722 172294 531778 172350
rect 531846 172294 531902 172350
rect 531474 172170 531530 172226
rect 531598 172170 531654 172226
rect 531722 172170 531778 172226
rect 531846 172170 531902 172226
rect 531474 172046 531530 172102
rect 531598 172046 531654 172102
rect 531722 172046 531778 172102
rect 531846 172046 531902 172102
rect 531474 171922 531530 171978
rect 531598 171922 531654 171978
rect 531722 171922 531778 171978
rect 531846 171922 531902 171978
rect 531474 154294 531530 154350
rect 531598 154294 531654 154350
rect 531722 154294 531778 154350
rect 531846 154294 531902 154350
rect 531474 154170 531530 154226
rect 531598 154170 531654 154226
rect 531722 154170 531778 154226
rect 531846 154170 531902 154226
rect 531474 154046 531530 154102
rect 531598 154046 531654 154102
rect 531722 154046 531778 154102
rect 531846 154046 531902 154102
rect 531474 153922 531530 153978
rect 531598 153922 531654 153978
rect 531722 153922 531778 153978
rect 531846 153922 531902 153978
rect 531474 136294 531530 136350
rect 531598 136294 531654 136350
rect 531722 136294 531778 136350
rect 531846 136294 531902 136350
rect 531474 136170 531530 136226
rect 531598 136170 531654 136226
rect 531722 136170 531778 136226
rect 531846 136170 531902 136226
rect 531474 136046 531530 136102
rect 531598 136046 531654 136102
rect 531722 136046 531778 136102
rect 531846 136046 531902 136102
rect 531474 135922 531530 135978
rect 531598 135922 531654 135978
rect 531722 135922 531778 135978
rect 531846 135922 531902 135978
rect 531474 118294 531530 118350
rect 531598 118294 531654 118350
rect 531722 118294 531778 118350
rect 531846 118294 531902 118350
rect 531474 118170 531530 118226
rect 531598 118170 531654 118226
rect 531722 118170 531778 118226
rect 531846 118170 531902 118226
rect 531474 118046 531530 118102
rect 531598 118046 531654 118102
rect 531722 118046 531778 118102
rect 531846 118046 531902 118102
rect 531474 117922 531530 117978
rect 531598 117922 531654 117978
rect 531722 117922 531778 117978
rect 531846 117922 531902 117978
rect 531474 100294 531530 100350
rect 531598 100294 531654 100350
rect 531722 100294 531778 100350
rect 531846 100294 531902 100350
rect 531474 100170 531530 100226
rect 531598 100170 531654 100226
rect 531722 100170 531778 100226
rect 531846 100170 531902 100226
rect 531474 100046 531530 100102
rect 531598 100046 531654 100102
rect 531722 100046 531778 100102
rect 531846 100046 531902 100102
rect 531474 99922 531530 99978
rect 531598 99922 531654 99978
rect 531722 99922 531778 99978
rect 531846 99922 531902 99978
rect 531474 82294 531530 82350
rect 531598 82294 531654 82350
rect 531722 82294 531778 82350
rect 531846 82294 531902 82350
rect 531474 82170 531530 82226
rect 531598 82170 531654 82226
rect 531722 82170 531778 82226
rect 531846 82170 531902 82226
rect 531474 82046 531530 82102
rect 531598 82046 531654 82102
rect 531722 82046 531778 82102
rect 531846 82046 531902 82102
rect 531474 81922 531530 81978
rect 531598 81922 531654 81978
rect 531722 81922 531778 81978
rect 531846 81922 531902 81978
rect 531474 64294 531530 64350
rect 531598 64294 531654 64350
rect 531722 64294 531778 64350
rect 531846 64294 531902 64350
rect 531474 64170 531530 64226
rect 531598 64170 531654 64226
rect 531722 64170 531778 64226
rect 531846 64170 531902 64226
rect 531474 64046 531530 64102
rect 531598 64046 531654 64102
rect 531722 64046 531778 64102
rect 531846 64046 531902 64102
rect 531474 63922 531530 63978
rect 531598 63922 531654 63978
rect 531722 63922 531778 63978
rect 531846 63922 531902 63978
rect 558474 597156 558530 597212
rect 558598 597156 558654 597212
rect 558722 597156 558778 597212
rect 558846 597156 558902 597212
rect 558474 597032 558530 597088
rect 558598 597032 558654 597088
rect 558722 597032 558778 597088
rect 558846 597032 558902 597088
rect 558474 596908 558530 596964
rect 558598 596908 558654 596964
rect 558722 596908 558778 596964
rect 558846 596908 558902 596964
rect 558474 596784 558530 596840
rect 558598 596784 558654 596840
rect 558722 596784 558778 596840
rect 558846 596784 558902 596840
rect 558474 580294 558530 580350
rect 558598 580294 558654 580350
rect 558722 580294 558778 580350
rect 558846 580294 558902 580350
rect 558474 580170 558530 580226
rect 558598 580170 558654 580226
rect 558722 580170 558778 580226
rect 558846 580170 558902 580226
rect 558474 580046 558530 580102
rect 558598 580046 558654 580102
rect 558722 580046 558778 580102
rect 558846 580046 558902 580102
rect 558474 579922 558530 579978
rect 558598 579922 558654 579978
rect 558722 579922 558778 579978
rect 558846 579922 558902 579978
rect 558474 562294 558530 562350
rect 558598 562294 558654 562350
rect 558722 562294 558778 562350
rect 558846 562294 558902 562350
rect 558474 562170 558530 562226
rect 558598 562170 558654 562226
rect 558722 562170 558778 562226
rect 558846 562170 558902 562226
rect 558474 562046 558530 562102
rect 558598 562046 558654 562102
rect 558722 562046 558778 562102
rect 558846 562046 558902 562102
rect 558474 561922 558530 561978
rect 558598 561922 558654 561978
rect 558722 561922 558778 561978
rect 558846 561922 558902 561978
rect 558474 544294 558530 544350
rect 558598 544294 558654 544350
rect 558722 544294 558778 544350
rect 558846 544294 558902 544350
rect 558474 544170 558530 544226
rect 558598 544170 558654 544226
rect 558722 544170 558778 544226
rect 558846 544170 558902 544226
rect 558474 544046 558530 544102
rect 558598 544046 558654 544102
rect 558722 544046 558778 544102
rect 558846 544046 558902 544102
rect 558474 543922 558530 543978
rect 558598 543922 558654 543978
rect 558722 543922 558778 543978
rect 558846 543922 558902 543978
rect 558474 526294 558530 526350
rect 558598 526294 558654 526350
rect 558722 526294 558778 526350
rect 558846 526294 558902 526350
rect 558474 526170 558530 526226
rect 558598 526170 558654 526226
rect 558722 526170 558778 526226
rect 558846 526170 558902 526226
rect 558474 526046 558530 526102
rect 558598 526046 558654 526102
rect 558722 526046 558778 526102
rect 558846 526046 558902 526102
rect 558474 525922 558530 525978
rect 558598 525922 558654 525978
rect 558722 525922 558778 525978
rect 558846 525922 558902 525978
rect 558474 508294 558530 508350
rect 558598 508294 558654 508350
rect 558722 508294 558778 508350
rect 558846 508294 558902 508350
rect 558474 508170 558530 508226
rect 558598 508170 558654 508226
rect 558722 508170 558778 508226
rect 558846 508170 558902 508226
rect 558474 508046 558530 508102
rect 558598 508046 558654 508102
rect 558722 508046 558778 508102
rect 558846 508046 558902 508102
rect 558474 507922 558530 507978
rect 558598 507922 558654 507978
rect 558722 507922 558778 507978
rect 558846 507922 558902 507978
rect 558474 490294 558530 490350
rect 558598 490294 558654 490350
rect 558722 490294 558778 490350
rect 558846 490294 558902 490350
rect 558474 490170 558530 490226
rect 558598 490170 558654 490226
rect 558722 490170 558778 490226
rect 558846 490170 558902 490226
rect 558474 490046 558530 490102
rect 558598 490046 558654 490102
rect 558722 490046 558778 490102
rect 558846 490046 558902 490102
rect 558474 489922 558530 489978
rect 558598 489922 558654 489978
rect 558722 489922 558778 489978
rect 558846 489922 558902 489978
rect 558474 472294 558530 472350
rect 558598 472294 558654 472350
rect 558722 472294 558778 472350
rect 558846 472294 558902 472350
rect 558474 472170 558530 472226
rect 558598 472170 558654 472226
rect 558722 472170 558778 472226
rect 558846 472170 558902 472226
rect 558474 472046 558530 472102
rect 558598 472046 558654 472102
rect 558722 472046 558778 472102
rect 558846 472046 558902 472102
rect 558474 471922 558530 471978
rect 558598 471922 558654 471978
rect 558722 471922 558778 471978
rect 558846 471922 558902 471978
rect 558474 454294 558530 454350
rect 558598 454294 558654 454350
rect 558722 454294 558778 454350
rect 558846 454294 558902 454350
rect 558474 454170 558530 454226
rect 558598 454170 558654 454226
rect 558722 454170 558778 454226
rect 558846 454170 558902 454226
rect 558474 454046 558530 454102
rect 558598 454046 558654 454102
rect 558722 454046 558778 454102
rect 558846 454046 558902 454102
rect 558474 453922 558530 453978
rect 558598 453922 558654 453978
rect 558722 453922 558778 453978
rect 558846 453922 558902 453978
rect 558474 436294 558530 436350
rect 558598 436294 558654 436350
rect 558722 436294 558778 436350
rect 558846 436294 558902 436350
rect 558474 436170 558530 436226
rect 558598 436170 558654 436226
rect 558722 436170 558778 436226
rect 558846 436170 558902 436226
rect 558474 436046 558530 436102
rect 558598 436046 558654 436102
rect 558722 436046 558778 436102
rect 558846 436046 558902 436102
rect 558474 435922 558530 435978
rect 558598 435922 558654 435978
rect 558722 435922 558778 435978
rect 558846 435922 558902 435978
rect 558474 418294 558530 418350
rect 558598 418294 558654 418350
rect 558722 418294 558778 418350
rect 558846 418294 558902 418350
rect 558474 418170 558530 418226
rect 558598 418170 558654 418226
rect 558722 418170 558778 418226
rect 558846 418170 558902 418226
rect 558474 418046 558530 418102
rect 558598 418046 558654 418102
rect 558722 418046 558778 418102
rect 558846 418046 558902 418102
rect 558474 417922 558530 417978
rect 558598 417922 558654 417978
rect 558722 417922 558778 417978
rect 558846 417922 558902 417978
rect 558474 400294 558530 400350
rect 558598 400294 558654 400350
rect 558722 400294 558778 400350
rect 558846 400294 558902 400350
rect 558474 400170 558530 400226
rect 558598 400170 558654 400226
rect 558722 400170 558778 400226
rect 558846 400170 558902 400226
rect 558474 400046 558530 400102
rect 558598 400046 558654 400102
rect 558722 400046 558778 400102
rect 558846 400046 558902 400102
rect 558474 399922 558530 399978
rect 558598 399922 558654 399978
rect 558722 399922 558778 399978
rect 558846 399922 558902 399978
rect 558474 382294 558530 382350
rect 558598 382294 558654 382350
rect 558722 382294 558778 382350
rect 558846 382294 558902 382350
rect 558474 382170 558530 382226
rect 558598 382170 558654 382226
rect 558722 382170 558778 382226
rect 558846 382170 558902 382226
rect 558474 382046 558530 382102
rect 558598 382046 558654 382102
rect 558722 382046 558778 382102
rect 558846 382046 558902 382102
rect 558474 381922 558530 381978
rect 558598 381922 558654 381978
rect 558722 381922 558778 381978
rect 558846 381922 558902 381978
rect 558474 364294 558530 364350
rect 558598 364294 558654 364350
rect 558722 364294 558778 364350
rect 558846 364294 558902 364350
rect 558474 364170 558530 364226
rect 558598 364170 558654 364226
rect 558722 364170 558778 364226
rect 558846 364170 558902 364226
rect 558474 364046 558530 364102
rect 558598 364046 558654 364102
rect 558722 364046 558778 364102
rect 558846 364046 558902 364102
rect 558474 363922 558530 363978
rect 558598 363922 558654 363978
rect 558722 363922 558778 363978
rect 558846 363922 558902 363978
rect 558474 346294 558530 346350
rect 558598 346294 558654 346350
rect 558722 346294 558778 346350
rect 558846 346294 558902 346350
rect 558474 346170 558530 346226
rect 558598 346170 558654 346226
rect 558722 346170 558778 346226
rect 558846 346170 558902 346226
rect 558474 346046 558530 346102
rect 558598 346046 558654 346102
rect 558722 346046 558778 346102
rect 558846 346046 558902 346102
rect 558474 345922 558530 345978
rect 558598 345922 558654 345978
rect 558722 345922 558778 345978
rect 558846 345922 558902 345978
rect 558474 328294 558530 328350
rect 558598 328294 558654 328350
rect 558722 328294 558778 328350
rect 558846 328294 558902 328350
rect 558474 328170 558530 328226
rect 558598 328170 558654 328226
rect 558722 328170 558778 328226
rect 558846 328170 558902 328226
rect 558474 328046 558530 328102
rect 558598 328046 558654 328102
rect 558722 328046 558778 328102
rect 558846 328046 558902 328102
rect 558474 327922 558530 327978
rect 558598 327922 558654 327978
rect 558722 327922 558778 327978
rect 558846 327922 558902 327978
rect 558474 310294 558530 310350
rect 558598 310294 558654 310350
rect 558722 310294 558778 310350
rect 558846 310294 558902 310350
rect 558474 310170 558530 310226
rect 558598 310170 558654 310226
rect 558722 310170 558778 310226
rect 558846 310170 558902 310226
rect 558474 310046 558530 310102
rect 558598 310046 558654 310102
rect 558722 310046 558778 310102
rect 558846 310046 558902 310102
rect 558474 309922 558530 309978
rect 558598 309922 558654 309978
rect 558722 309922 558778 309978
rect 558846 309922 558902 309978
rect 558474 292294 558530 292350
rect 558598 292294 558654 292350
rect 558722 292294 558778 292350
rect 558846 292294 558902 292350
rect 558474 292170 558530 292226
rect 558598 292170 558654 292226
rect 558722 292170 558778 292226
rect 558846 292170 558902 292226
rect 558474 292046 558530 292102
rect 558598 292046 558654 292102
rect 558722 292046 558778 292102
rect 558846 292046 558902 292102
rect 558474 291922 558530 291978
rect 558598 291922 558654 291978
rect 558722 291922 558778 291978
rect 558846 291922 558902 291978
rect 558474 274294 558530 274350
rect 558598 274294 558654 274350
rect 558722 274294 558778 274350
rect 558846 274294 558902 274350
rect 558474 274170 558530 274226
rect 558598 274170 558654 274226
rect 558722 274170 558778 274226
rect 558846 274170 558902 274226
rect 558474 274046 558530 274102
rect 558598 274046 558654 274102
rect 558722 274046 558778 274102
rect 558846 274046 558902 274102
rect 558474 273922 558530 273978
rect 558598 273922 558654 273978
rect 558722 273922 558778 273978
rect 558846 273922 558902 273978
rect 558474 256294 558530 256350
rect 558598 256294 558654 256350
rect 558722 256294 558778 256350
rect 558846 256294 558902 256350
rect 558474 256170 558530 256226
rect 558598 256170 558654 256226
rect 558722 256170 558778 256226
rect 558846 256170 558902 256226
rect 558474 256046 558530 256102
rect 558598 256046 558654 256102
rect 558722 256046 558778 256102
rect 558846 256046 558902 256102
rect 558474 255922 558530 255978
rect 558598 255922 558654 255978
rect 558722 255922 558778 255978
rect 558846 255922 558902 255978
rect 558474 238294 558530 238350
rect 558598 238294 558654 238350
rect 558722 238294 558778 238350
rect 558846 238294 558902 238350
rect 558474 238170 558530 238226
rect 558598 238170 558654 238226
rect 558722 238170 558778 238226
rect 558846 238170 558902 238226
rect 558474 238046 558530 238102
rect 558598 238046 558654 238102
rect 558722 238046 558778 238102
rect 558846 238046 558902 238102
rect 558474 237922 558530 237978
rect 558598 237922 558654 237978
rect 558722 237922 558778 237978
rect 558846 237922 558902 237978
rect 558474 220294 558530 220350
rect 558598 220294 558654 220350
rect 558722 220294 558778 220350
rect 558846 220294 558902 220350
rect 558474 220170 558530 220226
rect 558598 220170 558654 220226
rect 558722 220170 558778 220226
rect 558846 220170 558902 220226
rect 558474 220046 558530 220102
rect 558598 220046 558654 220102
rect 558722 220046 558778 220102
rect 558846 220046 558902 220102
rect 558474 219922 558530 219978
rect 558598 219922 558654 219978
rect 558722 219922 558778 219978
rect 558846 219922 558902 219978
rect 558474 202294 558530 202350
rect 558598 202294 558654 202350
rect 558722 202294 558778 202350
rect 558846 202294 558902 202350
rect 558474 202170 558530 202226
rect 558598 202170 558654 202226
rect 558722 202170 558778 202226
rect 558846 202170 558902 202226
rect 558474 202046 558530 202102
rect 558598 202046 558654 202102
rect 558722 202046 558778 202102
rect 558846 202046 558902 202102
rect 558474 201922 558530 201978
rect 558598 201922 558654 201978
rect 558722 201922 558778 201978
rect 558846 201922 558902 201978
rect 558474 184294 558530 184350
rect 558598 184294 558654 184350
rect 558722 184294 558778 184350
rect 558846 184294 558902 184350
rect 558474 184170 558530 184226
rect 558598 184170 558654 184226
rect 558722 184170 558778 184226
rect 558846 184170 558902 184226
rect 558474 184046 558530 184102
rect 558598 184046 558654 184102
rect 558722 184046 558778 184102
rect 558846 184046 558902 184102
rect 558474 183922 558530 183978
rect 558598 183922 558654 183978
rect 558722 183922 558778 183978
rect 558846 183922 558902 183978
rect 558474 166294 558530 166350
rect 558598 166294 558654 166350
rect 558722 166294 558778 166350
rect 558846 166294 558902 166350
rect 558474 166170 558530 166226
rect 558598 166170 558654 166226
rect 558722 166170 558778 166226
rect 558846 166170 558902 166226
rect 558474 166046 558530 166102
rect 558598 166046 558654 166102
rect 558722 166046 558778 166102
rect 558846 166046 558902 166102
rect 558474 165922 558530 165978
rect 558598 165922 558654 165978
rect 558722 165922 558778 165978
rect 558846 165922 558902 165978
rect 558474 148294 558530 148350
rect 558598 148294 558654 148350
rect 558722 148294 558778 148350
rect 558846 148294 558902 148350
rect 558474 148170 558530 148226
rect 558598 148170 558654 148226
rect 558722 148170 558778 148226
rect 558846 148170 558902 148226
rect 558474 148046 558530 148102
rect 558598 148046 558654 148102
rect 558722 148046 558778 148102
rect 558846 148046 558902 148102
rect 558474 147922 558530 147978
rect 558598 147922 558654 147978
rect 558722 147922 558778 147978
rect 558846 147922 558902 147978
rect 558474 130294 558530 130350
rect 558598 130294 558654 130350
rect 558722 130294 558778 130350
rect 558846 130294 558902 130350
rect 558474 130170 558530 130226
rect 558598 130170 558654 130226
rect 558722 130170 558778 130226
rect 558846 130170 558902 130226
rect 558474 130046 558530 130102
rect 558598 130046 558654 130102
rect 558722 130046 558778 130102
rect 558846 130046 558902 130102
rect 558474 129922 558530 129978
rect 558598 129922 558654 129978
rect 558722 129922 558778 129978
rect 558846 129922 558902 129978
rect 558474 112294 558530 112350
rect 558598 112294 558654 112350
rect 558722 112294 558778 112350
rect 558846 112294 558902 112350
rect 558474 112170 558530 112226
rect 558598 112170 558654 112226
rect 558722 112170 558778 112226
rect 558846 112170 558902 112226
rect 558474 112046 558530 112102
rect 558598 112046 558654 112102
rect 558722 112046 558778 112102
rect 558846 112046 558902 112102
rect 558474 111922 558530 111978
rect 558598 111922 558654 111978
rect 558722 111922 558778 111978
rect 558846 111922 558902 111978
rect 558474 94294 558530 94350
rect 558598 94294 558654 94350
rect 558722 94294 558778 94350
rect 558846 94294 558902 94350
rect 558474 94170 558530 94226
rect 558598 94170 558654 94226
rect 558722 94170 558778 94226
rect 558846 94170 558902 94226
rect 558474 94046 558530 94102
rect 558598 94046 558654 94102
rect 558722 94046 558778 94102
rect 558846 94046 558902 94102
rect 558474 93922 558530 93978
rect 558598 93922 558654 93978
rect 558722 93922 558778 93978
rect 558846 93922 558902 93978
rect 558474 76294 558530 76350
rect 558598 76294 558654 76350
rect 558722 76294 558778 76350
rect 558846 76294 558902 76350
rect 558474 76170 558530 76226
rect 558598 76170 558654 76226
rect 558722 76170 558778 76226
rect 558846 76170 558902 76226
rect 558474 76046 558530 76102
rect 558598 76046 558654 76102
rect 558722 76046 558778 76102
rect 558846 76046 558902 76102
rect 558474 75922 558530 75978
rect 558598 75922 558654 75978
rect 558722 75922 558778 75978
rect 558846 75922 558902 75978
rect 558474 58294 558530 58350
rect 558598 58294 558654 58350
rect 558722 58294 558778 58350
rect 558846 58294 558902 58350
rect 558474 58170 558530 58226
rect 558598 58170 558654 58226
rect 558722 58170 558778 58226
rect 558846 58170 558902 58226
rect 558474 58046 558530 58102
rect 558598 58046 558654 58102
rect 558722 58046 558778 58102
rect 558846 58046 558902 58102
rect 558474 57922 558530 57978
rect 558598 57922 558654 57978
rect 558722 57922 558778 57978
rect 558846 57922 558902 57978
rect 539308 57122 539364 57178
rect 534268 50642 534324 50698
rect 531474 46294 531530 46350
rect 531598 46294 531654 46350
rect 531722 46294 531778 46350
rect 531846 46294 531902 46350
rect 531474 46170 531530 46226
rect 531598 46170 531654 46226
rect 531722 46170 531778 46226
rect 531846 46170 531902 46226
rect 531474 46046 531530 46102
rect 531598 46046 531654 46102
rect 531722 46046 531778 46102
rect 531846 46046 531902 46102
rect 531474 45922 531530 45978
rect 531598 45922 531654 45978
rect 531722 45922 531778 45978
rect 531846 45922 531902 45978
rect 531474 28294 531530 28350
rect 531598 28294 531654 28350
rect 531722 28294 531778 28350
rect 531846 28294 531902 28350
rect 531474 28170 531530 28226
rect 531598 28170 531654 28226
rect 531722 28170 531778 28226
rect 531846 28170 531902 28226
rect 531474 28046 531530 28102
rect 531598 28046 531654 28102
rect 531722 28046 531778 28102
rect 531846 28046 531902 28102
rect 531474 27922 531530 27978
rect 531598 27922 531654 27978
rect 531722 27922 531778 27978
rect 531846 27922 531902 27978
rect 527754 4294 527810 4350
rect 527878 4294 527934 4350
rect 528002 4294 528058 4350
rect 528126 4294 528182 4350
rect 527754 4170 527810 4226
rect 527878 4170 527934 4226
rect 528002 4170 528058 4226
rect 528126 4170 528182 4226
rect 500754 -1176 500810 -1120
rect 500878 -1176 500934 -1120
rect 501002 -1176 501058 -1120
rect 501126 -1176 501182 -1120
rect 500754 -1300 500810 -1244
rect 500878 -1300 500934 -1244
rect 501002 -1300 501058 -1244
rect 501126 -1300 501182 -1244
rect 500754 -1424 500810 -1368
rect 500878 -1424 500934 -1368
rect 501002 -1424 501058 -1368
rect 501126 -1424 501182 -1368
rect 500754 -1548 500810 -1492
rect 500878 -1548 500934 -1492
rect 501002 -1548 501058 -1492
rect 501126 -1548 501182 -1492
rect 531132 15182 531188 15238
rect 531474 10294 531530 10350
rect 531598 10294 531654 10350
rect 531722 10294 531778 10350
rect 531846 10294 531902 10350
rect 531474 10170 531530 10226
rect 531598 10170 531654 10226
rect 531722 10170 531778 10226
rect 531846 10170 531902 10226
rect 531474 10046 531530 10102
rect 531598 10046 531654 10102
rect 531722 10046 531778 10102
rect 531846 10046 531902 10102
rect 531474 9922 531530 9978
rect 531598 9922 531654 9978
rect 531722 9922 531778 9978
rect 531846 9922 531902 9978
rect 527754 4046 527810 4102
rect 527878 4046 527934 4102
rect 528002 4046 528058 4102
rect 528126 4046 528182 4102
rect 527754 3922 527810 3978
rect 527878 3922 527934 3978
rect 528002 3922 528058 3978
rect 528126 3922 528182 3978
rect 527754 -216 527810 -160
rect 527878 -216 527934 -160
rect 528002 -216 528058 -160
rect 528126 -216 528182 -160
rect 527754 -340 527810 -284
rect 527878 -340 527934 -284
rect 528002 -340 528058 -284
rect 528126 -340 528182 -284
rect 527754 -464 527810 -408
rect 527878 -464 527934 -408
rect 528002 -464 528058 -408
rect 528126 -464 528182 -408
rect 527754 -588 527810 -532
rect 527878 -588 527934 -532
rect 528002 -588 528058 -532
rect 528126 -588 528182 -532
rect 532588 47042 532644 47098
rect 537628 50462 537684 50518
rect 554428 52082 554484 52138
rect 549388 48842 549444 48898
rect 544348 40562 544404 40618
rect 562194 598116 562250 598172
rect 562318 598116 562374 598172
rect 562442 598116 562498 598172
rect 562566 598116 562622 598172
rect 562194 597992 562250 598048
rect 562318 597992 562374 598048
rect 562442 597992 562498 598048
rect 562566 597992 562622 598048
rect 562194 597868 562250 597924
rect 562318 597868 562374 597924
rect 562442 597868 562498 597924
rect 562566 597868 562622 597924
rect 562194 597744 562250 597800
rect 562318 597744 562374 597800
rect 562442 597744 562498 597800
rect 562566 597744 562622 597800
rect 562194 586294 562250 586350
rect 562318 586294 562374 586350
rect 562442 586294 562498 586350
rect 562566 586294 562622 586350
rect 562194 586170 562250 586226
rect 562318 586170 562374 586226
rect 562442 586170 562498 586226
rect 562566 586170 562622 586226
rect 562194 586046 562250 586102
rect 562318 586046 562374 586102
rect 562442 586046 562498 586102
rect 562566 586046 562622 586102
rect 562194 585922 562250 585978
rect 562318 585922 562374 585978
rect 562442 585922 562498 585978
rect 562566 585922 562622 585978
rect 562194 568294 562250 568350
rect 562318 568294 562374 568350
rect 562442 568294 562498 568350
rect 562566 568294 562622 568350
rect 562194 568170 562250 568226
rect 562318 568170 562374 568226
rect 562442 568170 562498 568226
rect 562566 568170 562622 568226
rect 562194 568046 562250 568102
rect 562318 568046 562374 568102
rect 562442 568046 562498 568102
rect 562566 568046 562622 568102
rect 562194 567922 562250 567978
rect 562318 567922 562374 567978
rect 562442 567922 562498 567978
rect 562566 567922 562622 567978
rect 562194 550294 562250 550350
rect 562318 550294 562374 550350
rect 562442 550294 562498 550350
rect 562566 550294 562622 550350
rect 562194 550170 562250 550226
rect 562318 550170 562374 550226
rect 562442 550170 562498 550226
rect 562566 550170 562622 550226
rect 562194 550046 562250 550102
rect 562318 550046 562374 550102
rect 562442 550046 562498 550102
rect 562566 550046 562622 550102
rect 562194 549922 562250 549978
rect 562318 549922 562374 549978
rect 562442 549922 562498 549978
rect 562566 549922 562622 549978
rect 562194 532294 562250 532350
rect 562318 532294 562374 532350
rect 562442 532294 562498 532350
rect 562566 532294 562622 532350
rect 562194 532170 562250 532226
rect 562318 532170 562374 532226
rect 562442 532170 562498 532226
rect 562566 532170 562622 532226
rect 562194 532046 562250 532102
rect 562318 532046 562374 532102
rect 562442 532046 562498 532102
rect 562566 532046 562622 532102
rect 562194 531922 562250 531978
rect 562318 531922 562374 531978
rect 562442 531922 562498 531978
rect 562566 531922 562622 531978
rect 562194 514294 562250 514350
rect 562318 514294 562374 514350
rect 562442 514294 562498 514350
rect 562566 514294 562622 514350
rect 562194 514170 562250 514226
rect 562318 514170 562374 514226
rect 562442 514170 562498 514226
rect 562566 514170 562622 514226
rect 562194 514046 562250 514102
rect 562318 514046 562374 514102
rect 562442 514046 562498 514102
rect 562566 514046 562622 514102
rect 562194 513922 562250 513978
rect 562318 513922 562374 513978
rect 562442 513922 562498 513978
rect 562566 513922 562622 513978
rect 562194 496294 562250 496350
rect 562318 496294 562374 496350
rect 562442 496294 562498 496350
rect 562566 496294 562622 496350
rect 562194 496170 562250 496226
rect 562318 496170 562374 496226
rect 562442 496170 562498 496226
rect 562566 496170 562622 496226
rect 562194 496046 562250 496102
rect 562318 496046 562374 496102
rect 562442 496046 562498 496102
rect 562566 496046 562622 496102
rect 562194 495922 562250 495978
rect 562318 495922 562374 495978
rect 562442 495922 562498 495978
rect 562566 495922 562622 495978
rect 562194 478294 562250 478350
rect 562318 478294 562374 478350
rect 562442 478294 562498 478350
rect 562566 478294 562622 478350
rect 562194 478170 562250 478226
rect 562318 478170 562374 478226
rect 562442 478170 562498 478226
rect 562566 478170 562622 478226
rect 562194 478046 562250 478102
rect 562318 478046 562374 478102
rect 562442 478046 562498 478102
rect 562566 478046 562622 478102
rect 562194 477922 562250 477978
rect 562318 477922 562374 477978
rect 562442 477922 562498 477978
rect 562566 477922 562622 477978
rect 562194 460294 562250 460350
rect 562318 460294 562374 460350
rect 562442 460294 562498 460350
rect 562566 460294 562622 460350
rect 562194 460170 562250 460226
rect 562318 460170 562374 460226
rect 562442 460170 562498 460226
rect 562566 460170 562622 460226
rect 562194 460046 562250 460102
rect 562318 460046 562374 460102
rect 562442 460046 562498 460102
rect 562566 460046 562622 460102
rect 562194 459922 562250 459978
rect 562318 459922 562374 459978
rect 562442 459922 562498 459978
rect 562566 459922 562622 459978
rect 562194 442294 562250 442350
rect 562318 442294 562374 442350
rect 562442 442294 562498 442350
rect 562566 442294 562622 442350
rect 562194 442170 562250 442226
rect 562318 442170 562374 442226
rect 562442 442170 562498 442226
rect 562566 442170 562622 442226
rect 562194 442046 562250 442102
rect 562318 442046 562374 442102
rect 562442 442046 562498 442102
rect 562566 442046 562622 442102
rect 562194 441922 562250 441978
rect 562318 441922 562374 441978
rect 562442 441922 562498 441978
rect 562566 441922 562622 441978
rect 562194 424294 562250 424350
rect 562318 424294 562374 424350
rect 562442 424294 562498 424350
rect 562566 424294 562622 424350
rect 562194 424170 562250 424226
rect 562318 424170 562374 424226
rect 562442 424170 562498 424226
rect 562566 424170 562622 424226
rect 562194 424046 562250 424102
rect 562318 424046 562374 424102
rect 562442 424046 562498 424102
rect 562566 424046 562622 424102
rect 562194 423922 562250 423978
rect 562318 423922 562374 423978
rect 562442 423922 562498 423978
rect 562566 423922 562622 423978
rect 562194 406294 562250 406350
rect 562318 406294 562374 406350
rect 562442 406294 562498 406350
rect 562566 406294 562622 406350
rect 562194 406170 562250 406226
rect 562318 406170 562374 406226
rect 562442 406170 562498 406226
rect 562566 406170 562622 406226
rect 562194 406046 562250 406102
rect 562318 406046 562374 406102
rect 562442 406046 562498 406102
rect 562566 406046 562622 406102
rect 562194 405922 562250 405978
rect 562318 405922 562374 405978
rect 562442 405922 562498 405978
rect 562566 405922 562622 405978
rect 562194 388294 562250 388350
rect 562318 388294 562374 388350
rect 562442 388294 562498 388350
rect 562566 388294 562622 388350
rect 562194 388170 562250 388226
rect 562318 388170 562374 388226
rect 562442 388170 562498 388226
rect 562566 388170 562622 388226
rect 562194 388046 562250 388102
rect 562318 388046 562374 388102
rect 562442 388046 562498 388102
rect 562566 388046 562622 388102
rect 562194 387922 562250 387978
rect 562318 387922 562374 387978
rect 562442 387922 562498 387978
rect 562566 387922 562622 387978
rect 562194 370294 562250 370350
rect 562318 370294 562374 370350
rect 562442 370294 562498 370350
rect 562566 370294 562622 370350
rect 562194 370170 562250 370226
rect 562318 370170 562374 370226
rect 562442 370170 562498 370226
rect 562566 370170 562622 370226
rect 562194 370046 562250 370102
rect 562318 370046 562374 370102
rect 562442 370046 562498 370102
rect 562566 370046 562622 370102
rect 562194 369922 562250 369978
rect 562318 369922 562374 369978
rect 562442 369922 562498 369978
rect 562566 369922 562622 369978
rect 589194 597156 589250 597212
rect 589318 597156 589374 597212
rect 589442 597156 589498 597212
rect 589566 597156 589622 597212
rect 589194 597032 589250 597088
rect 589318 597032 589374 597088
rect 589442 597032 589498 597088
rect 589566 597032 589622 597088
rect 589194 596908 589250 596964
rect 589318 596908 589374 596964
rect 589442 596908 589498 596964
rect 589566 596908 589622 596964
rect 589194 596784 589250 596840
rect 589318 596784 589374 596840
rect 589442 596784 589498 596840
rect 589566 596784 589622 596840
rect 589194 580294 589250 580350
rect 589318 580294 589374 580350
rect 589442 580294 589498 580350
rect 589566 580294 589622 580350
rect 589194 580170 589250 580226
rect 589318 580170 589374 580226
rect 589442 580170 589498 580226
rect 589566 580170 589622 580226
rect 589194 580046 589250 580102
rect 589318 580046 589374 580102
rect 589442 580046 589498 580102
rect 589566 580046 589622 580102
rect 589194 579922 589250 579978
rect 589318 579922 589374 579978
rect 589442 579922 589498 579978
rect 589566 579922 589622 579978
rect 589194 562294 589250 562350
rect 589318 562294 589374 562350
rect 589442 562294 589498 562350
rect 589566 562294 589622 562350
rect 589194 562170 589250 562226
rect 589318 562170 589374 562226
rect 589442 562170 589498 562226
rect 589566 562170 589622 562226
rect 592914 598116 592970 598172
rect 593038 598116 593094 598172
rect 593162 598116 593218 598172
rect 593286 598116 593342 598172
rect 592914 597992 592970 598048
rect 593038 597992 593094 598048
rect 593162 597992 593218 598048
rect 593286 597992 593342 598048
rect 592914 597868 592970 597924
rect 593038 597868 593094 597924
rect 593162 597868 593218 597924
rect 593286 597868 593342 597924
rect 592914 597744 592970 597800
rect 593038 597744 593094 597800
rect 593162 597744 593218 597800
rect 593286 597744 593342 597800
rect 597456 598116 597512 598172
rect 597580 598116 597636 598172
rect 597704 598116 597760 598172
rect 597828 598116 597884 598172
rect 597456 597992 597512 598048
rect 597580 597992 597636 598048
rect 597704 597992 597760 598048
rect 597828 597992 597884 598048
rect 597456 597868 597512 597924
rect 597580 597868 597636 597924
rect 597704 597868 597760 597924
rect 597828 597868 597884 597924
rect 597456 597744 597512 597800
rect 597580 597744 597636 597800
rect 597704 597744 597760 597800
rect 597828 597744 597884 597800
rect 592914 586294 592970 586350
rect 593038 586294 593094 586350
rect 593162 586294 593218 586350
rect 593286 586294 593342 586350
rect 592914 586170 592970 586226
rect 593038 586170 593094 586226
rect 593162 586170 593218 586226
rect 593286 586170 593342 586226
rect 592914 586046 592970 586102
rect 593038 586046 593094 586102
rect 593162 586046 593218 586102
rect 593286 586046 593342 586102
rect 592914 585922 592970 585978
rect 593038 585922 593094 585978
rect 593162 585922 593218 585978
rect 593286 585922 593342 585978
rect 592914 568294 592970 568350
rect 593038 568294 593094 568350
rect 593162 568294 593218 568350
rect 593286 568294 593342 568350
rect 592914 568170 592970 568226
rect 593038 568170 593094 568226
rect 593162 568170 593218 568226
rect 593286 568170 593342 568226
rect 592914 568046 592970 568102
rect 593038 568046 593094 568102
rect 593162 568046 593218 568102
rect 593286 568046 593342 568102
rect 592914 567922 592970 567978
rect 593038 567922 593094 567978
rect 593162 567922 593218 567978
rect 593286 567922 593342 567978
rect 589194 562046 589250 562102
rect 589318 562046 589374 562102
rect 589442 562046 589498 562102
rect 589566 562046 589622 562102
rect 589194 561922 589250 561978
rect 589318 561922 589374 561978
rect 589442 561922 589498 561978
rect 589566 561922 589622 561978
rect 589194 544294 589250 544350
rect 589318 544294 589374 544350
rect 589442 544294 589498 544350
rect 589566 544294 589622 544350
rect 589194 544170 589250 544226
rect 589318 544170 589374 544226
rect 589442 544170 589498 544226
rect 589566 544170 589622 544226
rect 589194 544046 589250 544102
rect 589318 544046 589374 544102
rect 589442 544046 589498 544102
rect 589566 544046 589622 544102
rect 589194 543922 589250 543978
rect 589318 543922 589374 543978
rect 589442 543922 589498 543978
rect 589566 543922 589622 543978
rect 589194 526294 589250 526350
rect 589318 526294 589374 526350
rect 589442 526294 589498 526350
rect 589566 526294 589622 526350
rect 589194 526170 589250 526226
rect 589318 526170 589374 526226
rect 589442 526170 589498 526226
rect 589566 526170 589622 526226
rect 589194 526046 589250 526102
rect 589318 526046 589374 526102
rect 589442 526046 589498 526102
rect 589566 526046 589622 526102
rect 589194 525922 589250 525978
rect 589318 525922 589374 525978
rect 589442 525922 589498 525978
rect 589566 525922 589622 525978
rect 592914 550294 592970 550350
rect 593038 550294 593094 550350
rect 593162 550294 593218 550350
rect 593286 550294 593342 550350
rect 592914 550170 592970 550226
rect 593038 550170 593094 550226
rect 593162 550170 593218 550226
rect 593286 550170 593342 550226
rect 592914 550046 592970 550102
rect 593038 550046 593094 550102
rect 593162 550046 593218 550102
rect 593286 550046 593342 550102
rect 592914 549922 592970 549978
rect 593038 549922 593094 549978
rect 593162 549922 593218 549978
rect 593286 549922 593342 549978
rect 592914 532294 592970 532350
rect 593038 532294 593094 532350
rect 593162 532294 593218 532350
rect 593286 532294 593342 532350
rect 592914 532170 592970 532226
rect 593038 532170 593094 532226
rect 593162 532170 593218 532226
rect 593286 532170 593342 532226
rect 592914 532046 592970 532102
rect 593038 532046 593094 532102
rect 593162 532046 593218 532102
rect 593286 532046 593342 532102
rect 592914 531922 592970 531978
rect 593038 531922 593094 531978
rect 593162 531922 593218 531978
rect 593286 531922 593342 531978
rect 589194 508294 589250 508350
rect 589318 508294 589374 508350
rect 589442 508294 589498 508350
rect 589566 508294 589622 508350
rect 589194 508170 589250 508226
rect 589318 508170 589374 508226
rect 589442 508170 589498 508226
rect 589566 508170 589622 508226
rect 589194 508046 589250 508102
rect 589318 508046 589374 508102
rect 589442 508046 589498 508102
rect 589566 508046 589622 508102
rect 589194 507922 589250 507978
rect 589318 507922 589374 507978
rect 589442 507922 589498 507978
rect 589566 507922 589622 507978
rect 589194 490294 589250 490350
rect 589318 490294 589374 490350
rect 589442 490294 589498 490350
rect 589566 490294 589622 490350
rect 589194 490170 589250 490226
rect 589318 490170 589374 490226
rect 589442 490170 589498 490226
rect 589566 490170 589622 490226
rect 589194 490046 589250 490102
rect 589318 490046 589374 490102
rect 589442 490046 589498 490102
rect 589566 490046 589622 490102
rect 589194 489922 589250 489978
rect 589318 489922 589374 489978
rect 589442 489922 589498 489978
rect 589566 489922 589622 489978
rect 589194 472294 589250 472350
rect 589318 472294 589374 472350
rect 589442 472294 589498 472350
rect 589566 472294 589622 472350
rect 589194 472170 589250 472226
rect 589318 472170 589374 472226
rect 589442 472170 589498 472226
rect 589566 472170 589622 472226
rect 589194 472046 589250 472102
rect 589318 472046 589374 472102
rect 589442 472046 589498 472102
rect 589566 472046 589622 472102
rect 589194 471922 589250 471978
rect 589318 471922 589374 471978
rect 589442 471922 589498 471978
rect 589566 471922 589622 471978
rect 589194 454294 589250 454350
rect 589318 454294 589374 454350
rect 589442 454294 589498 454350
rect 589566 454294 589622 454350
rect 589194 454170 589250 454226
rect 589318 454170 589374 454226
rect 589442 454170 589498 454226
rect 589566 454170 589622 454226
rect 589194 454046 589250 454102
rect 589318 454046 589374 454102
rect 589442 454046 589498 454102
rect 589566 454046 589622 454102
rect 589194 453922 589250 453978
rect 589318 453922 589374 453978
rect 589442 453922 589498 453978
rect 589566 453922 589622 453978
rect 589194 436294 589250 436350
rect 589318 436294 589374 436350
rect 589442 436294 589498 436350
rect 589566 436294 589622 436350
rect 589194 436170 589250 436226
rect 589318 436170 589374 436226
rect 589442 436170 589498 436226
rect 589566 436170 589622 436226
rect 589194 436046 589250 436102
rect 589318 436046 589374 436102
rect 589442 436046 589498 436102
rect 589566 436046 589622 436102
rect 589194 435922 589250 435978
rect 589318 435922 589374 435978
rect 589442 435922 589498 435978
rect 589566 435922 589622 435978
rect 589194 418294 589250 418350
rect 589318 418294 589374 418350
rect 589442 418294 589498 418350
rect 589566 418294 589622 418350
rect 589194 418170 589250 418226
rect 589318 418170 589374 418226
rect 589442 418170 589498 418226
rect 589566 418170 589622 418226
rect 589194 418046 589250 418102
rect 589318 418046 589374 418102
rect 589442 418046 589498 418102
rect 589566 418046 589622 418102
rect 589194 417922 589250 417978
rect 589318 417922 589374 417978
rect 589442 417922 589498 417978
rect 589566 417922 589622 417978
rect 589194 400294 589250 400350
rect 589318 400294 589374 400350
rect 589442 400294 589498 400350
rect 589566 400294 589622 400350
rect 589194 400170 589250 400226
rect 589318 400170 589374 400226
rect 589442 400170 589498 400226
rect 589566 400170 589622 400226
rect 589194 400046 589250 400102
rect 589318 400046 589374 400102
rect 589442 400046 589498 400102
rect 589566 400046 589622 400102
rect 589194 399922 589250 399978
rect 589318 399922 589374 399978
rect 589442 399922 589498 399978
rect 589566 399922 589622 399978
rect 589194 382294 589250 382350
rect 589318 382294 589374 382350
rect 589442 382294 589498 382350
rect 589566 382294 589622 382350
rect 589194 382170 589250 382226
rect 589318 382170 589374 382226
rect 589442 382170 589498 382226
rect 589566 382170 589622 382226
rect 589194 382046 589250 382102
rect 589318 382046 589374 382102
rect 589442 382046 589498 382102
rect 589566 382046 589622 382102
rect 589194 381922 589250 381978
rect 589318 381922 589374 381978
rect 589442 381922 589498 381978
rect 589566 381922 589622 381978
rect 589194 364294 589250 364350
rect 589318 364294 589374 364350
rect 589442 364294 589498 364350
rect 589566 364294 589622 364350
rect 589194 364170 589250 364226
rect 589318 364170 589374 364226
rect 589442 364170 589498 364226
rect 589566 364170 589622 364226
rect 589194 364046 589250 364102
rect 589318 364046 589374 364102
rect 589442 364046 589498 364102
rect 589566 364046 589622 364102
rect 562194 352294 562250 352350
rect 562318 352294 562374 352350
rect 562442 352294 562498 352350
rect 562566 352294 562622 352350
rect 562194 352170 562250 352226
rect 562318 352170 562374 352226
rect 562442 352170 562498 352226
rect 562566 352170 562622 352226
rect 562194 352046 562250 352102
rect 562318 352046 562374 352102
rect 562442 352046 562498 352102
rect 562566 352046 562622 352102
rect 562194 351922 562250 351978
rect 562318 351922 562374 351978
rect 562442 351922 562498 351978
rect 562566 351922 562622 351978
rect 562194 334294 562250 334350
rect 562318 334294 562374 334350
rect 562442 334294 562498 334350
rect 562566 334294 562622 334350
rect 562194 334170 562250 334226
rect 562318 334170 562374 334226
rect 562442 334170 562498 334226
rect 562566 334170 562622 334226
rect 562194 334046 562250 334102
rect 562318 334046 562374 334102
rect 562442 334046 562498 334102
rect 562566 334046 562622 334102
rect 562194 333922 562250 333978
rect 562318 333922 562374 333978
rect 562442 333922 562498 333978
rect 562566 333922 562622 333978
rect 562194 316294 562250 316350
rect 562318 316294 562374 316350
rect 562442 316294 562498 316350
rect 562566 316294 562622 316350
rect 562194 316170 562250 316226
rect 562318 316170 562374 316226
rect 562442 316170 562498 316226
rect 562566 316170 562622 316226
rect 562194 316046 562250 316102
rect 562318 316046 562374 316102
rect 562442 316046 562498 316102
rect 562566 316046 562622 316102
rect 562194 315922 562250 315978
rect 562318 315922 562374 315978
rect 562442 315922 562498 315978
rect 562566 315922 562622 315978
rect 562194 298294 562250 298350
rect 562318 298294 562374 298350
rect 562442 298294 562498 298350
rect 562566 298294 562622 298350
rect 562194 298170 562250 298226
rect 562318 298170 562374 298226
rect 562442 298170 562498 298226
rect 562566 298170 562622 298226
rect 562194 298046 562250 298102
rect 562318 298046 562374 298102
rect 562442 298046 562498 298102
rect 562566 298046 562622 298102
rect 562194 297922 562250 297978
rect 562318 297922 562374 297978
rect 562442 297922 562498 297978
rect 562566 297922 562622 297978
rect 562194 280294 562250 280350
rect 562318 280294 562374 280350
rect 562442 280294 562498 280350
rect 562566 280294 562622 280350
rect 562194 280170 562250 280226
rect 562318 280170 562374 280226
rect 562442 280170 562498 280226
rect 562566 280170 562622 280226
rect 562194 280046 562250 280102
rect 562318 280046 562374 280102
rect 562442 280046 562498 280102
rect 562566 280046 562622 280102
rect 562194 279922 562250 279978
rect 562318 279922 562374 279978
rect 562442 279922 562498 279978
rect 562566 279922 562622 279978
rect 562194 262294 562250 262350
rect 562318 262294 562374 262350
rect 562442 262294 562498 262350
rect 562566 262294 562622 262350
rect 562194 262170 562250 262226
rect 562318 262170 562374 262226
rect 562442 262170 562498 262226
rect 562566 262170 562622 262226
rect 562194 262046 562250 262102
rect 562318 262046 562374 262102
rect 562442 262046 562498 262102
rect 562566 262046 562622 262102
rect 562194 261922 562250 261978
rect 562318 261922 562374 261978
rect 562442 261922 562498 261978
rect 562566 261922 562622 261978
rect 562194 244294 562250 244350
rect 562318 244294 562374 244350
rect 562442 244294 562498 244350
rect 562566 244294 562622 244350
rect 562194 244170 562250 244226
rect 562318 244170 562374 244226
rect 562442 244170 562498 244226
rect 562566 244170 562622 244226
rect 562194 244046 562250 244102
rect 562318 244046 562374 244102
rect 562442 244046 562498 244102
rect 562566 244046 562622 244102
rect 562194 243922 562250 243978
rect 562318 243922 562374 243978
rect 562442 243922 562498 243978
rect 562566 243922 562622 243978
rect 562194 226294 562250 226350
rect 562318 226294 562374 226350
rect 562442 226294 562498 226350
rect 562566 226294 562622 226350
rect 562194 226170 562250 226226
rect 562318 226170 562374 226226
rect 562442 226170 562498 226226
rect 562566 226170 562622 226226
rect 562194 226046 562250 226102
rect 562318 226046 562374 226102
rect 562442 226046 562498 226102
rect 562566 226046 562622 226102
rect 562194 225922 562250 225978
rect 562318 225922 562374 225978
rect 562442 225922 562498 225978
rect 562566 225922 562622 225978
rect 562194 208294 562250 208350
rect 562318 208294 562374 208350
rect 562442 208294 562498 208350
rect 562566 208294 562622 208350
rect 562194 208170 562250 208226
rect 562318 208170 562374 208226
rect 562442 208170 562498 208226
rect 562566 208170 562622 208226
rect 562194 208046 562250 208102
rect 562318 208046 562374 208102
rect 562442 208046 562498 208102
rect 562566 208046 562622 208102
rect 562194 207922 562250 207978
rect 562318 207922 562374 207978
rect 562442 207922 562498 207978
rect 562566 207922 562622 207978
rect 562194 190294 562250 190350
rect 562318 190294 562374 190350
rect 562442 190294 562498 190350
rect 562566 190294 562622 190350
rect 562194 190170 562250 190226
rect 562318 190170 562374 190226
rect 562442 190170 562498 190226
rect 562566 190170 562622 190226
rect 562194 190046 562250 190102
rect 562318 190046 562374 190102
rect 562442 190046 562498 190102
rect 562566 190046 562622 190102
rect 562194 189922 562250 189978
rect 562318 189922 562374 189978
rect 562442 189922 562498 189978
rect 562566 189922 562622 189978
rect 562194 172294 562250 172350
rect 562318 172294 562374 172350
rect 562442 172294 562498 172350
rect 562566 172294 562622 172350
rect 562194 172170 562250 172226
rect 562318 172170 562374 172226
rect 562442 172170 562498 172226
rect 562566 172170 562622 172226
rect 562194 172046 562250 172102
rect 562318 172046 562374 172102
rect 562442 172046 562498 172102
rect 562566 172046 562622 172102
rect 562194 171922 562250 171978
rect 562318 171922 562374 171978
rect 562442 171922 562498 171978
rect 562566 171922 562622 171978
rect 562194 154294 562250 154350
rect 562318 154294 562374 154350
rect 562442 154294 562498 154350
rect 562566 154294 562622 154350
rect 562194 154170 562250 154226
rect 562318 154170 562374 154226
rect 562442 154170 562498 154226
rect 562566 154170 562622 154226
rect 562194 154046 562250 154102
rect 562318 154046 562374 154102
rect 562442 154046 562498 154102
rect 562566 154046 562622 154102
rect 562194 153922 562250 153978
rect 562318 153922 562374 153978
rect 562442 153922 562498 153978
rect 562566 153922 562622 153978
rect 562194 136294 562250 136350
rect 562318 136294 562374 136350
rect 562442 136294 562498 136350
rect 562566 136294 562622 136350
rect 562194 136170 562250 136226
rect 562318 136170 562374 136226
rect 562442 136170 562498 136226
rect 562566 136170 562622 136226
rect 562194 136046 562250 136102
rect 562318 136046 562374 136102
rect 562442 136046 562498 136102
rect 562566 136046 562622 136102
rect 562194 135922 562250 135978
rect 562318 135922 562374 135978
rect 562442 135922 562498 135978
rect 562566 135922 562622 135978
rect 562194 118294 562250 118350
rect 562318 118294 562374 118350
rect 562442 118294 562498 118350
rect 562566 118294 562622 118350
rect 562194 118170 562250 118226
rect 562318 118170 562374 118226
rect 562442 118170 562498 118226
rect 562566 118170 562622 118226
rect 562194 118046 562250 118102
rect 562318 118046 562374 118102
rect 562442 118046 562498 118102
rect 562566 118046 562622 118102
rect 562194 117922 562250 117978
rect 562318 117922 562374 117978
rect 562442 117922 562498 117978
rect 562566 117922 562622 117978
rect 589194 363922 589250 363978
rect 589318 363922 589374 363978
rect 589442 363922 589498 363978
rect 589566 363922 589622 363978
rect 589194 346294 589250 346350
rect 589318 346294 589374 346350
rect 589442 346294 589498 346350
rect 589566 346294 589622 346350
rect 589194 346170 589250 346226
rect 589318 346170 589374 346226
rect 589442 346170 589498 346226
rect 589566 346170 589622 346226
rect 589194 346046 589250 346102
rect 589318 346046 589374 346102
rect 589442 346046 589498 346102
rect 589566 346046 589622 346102
rect 589194 345922 589250 345978
rect 589318 345922 589374 345978
rect 589442 345922 589498 345978
rect 589566 345922 589622 345978
rect 589194 328294 589250 328350
rect 589318 328294 589374 328350
rect 589442 328294 589498 328350
rect 589566 328294 589622 328350
rect 589194 328170 589250 328226
rect 589318 328170 589374 328226
rect 589442 328170 589498 328226
rect 589566 328170 589622 328226
rect 589194 328046 589250 328102
rect 589318 328046 589374 328102
rect 589442 328046 589498 328102
rect 589566 328046 589622 328102
rect 589194 327922 589250 327978
rect 589318 327922 589374 327978
rect 589442 327922 589498 327978
rect 589566 327922 589622 327978
rect 589194 310294 589250 310350
rect 589318 310294 589374 310350
rect 589442 310294 589498 310350
rect 589566 310294 589622 310350
rect 589194 310170 589250 310226
rect 589318 310170 589374 310226
rect 589442 310170 589498 310226
rect 589566 310170 589622 310226
rect 589194 310046 589250 310102
rect 589318 310046 589374 310102
rect 589442 310046 589498 310102
rect 589566 310046 589622 310102
rect 589194 309922 589250 309978
rect 589318 309922 589374 309978
rect 589442 309922 589498 309978
rect 589566 309922 589622 309978
rect 589194 292294 589250 292350
rect 589318 292294 589374 292350
rect 589442 292294 589498 292350
rect 589566 292294 589622 292350
rect 589194 292170 589250 292226
rect 589318 292170 589374 292226
rect 589442 292170 589498 292226
rect 589566 292170 589622 292226
rect 589194 292046 589250 292102
rect 589318 292046 589374 292102
rect 589442 292046 589498 292102
rect 589566 292046 589622 292102
rect 589194 291922 589250 291978
rect 589318 291922 589374 291978
rect 589442 291922 589498 291978
rect 589566 291922 589622 291978
rect 589194 274294 589250 274350
rect 589318 274294 589374 274350
rect 589442 274294 589498 274350
rect 589566 274294 589622 274350
rect 589194 274170 589250 274226
rect 589318 274170 589374 274226
rect 589442 274170 589498 274226
rect 589566 274170 589622 274226
rect 589194 274046 589250 274102
rect 589318 274046 589374 274102
rect 589442 274046 589498 274102
rect 589566 274046 589622 274102
rect 589194 273922 589250 273978
rect 589318 273922 589374 273978
rect 589442 273922 589498 273978
rect 589566 273922 589622 273978
rect 589194 256294 589250 256350
rect 589318 256294 589374 256350
rect 589442 256294 589498 256350
rect 589566 256294 589622 256350
rect 589194 256170 589250 256226
rect 589318 256170 589374 256226
rect 589442 256170 589498 256226
rect 589566 256170 589622 256226
rect 589194 256046 589250 256102
rect 589318 256046 589374 256102
rect 589442 256046 589498 256102
rect 589566 256046 589622 256102
rect 589194 255922 589250 255978
rect 589318 255922 589374 255978
rect 589442 255922 589498 255978
rect 589566 255922 589622 255978
rect 589194 238294 589250 238350
rect 589318 238294 589374 238350
rect 589442 238294 589498 238350
rect 589566 238294 589622 238350
rect 589194 238170 589250 238226
rect 589318 238170 589374 238226
rect 589442 238170 589498 238226
rect 589566 238170 589622 238226
rect 589194 238046 589250 238102
rect 589318 238046 589374 238102
rect 589442 238046 589498 238102
rect 589566 238046 589622 238102
rect 589194 237922 589250 237978
rect 589318 237922 589374 237978
rect 589442 237922 589498 237978
rect 589566 237922 589622 237978
rect 589194 220294 589250 220350
rect 589318 220294 589374 220350
rect 589442 220294 589498 220350
rect 589566 220294 589622 220350
rect 589194 220170 589250 220226
rect 589318 220170 589374 220226
rect 589442 220170 589498 220226
rect 589566 220170 589622 220226
rect 589194 220046 589250 220102
rect 589318 220046 589374 220102
rect 589442 220046 589498 220102
rect 589566 220046 589622 220102
rect 589194 219922 589250 219978
rect 589318 219922 589374 219978
rect 589442 219922 589498 219978
rect 589566 219922 589622 219978
rect 589194 202294 589250 202350
rect 589318 202294 589374 202350
rect 589442 202294 589498 202350
rect 589566 202294 589622 202350
rect 589194 202170 589250 202226
rect 589318 202170 589374 202226
rect 589442 202170 589498 202226
rect 589566 202170 589622 202226
rect 589194 202046 589250 202102
rect 589318 202046 589374 202102
rect 589442 202046 589498 202102
rect 589566 202046 589622 202102
rect 589194 201922 589250 201978
rect 589318 201922 589374 201978
rect 589442 201922 589498 201978
rect 589566 201922 589622 201978
rect 589194 184294 589250 184350
rect 589318 184294 589374 184350
rect 589442 184294 589498 184350
rect 589566 184294 589622 184350
rect 589194 184170 589250 184226
rect 589318 184170 589374 184226
rect 589442 184170 589498 184226
rect 589566 184170 589622 184226
rect 589194 184046 589250 184102
rect 589318 184046 589374 184102
rect 589442 184046 589498 184102
rect 589566 184046 589622 184102
rect 589194 183922 589250 183978
rect 589318 183922 589374 183978
rect 589442 183922 589498 183978
rect 589566 183922 589622 183978
rect 589194 166294 589250 166350
rect 589318 166294 589374 166350
rect 589442 166294 589498 166350
rect 589566 166294 589622 166350
rect 589194 166170 589250 166226
rect 589318 166170 589374 166226
rect 589442 166170 589498 166226
rect 589566 166170 589622 166226
rect 589194 166046 589250 166102
rect 589318 166046 589374 166102
rect 589442 166046 589498 166102
rect 589566 166046 589622 166102
rect 589194 165922 589250 165978
rect 589318 165922 589374 165978
rect 589442 165922 589498 165978
rect 589566 165922 589622 165978
rect 589194 148294 589250 148350
rect 589318 148294 589374 148350
rect 589442 148294 589498 148350
rect 589566 148294 589622 148350
rect 589194 148170 589250 148226
rect 589318 148170 589374 148226
rect 589442 148170 589498 148226
rect 589566 148170 589622 148226
rect 589194 148046 589250 148102
rect 589318 148046 589374 148102
rect 589442 148046 589498 148102
rect 589566 148046 589622 148102
rect 589194 147922 589250 147978
rect 589318 147922 589374 147978
rect 589442 147922 589498 147978
rect 589566 147922 589622 147978
rect 589194 130294 589250 130350
rect 589318 130294 589374 130350
rect 589442 130294 589498 130350
rect 589566 130294 589622 130350
rect 589194 130170 589250 130226
rect 589318 130170 589374 130226
rect 589442 130170 589498 130226
rect 589566 130170 589622 130226
rect 589194 130046 589250 130102
rect 589318 130046 589374 130102
rect 589442 130046 589498 130102
rect 589566 130046 589622 130102
rect 589194 129922 589250 129978
rect 589318 129922 589374 129978
rect 589442 129922 589498 129978
rect 589566 129922 589622 129978
rect 589194 112294 589250 112350
rect 589318 112294 589374 112350
rect 589442 112294 589498 112350
rect 589566 112294 589622 112350
rect 589194 112170 589250 112226
rect 589318 112170 589374 112226
rect 589442 112170 589498 112226
rect 589566 112170 589622 112226
rect 589194 112046 589250 112102
rect 589318 112046 589374 112102
rect 589442 112046 589498 112102
rect 589566 112046 589622 112102
rect 589194 111922 589250 111978
rect 589318 111922 589374 111978
rect 589442 111922 589498 111978
rect 589566 111922 589622 111978
rect 562194 100294 562250 100350
rect 562318 100294 562374 100350
rect 562442 100294 562498 100350
rect 562566 100294 562622 100350
rect 562194 100170 562250 100226
rect 562318 100170 562374 100226
rect 562442 100170 562498 100226
rect 562566 100170 562622 100226
rect 562194 100046 562250 100102
rect 562318 100046 562374 100102
rect 562442 100046 562498 100102
rect 562566 100046 562622 100102
rect 562194 99922 562250 99978
rect 562318 99922 562374 99978
rect 562442 99922 562498 99978
rect 562566 99922 562622 99978
rect 562194 82294 562250 82350
rect 562318 82294 562374 82350
rect 562442 82294 562498 82350
rect 562566 82294 562622 82350
rect 562194 82170 562250 82226
rect 562318 82170 562374 82226
rect 562442 82170 562498 82226
rect 562566 82170 562622 82226
rect 562194 82046 562250 82102
rect 562318 82046 562374 82102
rect 562442 82046 562498 82102
rect 562566 82046 562622 82102
rect 562194 81922 562250 81978
rect 562318 81922 562374 81978
rect 562442 81922 562498 81978
rect 562566 81922 562622 81978
rect 589194 94294 589250 94350
rect 589318 94294 589374 94350
rect 589442 94294 589498 94350
rect 589566 94294 589622 94350
rect 589194 94170 589250 94226
rect 589318 94170 589374 94226
rect 589442 94170 589498 94226
rect 589566 94170 589622 94226
rect 589194 94046 589250 94102
rect 589318 94046 589374 94102
rect 589442 94046 589498 94102
rect 589566 94046 589622 94102
rect 589194 93922 589250 93978
rect 589318 93922 589374 93978
rect 589442 93922 589498 93978
rect 589566 93922 589622 93978
rect 592914 514294 592970 514350
rect 593038 514294 593094 514350
rect 593162 514294 593218 514350
rect 593286 514294 593342 514350
rect 592914 514170 592970 514226
rect 593038 514170 593094 514226
rect 593162 514170 593218 514226
rect 593286 514170 593342 514226
rect 592914 514046 592970 514102
rect 593038 514046 593094 514102
rect 593162 514046 593218 514102
rect 593286 514046 593342 514102
rect 592914 513922 592970 513978
rect 593038 513922 593094 513978
rect 593162 513922 593218 513978
rect 593286 513922 593342 513978
rect 592914 496294 592970 496350
rect 593038 496294 593094 496350
rect 593162 496294 593218 496350
rect 593286 496294 593342 496350
rect 592914 496170 592970 496226
rect 593038 496170 593094 496226
rect 593162 496170 593218 496226
rect 593286 496170 593342 496226
rect 592914 496046 592970 496102
rect 593038 496046 593094 496102
rect 593162 496046 593218 496102
rect 593286 496046 593342 496102
rect 592914 495922 592970 495978
rect 593038 495922 593094 495978
rect 593162 495922 593218 495978
rect 593286 495922 593342 495978
rect 592914 478294 592970 478350
rect 593038 478294 593094 478350
rect 593162 478294 593218 478350
rect 593286 478294 593342 478350
rect 592914 478170 592970 478226
rect 593038 478170 593094 478226
rect 593162 478170 593218 478226
rect 593286 478170 593342 478226
rect 592914 478046 592970 478102
rect 593038 478046 593094 478102
rect 593162 478046 593218 478102
rect 593286 478046 593342 478102
rect 592914 477922 592970 477978
rect 593038 477922 593094 477978
rect 593162 477922 593218 477978
rect 593286 477922 593342 477978
rect 592914 460294 592970 460350
rect 593038 460294 593094 460350
rect 593162 460294 593218 460350
rect 593286 460294 593342 460350
rect 592914 460170 592970 460226
rect 593038 460170 593094 460226
rect 593162 460170 593218 460226
rect 593286 460170 593342 460226
rect 592914 460046 592970 460102
rect 593038 460046 593094 460102
rect 593162 460046 593218 460102
rect 593286 460046 593342 460102
rect 592914 459922 592970 459978
rect 593038 459922 593094 459978
rect 593162 459922 593218 459978
rect 593286 459922 593342 459978
rect 592914 442294 592970 442350
rect 593038 442294 593094 442350
rect 593162 442294 593218 442350
rect 593286 442294 593342 442350
rect 592914 442170 592970 442226
rect 593038 442170 593094 442226
rect 593162 442170 593218 442226
rect 593286 442170 593342 442226
rect 592914 442046 592970 442102
rect 593038 442046 593094 442102
rect 593162 442046 593218 442102
rect 593286 442046 593342 442102
rect 592914 441922 592970 441978
rect 593038 441922 593094 441978
rect 593162 441922 593218 441978
rect 593286 441922 593342 441978
rect 592914 424294 592970 424350
rect 593038 424294 593094 424350
rect 593162 424294 593218 424350
rect 593286 424294 593342 424350
rect 592914 424170 592970 424226
rect 593038 424170 593094 424226
rect 593162 424170 593218 424226
rect 593286 424170 593342 424226
rect 592914 424046 592970 424102
rect 593038 424046 593094 424102
rect 593162 424046 593218 424102
rect 593286 424046 593342 424102
rect 592914 423922 592970 423978
rect 593038 423922 593094 423978
rect 593162 423922 593218 423978
rect 593286 423922 593342 423978
rect 592914 406294 592970 406350
rect 593038 406294 593094 406350
rect 593162 406294 593218 406350
rect 593286 406294 593342 406350
rect 592914 406170 592970 406226
rect 593038 406170 593094 406226
rect 593162 406170 593218 406226
rect 593286 406170 593342 406226
rect 592914 406046 592970 406102
rect 593038 406046 593094 406102
rect 593162 406046 593218 406102
rect 593286 406046 593342 406102
rect 592914 405922 592970 405978
rect 593038 405922 593094 405978
rect 593162 405922 593218 405978
rect 593286 405922 593342 405978
rect 592914 388294 592970 388350
rect 593038 388294 593094 388350
rect 593162 388294 593218 388350
rect 593286 388294 593342 388350
rect 592914 388170 592970 388226
rect 593038 388170 593094 388226
rect 593162 388170 593218 388226
rect 593286 388170 593342 388226
rect 592914 388046 592970 388102
rect 593038 388046 593094 388102
rect 593162 388046 593218 388102
rect 593286 388046 593342 388102
rect 592914 387922 592970 387978
rect 593038 387922 593094 387978
rect 593162 387922 593218 387978
rect 593286 387922 593342 387978
rect 592914 370294 592970 370350
rect 593038 370294 593094 370350
rect 593162 370294 593218 370350
rect 593286 370294 593342 370350
rect 592914 370170 592970 370226
rect 593038 370170 593094 370226
rect 593162 370170 593218 370226
rect 593286 370170 593342 370226
rect 592914 370046 592970 370102
rect 593038 370046 593094 370102
rect 593162 370046 593218 370102
rect 593286 370046 593342 370102
rect 592914 369922 592970 369978
rect 593038 369922 593094 369978
rect 593162 369922 593218 369978
rect 593286 369922 593342 369978
rect 592914 352294 592970 352350
rect 593038 352294 593094 352350
rect 593162 352294 593218 352350
rect 593286 352294 593342 352350
rect 592914 352170 592970 352226
rect 593038 352170 593094 352226
rect 593162 352170 593218 352226
rect 593286 352170 593342 352226
rect 592914 352046 592970 352102
rect 593038 352046 593094 352102
rect 593162 352046 593218 352102
rect 593286 352046 593342 352102
rect 592914 351922 592970 351978
rect 593038 351922 593094 351978
rect 593162 351922 593218 351978
rect 593286 351922 593342 351978
rect 592914 334294 592970 334350
rect 593038 334294 593094 334350
rect 593162 334294 593218 334350
rect 593286 334294 593342 334350
rect 592914 334170 592970 334226
rect 593038 334170 593094 334226
rect 593162 334170 593218 334226
rect 593286 334170 593342 334226
rect 592914 334046 592970 334102
rect 593038 334046 593094 334102
rect 593162 334046 593218 334102
rect 593286 334046 593342 334102
rect 592914 333922 592970 333978
rect 593038 333922 593094 333978
rect 593162 333922 593218 333978
rect 593286 333922 593342 333978
rect 592914 316294 592970 316350
rect 593038 316294 593094 316350
rect 593162 316294 593218 316350
rect 593286 316294 593342 316350
rect 592914 316170 592970 316226
rect 593038 316170 593094 316226
rect 593162 316170 593218 316226
rect 593286 316170 593342 316226
rect 592914 316046 592970 316102
rect 593038 316046 593094 316102
rect 593162 316046 593218 316102
rect 593286 316046 593342 316102
rect 592914 315922 592970 315978
rect 593038 315922 593094 315978
rect 593162 315922 593218 315978
rect 593286 315922 593342 315978
rect 592914 298294 592970 298350
rect 593038 298294 593094 298350
rect 593162 298294 593218 298350
rect 593286 298294 593342 298350
rect 592914 298170 592970 298226
rect 593038 298170 593094 298226
rect 593162 298170 593218 298226
rect 593286 298170 593342 298226
rect 592914 298046 592970 298102
rect 593038 298046 593094 298102
rect 593162 298046 593218 298102
rect 593286 298046 593342 298102
rect 592914 297922 592970 297978
rect 593038 297922 593094 297978
rect 593162 297922 593218 297978
rect 593286 297922 593342 297978
rect 592914 280294 592970 280350
rect 593038 280294 593094 280350
rect 593162 280294 593218 280350
rect 593286 280294 593342 280350
rect 592914 280170 592970 280226
rect 593038 280170 593094 280226
rect 593162 280170 593218 280226
rect 593286 280170 593342 280226
rect 592914 280046 592970 280102
rect 593038 280046 593094 280102
rect 593162 280046 593218 280102
rect 593286 280046 593342 280102
rect 592914 279922 592970 279978
rect 593038 279922 593094 279978
rect 593162 279922 593218 279978
rect 593286 279922 593342 279978
rect 592914 262294 592970 262350
rect 593038 262294 593094 262350
rect 593162 262294 593218 262350
rect 593286 262294 593342 262350
rect 592914 262170 592970 262226
rect 593038 262170 593094 262226
rect 593162 262170 593218 262226
rect 593286 262170 593342 262226
rect 592914 262046 592970 262102
rect 593038 262046 593094 262102
rect 593162 262046 593218 262102
rect 593286 262046 593342 262102
rect 592914 261922 592970 261978
rect 593038 261922 593094 261978
rect 593162 261922 593218 261978
rect 593286 261922 593342 261978
rect 592914 244294 592970 244350
rect 593038 244294 593094 244350
rect 593162 244294 593218 244350
rect 593286 244294 593342 244350
rect 592914 244170 592970 244226
rect 593038 244170 593094 244226
rect 593162 244170 593218 244226
rect 593286 244170 593342 244226
rect 592914 244046 592970 244102
rect 593038 244046 593094 244102
rect 593162 244046 593218 244102
rect 593286 244046 593342 244102
rect 592914 243922 592970 243978
rect 593038 243922 593094 243978
rect 593162 243922 593218 243978
rect 593286 243922 593342 243978
rect 590492 78002 590548 78058
rect 592914 226294 592970 226350
rect 593038 226294 593094 226350
rect 593162 226294 593218 226350
rect 593286 226294 593342 226350
rect 592914 226170 592970 226226
rect 593038 226170 593094 226226
rect 593162 226170 593218 226226
rect 593286 226170 593342 226226
rect 592914 226046 592970 226102
rect 593038 226046 593094 226102
rect 593162 226046 593218 226102
rect 593286 226046 593342 226102
rect 592914 225922 592970 225978
rect 593038 225922 593094 225978
rect 593162 225922 593218 225978
rect 593286 225922 593342 225978
rect 592914 208294 592970 208350
rect 593038 208294 593094 208350
rect 593162 208294 593218 208350
rect 593286 208294 593342 208350
rect 592914 208170 592970 208226
rect 593038 208170 593094 208226
rect 593162 208170 593218 208226
rect 593286 208170 593342 208226
rect 592914 208046 592970 208102
rect 593038 208046 593094 208102
rect 593162 208046 593218 208102
rect 593286 208046 593342 208102
rect 592914 207922 592970 207978
rect 593038 207922 593094 207978
rect 593162 207922 593218 207978
rect 593286 207922 593342 207978
rect 592914 190294 592970 190350
rect 593038 190294 593094 190350
rect 593162 190294 593218 190350
rect 593286 190294 593342 190350
rect 592914 190170 592970 190226
rect 593038 190170 593094 190226
rect 593162 190170 593218 190226
rect 593286 190170 593342 190226
rect 592914 190046 592970 190102
rect 593038 190046 593094 190102
rect 593162 190046 593218 190102
rect 593286 190046 593342 190102
rect 592914 189922 592970 189978
rect 593038 189922 593094 189978
rect 593162 189922 593218 189978
rect 593286 189922 593342 189978
rect 592914 172294 592970 172350
rect 593038 172294 593094 172350
rect 593162 172294 593218 172350
rect 593286 172294 593342 172350
rect 592914 172170 592970 172226
rect 593038 172170 593094 172226
rect 593162 172170 593218 172226
rect 593286 172170 593342 172226
rect 592914 172046 592970 172102
rect 593038 172046 593094 172102
rect 593162 172046 593218 172102
rect 593286 172046 593342 172102
rect 592914 171922 592970 171978
rect 593038 171922 593094 171978
rect 593162 171922 593218 171978
rect 593286 171922 593342 171978
rect 592914 154294 592970 154350
rect 593038 154294 593094 154350
rect 593162 154294 593218 154350
rect 593286 154294 593342 154350
rect 592914 154170 592970 154226
rect 593038 154170 593094 154226
rect 593162 154170 593218 154226
rect 593286 154170 593342 154226
rect 592914 154046 592970 154102
rect 593038 154046 593094 154102
rect 593162 154046 593218 154102
rect 593286 154046 593342 154102
rect 592914 153922 592970 153978
rect 593038 153922 593094 153978
rect 593162 153922 593218 153978
rect 593286 153922 593342 153978
rect 592914 136294 592970 136350
rect 593038 136294 593094 136350
rect 593162 136294 593218 136350
rect 593286 136294 593342 136350
rect 592914 136170 592970 136226
rect 593038 136170 593094 136226
rect 593162 136170 593218 136226
rect 593286 136170 593342 136226
rect 592914 136046 592970 136102
rect 593038 136046 593094 136102
rect 593162 136046 593218 136102
rect 593286 136046 593342 136102
rect 592914 135922 592970 135978
rect 593038 135922 593094 135978
rect 593162 135922 593218 135978
rect 593286 135922 593342 135978
rect 592914 118294 592970 118350
rect 593038 118294 593094 118350
rect 593162 118294 593218 118350
rect 593286 118294 593342 118350
rect 592914 118170 592970 118226
rect 593038 118170 593094 118226
rect 593162 118170 593218 118226
rect 593286 118170 593342 118226
rect 592914 118046 592970 118102
rect 593038 118046 593094 118102
rect 593162 118046 593218 118102
rect 593286 118046 593342 118102
rect 592914 117922 592970 117978
rect 593038 117922 593094 117978
rect 593162 117922 593218 117978
rect 593286 117922 593342 117978
rect 592914 100294 592970 100350
rect 593038 100294 593094 100350
rect 593162 100294 593218 100350
rect 593286 100294 593342 100350
rect 592914 100170 592970 100226
rect 593038 100170 593094 100226
rect 593162 100170 593218 100226
rect 593286 100170 593342 100226
rect 592914 100046 592970 100102
rect 593038 100046 593094 100102
rect 593162 100046 593218 100102
rect 593286 100046 593342 100102
rect 592914 99922 592970 99978
rect 593038 99922 593094 99978
rect 593162 99922 593218 99978
rect 593286 99922 593342 99978
rect 592914 82294 592970 82350
rect 593038 82294 593094 82350
rect 593162 82294 593218 82350
rect 593286 82294 593342 82350
rect 592914 82170 592970 82226
rect 593038 82170 593094 82226
rect 593162 82170 593218 82226
rect 593286 82170 593342 82226
rect 592914 82046 592970 82102
rect 593038 82046 593094 82102
rect 593162 82046 593218 82102
rect 593286 82046 593342 82102
rect 592914 81922 592970 81978
rect 593038 81922 593094 81978
rect 593162 81922 593218 81978
rect 593286 81922 593342 81978
rect 589194 76294 589250 76350
rect 589318 76294 589374 76350
rect 589442 76294 589498 76350
rect 589566 76294 589622 76350
rect 589194 76170 589250 76226
rect 589318 76170 589374 76226
rect 589442 76170 589498 76226
rect 589566 76170 589622 76226
rect 589194 76046 589250 76102
rect 589318 76046 589374 76102
rect 589442 76046 589498 76102
rect 589566 76046 589622 76102
rect 589194 75922 589250 75978
rect 589318 75922 589374 75978
rect 589442 75922 589498 75978
rect 589566 75922 589622 75978
rect 562194 64294 562250 64350
rect 562318 64294 562374 64350
rect 562442 64294 562498 64350
rect 562566 64294 562622 64350
rect 562194 64170 562250 64226
rect 562318 64170 562374 64226
rect 562442 64170 562498 64226
rect 562566 64170 562622 64226
rect 562194 64046 562250 64102
rect 562318 64046 562374 64102
rect 562442 64046 562498 64102
rect 562566 64046 562622 64102
rect 562194 63922 562250 63978
rect 562318 63922 562374 63978
rect 562442 63922 562498 63978
rect 562566 63922 562622 63978
rect 558474 40294 558530 40350
rect 558598 40294 558654 40350
rect 558722 40294 558778 40350
rect 558846 40294 558902 40350
rect 558474 40170 558530 40226
rect 558598 40170 558654 40226
rect 558722 40170 558778 40226
rect 558846 40170 558902 40226
rect 558474 40046 558530 40102
rect 558598 40046 558654 40102
rect 558722 40046 558778 40102
rect 558846 40046 558902 40102
rect 558474 39922 558530 39978
rect 558598 39922 558654 39978
rect 558722 39922 558778 39978
rect 558846 39922 558902 39978
rect 558474 22294 558530 22350
rect 558598 22294 558654 22350
rect 558722 22294 558778 22350
rect 558846 22294 558902 22350
rect 558474 22170 558530 22226
rect 558598 22170 558654 22226
rect 558722 22170 558778 22226
rect 558846 22170 558902 22226
rect 558474 22046 558530 22102
rect 558598 22046 558654 22102
rect 558722 22046 558778 22102
rect 558846 22046 558902 22102
rect 558474 21922 558530 21978
rect 558598 21922 558654 21978
rect 558722 21922 558778 21978
rect 558846 21922 558902 21978
rect 558474 4294 558530 4350
rect 558598 4294 558654 4350
rect 558722 4294 558778 4350
rect 558846 4294 558902 4350
rect 558474 4170 558530 4226
rect 558598 4170 558654 4226
rect 558722 4170 558778 4226
rect 558846 4170 558902 4226
rect 561148 55502 561204 55558
rect 572908 67202 572964 67258
rect 562194 46294 562250 46350
rect 562318 46294 562374 46350
rect 562442 46294 562498 46350
rect 562566 46294 562622 46350
rect 562194 46170 562250 46226
rect 562318 46170 562374 46226
rect 562442 46170 562498 46226
rect 562566 46170 562622 46226
rect 562194 46046 562250 46102
rect 562318 46046 562374 46102
rect 562442 46046 562498 46102
rect 562566 46046 562622 46102
rect 562194 45922 562250 45978
rect 562318 45922 562374 45978
rect 562442 45922 562498 45978
rect 562566 45922 562622 45978
rect 566188 53882 566244 53938
rect 562194 28294 562250 28350
rect 562318 28294 562374 28350
rect 562442 28294 562498 28350
rect 562566 28294 562622 28350
rect 562194 28170 562250 28226
rect 562318 28170 562374 28226
rect 562442 28170 562498 28226
rect 562566 28170 562622 28226
rect 562194 28046 562250 28102
rect 562318 28046 562374 28102
rect 562442 28046 562498 28102
rect 562566 28046 562622 28102
rect 562194 27922 562250 27978
rect 562318 27922 562374 27978
rect 562442 27922 562498 27978
rect 562566 27922 562622 27978
rect 562194 10294 562250 10350
rect 562318 10294 562374 10350
rect 562442 10294 562498 10350
rect 562566 10294 562622 10350
rect 562194 10170 562250 10226
rect 562318 10170 562374 10226
rect 562442 10170 562498 10226
rect 562566 10170 562622 10226
rect 562194 10046 562250 10102
rect 562318 10046 562374 10102
rect 562442 10046 562498 10102
rect 562566 10046 562622 10102
rect 562194 9922 562250 9978
rect 562318 9922 562374 9978
rect 562442 9922 562498 9978
rect 562566 9922 562622 9978
rect 558474 4046 558530 4102
rect 558598 4046 558654 4102
rect 558722 4046 558778 4102
rect 558846 4046 558902 4102
rect 558474 3922 558530 3978
rect 558598 3922 558654 3978
rect 558722 3922 558778 3978
rect 558846 3922 558902 3978
rect 557788 3122 557844 3178
rect 542556 1322 542612 1378
rect 531474 -1176 531530 -1120
rect 531598 -1176 531654 -1120
rect 531722 -1176 531778 -1120
rect 531846 -1176 531902 -1120
rect 531474 -1300 531530 -1244
rect 531598 -1300 531654 -1244
rect 531722 -1300 531778 -1244
rect 531846 -1300 531902 -1244
rect 531474 -1424 531530 -1368
rect 531598 -1424 531654 -1368
rect 531722 -1424 531778 -1368
rect 531846 -1424 531902 -1368
rect 531474 -1548 531530 -1492
rect 531598 -1548 531654 -1492
rect 531722 -1548 531778 -1492
rect 531846 -1548 531902 -1492
rect 558474 -216 558530 -160
rect 558598 -216 558654 -160
rect 558722 -216 558778 -160
rect 558846 -216 558902 -160
rect 558474 -340 558530 -284
rect 558598 -340 558654 -284
rect 558722 -340 558778 -284
rect 558846 -340 558902 -284
rect 558474 -464 558530 -408
rect 558598 -464 558654 -408
rect 558722 -464 558778 -408
rect 558846 -464 558902 -408
rect 558474 -588 558530 -532
rect 558598 -588 558654 -532
rect 558722 -588 558778 -532
rect 558846 -588 558902 -532
rect 564508 31922 564564 31978
rect 563500 6722 563556 6778
rect 576268 65582 576324 65638
rect 574588 25262 574644 25318
rect 589194 58294 589250 58350
rect 589318 58294 589374 58350
rect 589442 58294 589498 58350
rect 589566 58294 589622 58350
rect 589194 58170 589250 58226
rect 589318 58170 589374 58226
rect 589442 58170 589498 58226
rect 589566 58170 589622 58226
rect 589194 58046 589250 58102
rect 589318 58046 589374 58102
rect 589442 58046 589498 58102
rect 589566 58046 589622 58102
rect 589194 57922 589250 57978
rect 589318 57922 589374 57978
rect 589442 57922 589498 57978
rect 589566 57922 589622 57978
rect 592914 64294 592970 64350
rect 593038 64294 593094 64350
rect 593162 64294 593218 64350
rect 593286 64294 593342 64350
rect 592914 64170 592970 64226
rect 593038 64170 593094 64226
rect 593162 64170 593218 64226
rect 593286 64170 593342 64226
rect 592914 64046 592970 64102
rect 593038 64046 593094 64102
rect 593162 64046 593218 64102
rect 593286 64046 593342 64102
rect 592914 63922 592970 63978
rect 593038 63922 593094 63978
rect 593162 63922 593218 63978
rect 593286 63922 593342 63978
rect 589194 40294 589250 40350
rect 589318 40294 589374 40350
rect 589442 40294 589498 40350
rect 589566 40294 589622 40350
rect 589194 40170 589250 40226
rect 589318 40170 589374 40226
rect 589442 40170 589498 40226
rect 589566 40170 589622 40226
rect 589194 40046 589250 40102
rect 589318 40046 589374 40102
rect 589442 40046 589498 40102
rect 589566 40046 589622 40102
rect 589194 39922 589250 39978
rect 589318 39922 589374 39978
rect 589442 39922 589498 39978
rect 589566 39922 589622 39978
rect 592914 46294 592970 46350
rect 593038 46294 593094 46350
rect 593162 46294 593218 46350
rect 593286 46294 593342 46350
rect 592914 46170 592970 46226
rect 593038 46170 593094 46226
rect 593162 46170 593218 46226
rect 593286 46170 593342 46226
rect 592914 46046 592970 46102
rect 593038 46046 593094 46102
rect 593162 46046 593218 46102
rect 593286 46046 593342 46102
rect 592914 45922 592970 45978
rect 593038 45922 593094 45978
rect 593162 45922 593218 45978
rect 593286 45922 593342 45978
rect 589194 22294 589250 22350
rect 589318 22294 589374 22350
rect 589442 22294 589498 22350
rect 589566 22294 589622 22350
rect 589194 22170 589250 22226
rect 589318 22170 589374 22226
rect 589442 22170 589498 22226
rect 589566 22170 589622 22226
rect 589194 22046 589250 22102
rect 589318 22046 589374 22102
rect 589442 22046 589498 22102
rect 589566 22046 589622 22102
rect 589194 21922 589250 21978
rect 589318 21922 589374 21978
rect 589442 21922 589498 21978
rect 589566 21922 589622 21978
rect 589194 4294 589250 4350
rect 589318 4294 589374 4350
rect 589442 4294 589498 4350
rect 589566 4294 589622 4350
rect 589194 4170 589250 4226
rect 589318 4170 589374 4226
rect 589442 4170 589498 4226
rect 589566 4170 589622 4226
rect 589194 4046 589250 4102
rect 589318 4046 589374 4102
rect 589442 4046 589498 4102
rect 589566 4046 589622 4102
rect 589194 3922 589250 3978
rect 589318 3922 589374 3978
rect 589442 3922 589498 3978
rect 589566 3922 589622 3978
rect 569548 1502 569604 1558
rect 562194 -1176 562250 -1120
rect 562318 -1176 562374 -1120
rect 562442 -1176 562498 -1120
rect 562566 -1176 562622 -1120
rect 562194 -1300 562250 -1244
rect 562318 -1300 562374 -1244
rect 562442 -1300 562498 -1244
rect 562566 -1300 562622 -1244
rect 562194 -1424 562250 -1368
rect 562318 -1424 562374 -1368
rect 562442 -1424 562498 -1368
rect 562566 -1424 562622 -1368
rect 562194 -1548 562250 -1492
rect 562318 -1548 562374 -1492
rect 562442 -1548 562498 -1492
rect 562566 -1548 562622 -1492
rect 589194 -216 589250 -160
rect 589318 -216 589374 -160
rect 589442 -216 589498 -160
rect 589566 -216 589622 -160
rect 589194 -340 589250 -284
rect 589318 -340 589374 -284
rect 589442 -340 589498 -284
rect 589566 -340 589622 -284
rect 589194 -464 589250 -408
rect 589318 -464 589374 -408
rect 589442 -464 589498 -408
rect 589566 -464 589622 -408
rect 589194 -588 589250 -532
rect 589318 -588 589374 -532
rect 589442 -588 589498 -532
rect 589566 -588 589622 -532
rect 592914 28294 592970 28350
rect 593038 28294 593094 28350
rect 593162 28294 593218 28350
rect 593286 28294 593342 28350
rect 592914 28170 592970 28226
rect 593038 28170 593094 28226
rect 593162 28170 593218 28226
rect 593286 28170 593342 28226
rect 592914 28046 592970 28102
rect 593038 28046 593094 28102
rect 593162 28046 593218 28102
rect 593286 28046 593342 28102
rect 592914 27922 592970 27978
rect 593038 27922 593094 27978
rect 593162 27922 593218 27978
rect 593286 27922 593342 27978
rect 592914 10294 592970 10350
rect 593038 10294 593094 10350
rect 593162 10294 593218 10350
rect 593286 10294 593342 10350
rect 592914 10170 592970 10226
rect 593038 10170 593094 10226
rect 593162 10170 593218 10226
rect 593286 10170 593342 10226
rect 592914 10046 592970 10102
rect 593038 10046 593094 10102
rect 593162 10046 593218 10102
rect 593286 10046 593342 10102
rect 592914 9922 592970 9978
rect 593038 9922 593094 9978
rect 593162 9922 593218 9978
rect 593286 9922 593342 9978
rect 596496 597156 596552 597212
rect 596620 597156 596676 597212
rect 596744 597156 596800 597212
rect 596868 597156 596924 597212
rect 596496 597032 596552 597088
rect 596620 597032 596676 597088
rect 596744 597032 596800 597088
rect 596868 597032 596924 597088
rect 596496 596908 596552 596964
rect 596620 596908 596676 596964
rect 596744 596908 596800 596964
rect 596868 596908 596924 596964
rect 596496 596784 596552 596840
rect 596620 596784 596676 596840
rect 596744 596784 596800 596840
rect 596868 596784 596924 596840
rect 596496 580294 596552 580350
rect 596620 580294 596676 580350
rect 596744 580294 596800 580350
rect 596868 580294 596924 580350
rect 596496 580170 596552 580226
rect 596620 580170 596676 580226
rect 596744 580170 596800 580226
rect 596868 580170 596924 580226
rect 596496 580046 596552 580102
rect 596620 580046 596676 580102
rect 596744 580046 596800 580102
rect 596868 580046 596924 580102
rect 596496 579922 596552 579978
rect 596620 579922 596676 579978
rect 596744 579922 596800 579978
rect 596868 579922 596924 579978
rect 596496 562294 596552 562350
rect 596620 562294 596676 562350
rect 596744 562294 596800 562350
rect 596868 562294 596924 562350
rect 596496 562170 596552 562226
rect 596620 562170 596676 562226
rect 596744 562170 596800 562226
rect 596868 562170 596924 562226
rect 596496 562046 596552 562102
rect 596620 562046 596676 562102
rect 596744 562046 596800 562102
rect 596868 562046 596924 562102
rect 596496 561922 596552 561978
rect 596620 561922 596676 561978
rect 596744 561922 596800 561978
rect 596868 561922 596924 561978
rect 596496 544294 596552 544350
rect 596620 544294 596676 544350
rect 596744 544294 596800 544350
rect 596868 544294 596924 544350
rect 596496 544170 596552 544226
rect 596620 544170 596676 544226
rect 596744 544170 596800 544226
rect 596868 544170 596924 544226
rect 596496 544046 596552 544102
rect 596620 544046 596676 544102
rect 596744 544046 596800 544102
rect 596868 544046 596924 544102
rect 596496 543922 596552 543978
rect 596620 543922 596676 543978
rect 596744 543922 596800 543978
rect 596868 543922 596924 543978
rect 596496 526294 596552 526350
rect 596620 526294 596676 526350
rect 596744 526294 596800 526350
rect 596868 526294 596924 526350
rect 596496 526170 596552 526226
rect 596620 526170 596676 526226
rect 596744 526170 596800 526226
rect 596868 526170 596924 526226
rect 596496 526046 596552 526102
rect 596620 526046 596676 526102
rect 596744 526046 596800 526102
rect 596868 526046 596924 526102
rect 596496 525922 596552 525978
rect 596620 525922 596676 525978
rect 596744 525922 596800 525978
rect 596868 525922 596924 525978
rect 596496 508294 596552 508350
rect 596620 508294 596676 508350
rect 596744 508294 596800 508350
rect 596868 508294 596924 508350
rect 596496 508170 596552 508226
rect 596620 508170 596676 508226
rect 596744 508170 596800 508226
rect 596868 508170 596924 508226
rect 596496 508046 596552 508102
rect 596620 508046 596676 508102
rect 596744 508046 596800 508102
rect 596868 508046 596924 508102
rect 596496 507922 596552 507978
rect 596620 507922 596676 507978
rect 596744 507922 596800 507978
rect 596868 507922 596924 507978
rect 596496 490294 596552 490350
rect 596620 490294 596676 490350
rect 596744 490294 596800 490350
rect 596868 490294 596924 490350
rect 596496 490170 596552 490226
rect 596620 490170 596676 490226
rect 596744 490170 596800 490226
rect 596868 490170 596924 490226
rect 596496 490046 596552 490102
rect 596620 490046 596676 490102
rect 596744 490046 596800 490102
rect 596868 490046 596924 490102
rect 596496 489922 596552 489978
rect 596620 489922 596676 489978
rect 596744 489922 596800 489978
rect 596868 489922 596924 489978
rect 596496 472294 596552 472350
rect 596620 472294 596676 472350
rect 596744 472294 596800 472350
rect 596868 472294 596924 472350
rect 596496 472170 596552 472226
rect 596620 472170 596676 472226
rect 596744 472170 596800 472226
rect 596868 472170 596924 472226
rect 596496 472046 596552 472102
rect 596620 472046 596676 472102
rect 596744 472046 596800 472102
rect 596868 472046 596924 472102
rect 596496 471922 596552 471978
rect 596620 471922 596676 471978
rect 596744 471922 596800 471978
rect 596868 471922 596924 471978
rect 596496 454294 596552 454350
rect 596620 454294 596676 454350
rect 596744 454294 596800 454350
rect 596868 454294 596924 454350
rect 596496 454170 596552 454226
rect 596620 454170 596676 454226
rect 596744 454170 596800 454226
rect 596868 454170 596924 454226
rect 596496 454046 596552 454102
rect 596620 454046 596676 454102
rect 596744 454046 596800 454102
rect 596868 454046 596924 454102
rect 596496 453922 596552 453978
rect 596620 453922 596676 453978
rect 596744 453922 596800 453978
rect 596868 453922 596924 453978
rect 596496 436294 596552 436350
rect 596620 436294 596676 436350
rect 596744 436294 596800 436350
rect 596868 436294 596924 436350
rect 596496 436170 596552 436226
rect 596620 436170 596676 436226
rect 596744 436170 596800 436226
rect 596868 436170 596924 436226
rect 596496 436046 596552 436102
rect 596620 436046 596676 436102
rect 596744 436046 596800 436102
rect 596868 436046 596924 436102
rect 596496 435922 596552 435978
rect 596620 435922 596676 435978
rect 596744 435922 596800 435978
rect 596868 435922 596924 435978
rect 596496 418294 596552 418350
rect 596620 418294 596676 418350
rect 596744 418294 596800 418350
rect 596868 418294 596924 418350
rect 596496 418170 596552 418226
rect 596620 418170 596676 418226
rect 596744 418170 596800 418226
rect 596868 418170 596924 418226
rect 596496 418046 596552 418102
rect 596620 418046 596676 418102
rect 596744 418046 596800 418102
rect 596868 418046 596924 418102
rect 596496 417922 596552 417978
rect 596620 417922 596676 417978
rect 596744 417922 596800 417978
rect 596868 417922 596924 417978
rect 596496 400294 596552 400350
rect 596620 400294 596676 400350
rect 596744 400294 596800 400350
rect 596868 400294 596924 400350
rect 596496 400170 596552 400226
rect 596620 400170 596676 400226
rect 596744 400170 596800 400226
rect 596868 400170 596924 400226
rect 596496 400046 596552 400102
rect 596620 400046 596676 400102
rect 596744 400046 596800 400102
rect 596868 400046 596924 400102
rect 596496 399922 596552 399978
rect 596620 399922 596676 399978
rect 596744 399922 596800 399978
rect 596868 399922 596924 399978
rect 596496 382294 596552 382350
rect 596620 382294 596676 382350
rect 596744 382294 596800 382350
rect 596868 382294 596924 382350
rect 596496 382170 596552 382226
rect 596620 382170 596676 382226
rect 596744 382170 596800 382226
rect 596868 382170 596924 382226
rect 596496 382046 596552 382102
rect 596620 382046 596676 382102
rect 596744 382046 596800 382102
rect 596868 382046 596924 382102
rect 596496 381922 596552 381978
rect 596620 381922 596676 381978
rect 596744 381922 596800 381978
rect 596868 381922 596924 381978
rect 596496 364294 596552 364350
rect 596620 364294 596676 364350
rect 596744 364294 596800 364350
rect 596868 364294 596924 364350
rect 596496 364170 596552 364226
rect 596620 364170 596676 364226
rect 596744 364170 596800 364226
rect 596868 364170 596924 364226
rect 596496 364046 596552 364102
rect 596620 364046 596676 364102
rect 596744 364046 596800 364102
rect 596868 364046 596924 364102
rect 596496 363922 596552 363978
rect 596620 363922 596676 363978
rect 596744 363922 596800 363978
rect 596868 363922 596924 363978
rect 596496 346294 596552 346350
rect 596620 346294 596676 346350
rect 596744 346294 596800 346350
rect 596868 346294 596924 346350
rect 596496 346170 596552 346226
rect 596620 346170 596676 346226
rect 596744 346170 596800 346226
rect 596868 346170 596924 346226
rect 596496 346046 596552 346102
rect 596620 346046 596676 346102
rect 596744 346046 596800 346102
rect 596868 346046 596924 346102
rect 596496 345922 596552 345978
rect 596620 345922 596676 345978
rect 596744 345922 596800 345978
rect 596868 345922 596924 345978
rect 596496 328294 596552 328350
rect 596620 328294 596676 328350
rect 596744 328294 596800 328350
rect 596868 328294 596924 328350
rect 596496 328170 596552 328226
rect 596620 328170 596676 328226
rect 596744 328170 596800 328226
rect 596868 328170 596924 328226
rect 596496 328046 596552 328102
rect 596620 328046 596676 328102
rect 596744 328046 596800 328102
rect 596868 328046 596924 328102
rect 596496 327922 596552 327978
rect 596620 327922 596676 327978
rect 596744 327922 596800 327978
rect 596868 327922 596924 327978
rect 596496 310294 596552 310350
rect 596620 310294 596676 310350
rect 596744 310294 596800 310350
rect 596868 310294 596924 310350
rect 596496 310170 596552 310226
rect 596620 310170 596676 310226
rect 596744 310170 596800 310226
rect 596868 310170 596924 310226
rect 596496 310046 596552 310102
rect 596620 310046 596676 310102
rect 596744 310046 596800 310102
rect 596868 310046 596924 310102
rect 596496 309922 596552 309978
rect 596620 309922 596676 309978
rect 596744 309922 596800 309978
rect 596868 309922 596924 309978
rect 596496 292294 596552 292350
rect 596620 292294 596676 292350
rect 596744 292294 596800 292350
rect 596868 292294 596924 292350
rect 596496 292170 596552 292226
rect 596620 292170 596676 292226
rect 596744 292170 596800 292226
rect 596868 292170 596924 292226
rect 596496 292046 596552 292102
rect 596620 292046 596676 292102
rect 596744 292046 596800 292102
rect 596868 292046 596924 292102
rect 596496 291922 596552 291978
rect 596620 291922 596676 291978
rect 596744 291922 596800 291978
rect 596868 291922 596924 291978
rect 596496 274294 596552 274350
rect 596620 274294 596676 274350
rect 596744 274294 596800 274350
rect 596868 274294 596924 274350
rect 596496 274170 596552 274226
rect 596620 274170 596676 274226
rect 596744 274170 596800 274226
rect 596868 274170 596924 274226
rect 596496 274046 596552 274102
rect 596620 274046 596676 274102
rect 596744 274046 596800 274102
rect 596868 274046 596924 274102
rect 596496 273922 596552 273978
rect 596620 273922 596676 273978
rect 596744 273922 596800 273978
rect 596868 273922 596924 273978
rect 596496 256294 596552 256350
rect 596620 256294 596676 256350
rect 596744 256294 596800 256350
rect 596868 256294 596924 256350
rect 596496 256170 596552 256226
rect 596620 256170 596676 256226
rect 596744 256170 596800 256226
rect 596868 256170 596924 256226
rect 596496 256046 596552 256102
rect 596620 256046 596676 256102
rect 596744 256046 596800 256102
rect 596868 256046 596924 256102
rect 596496 255922 596552 255978
rect 596620 255922 596676 255978
rect 596744 255922 596800 255978
rect 596868 255922 596924 255978
rect 596496 238294 596552 238350
rect 596620 238294 596676 238350
rect 596744 238294 596800 238350
rect 596868 238294 596924 238350
rect 596496 238170 596552 238226
rect 596620 238170 596676 238226
rect 596744 238170 596800 238226
rect 596868 238170 596924 238226
rect 596496 238046 596552 238102
rect 596620 238046 596676 238102
rect 596744 238046 596800 238102
rect 596868 238046 596924 238102
rect 596496 237922 596552 237978
rect 596620 237922 596676 237978
rect 596744 237922 596800 237978
rect 596868 237922 596924 237978
rect 596496 220294 596552 220350
rect 596620 220294 596676 220350
rect 596744 220294 596800 220350
rect 596868 220294 596924 220350
rect 596496 220170 596552 220226
rect 596620 220170 596676 220226
rect 596744 220170 596800 220226
rect 596868 220170 596924 220226
rect 596496 220046 596552 220102
rect 596620 220046 596676 220102
rect 596744 220046 596800 220102
rect 596868 220046 596924 220102
rect 596496 219922 596552 219978
rect 596620 219922 596676 219978
rect 596744 219922 596800 219978
rect 596868 219922 596924 219978
rect 596496 202294 596552 202350
rect 596620 202294 596676 202350
rect 596744 202294 596800 202350
rect 596868 202294 596924 202350
rect 596496 202170 596552 202226
rect 596620 202170 596676 202226
rect 596744 202170 596800 202226
rect 596868 202170 596924 202226
rect 596496 202046 596552 202102
rect 596620 202046 596676 202102
rect 596744 202046 596800 202102
rect 596868 202046 596924 202102
rect 596496 201922 596552 201978
rect 596620 201922 596676 201978
rect 596744 201922 596800 201978
rect 596868 201922 596924 201978
rect 596496 184294 596552 184350
rect 596620 184294 596676 184350
rect 596744 184294 596800 184350
rect 596868 184294 596924 184350
rect 596496 184170 596552 184226
rect 596620 184170 596676 184226
rect 596744 184170 596800 184226
rect 596868 184170 596924 184226
rect 596496 184046 596552 184102
rect 596620 184046 596676 184102
rect 596744 184046 596800 184102
rect 596868 184046 596924 184102
rect 596496 183922 596552 183978
rect 596620 183922 596676 183978
rect 596744 183922 596800 183978
rect 596868 183922 596924 183978
rect 596496 166294 596552 166350
rect 596620 166294 596676 166350
rect 596744 166294 596800 166350
rect 596868 166294 596924 166350
rect 596496 166170 596552 166226
rect 596620 166170 596676 166226
rect 596744 166170 596800 166226
rect 596868 166170 596924 166226
rect 596496 166046 596552 166102
rect 596620 166046 596676 166102
rect 596744 166046 596800 166102
rect 596868 166046 596924 166102
rect 596496 165922 596552 165978
rect 596620 165922 596676 165978
rect 596744 165922 596800 165978
rect 596868 165922 596924 165978
rect 596496 148294 596552 148350
rect 596620 148294 596676 148350
rect 596744 148294 596800 148350
rect 596868 148294 596924 148350
rect 596496 148170 596552 148226
rect 596620 148170 596676 148226
rect 596744 148170 596800 148226
rect 596868 148170 596924 148226
rect 596496 148046 596552 148102
rect 596620 148046 596676 148102
rect 596744 148046 596800 148102
rect 596868 148046 596924 148102
rect 596496 147922 596552 147978
rect 596620 147922 596676 147978
rect 596744 147922 596800 147978
rect 596868 147922 596924 147978
rect 596496 130294 596552 130350
rect 596620 130294 596676 130350
rect 596744 130294 596800 130350
rect 596868 130294 596924 130350
rect 596496 130170 596552 130226
rect 596620 130170 596676 130226
rect 596744 130170 596800 130226
rect 596868 130170 596924 130226
rect 596496 130046 596552 130102
rect 596620 130046 596676 130102
rect 596744 130046 596800 130102
rect 596868 130046 596924 130102
rect 596496 129922 596552 129978
rect 596620 129922 596676 129978
rect 596744 129922 596800 129978
rect 596868 129922 596924 129978
rect 596496 112294 596552 112350
rect 596620 112294 596676 112350
rect 596744 112294 596800 112350
rect 596868 112294 596924 112350
rect 596496 112170 596552 112226
rect 596620 112170 596676 112226
rect 596744 112170 596800 112226
rect 596868 112170 596924 112226
rect 596496 112046 596552 112102
rect 596620 112046 596676 112102
rect 596744 112046 596800 112102
rect 596868 112046 596924 112102
rect 596496 111922 596552 111978
rect 596620 111922 596676 111978
rect 596744 111922 596800 111978
rect 596868 111922 596924 111978
rect 596496 94294 596552 94350
rect 596620 94294 596676 94350
rect 596744 94294 596800 94350
rect 596868 94294 596924 94350
rect 596496 94170 596552 94226
rect 596620 94170 596676 94226
rect 596744 94170 596800 94226
rect 596868 94170 596924 94226
rect 596496 94046 596552 94102
rect 596620 94046 596676 94102
rect 596744 94046 596800 94102
rect 596868 94046 596924 94102
rect 596496 93922 596552 93978
rect 596620 93922 596676 93978
rect 596744 93922 596800 93978
rect 596868 93922 596924 93978
rect 596496 76294 596552 76350
rect 596620 76294 596676 76350
rect 596744 76294 596800 76350
rect 596868 76294 596924 76350
rect 596496 76170 596552 76226
rect 596620 76170 596676 76226
rect 596744 76170 596800 76226
rect 596868 76170 596924 76226
rect 596496 76046 596552 76102
rect 596620 76046 596676 76102
rect 596744 76046 596800 76102
rect 596868 76046 596924 76102
rect 596496 75922 596552 75978
rect 596620 75922 596676 75978
rect 596744 75922 596800 75978
rect 596868 75922 596924 75978
rect 596496 58294 596552 58350
rect 596620 58294 596676 58350
rect 596744 58294 596800 58350
rect 596868 58294 596924 58350
rect 596496 58170 596552 58226
rect 596620 58170 596676 58226
rect 596744 58170 596800 58226
rect 596868 58170 596924 58226
rect 596496 58046 596552 58102
rect 596620 58046 596676 58102
rect 596744 58046 596800 58102
rect 596868 58046 596924 58102
rect 596496 57922 596552 57978
rect 596620 57922 596676 57978
rect 596744 57922 596800 57978
rect 596868 57922 596924 57978
rect 596496 40294 596552 40350
rect 596620 40294 596676 40350
rect 596744 40294 596800 40350
rect 596868 40294 596924 40350
rect 596496 40170 596552 40226
rect 596620 40170 596676 40226
rect 596744 40170 596800 40226
rect 596868 40170 596924 40226
rect 596496 40046 596552 40102
rect 596620 40046 596676 40102
rect 596744 40046 596800 40102
rect 596868 40046 596924 40102
rect 596496 39922 596552 39978
rect 596620 39922 596676 39978
rect 596744 39922 596800 39978
rect 596868 39922 596924 39978
rect 596496 22294 596552 22350
rect 596620 22294 596676 22350
rect 596744 22294 596800 22350
rect 596868 22294 596924 22350
rect 596496 22170 596552 22226
rect 596620 22170 596676 22226
rect 596744 22170 596800 22226
rect 596868 22170 596924 22226
rect 596496 22046 596552 22102
rect 596620 22046 596676 22102
rect 596744 22046 596800 22102
rect 596868 22046 596924 22102
rect 596496 21922 596552 21978
rect 596620 21922 596676 21978
rect 596744 21922 596800 21978
rect 596868 21922 596924 21978
rect 596496 4294 596552 4350
rect 596620 4294 596676 4350
rect 596744 4294 596800 4350
rect 596868 4294 596924 4350
rect 596496 4170 596552 4226
rect 596620 4170 596676 4226
rect 596744 4170 596800 4226
rect 596868 4170 596924 4226
rect 596496 4046 596552 4102
rect 596620 4046 596676 4102
rect 596744 4046 596800 4102
rect 596868 4046 596924 4102
rect 596496 3922 596552 3978
rect 596620 3922 596676 3978
rect 596744 3922 596800 3978
rect 596868 3922 596924 3978
rect 596496 -216 596552 -160
rect 596620 -216 596676 -160
rect 596744 -216 596800 -160
rect 596868 -216 596924 -160
rect 596496 -340 596552 -284
rect 596620 -340 596676 -284
rect 596744 -340 596800 -284
rect 596868 -340 596924 -284
rect 596496 -464 596552 -408
rect 596620 -464 596676 -408
rect 596744 -464 596800 -408
rect 596868 -464 596924 -408
rect 596496 -588 596552 -532
rect 596620 -588 596676 -532
rect 596744 -588 596800 -532
rect 596868 -588 596924 -532
rect 597456 586294 597512 586350
rect 597580 586294 597636 586350
rect 597704 586294 597760 586350
rect 597828 586294 597884 586350
rect 597456 586170 597512 586226
rect 597580 586170 597636 586226
rect 597704 586170 597760 586226
rect 597828 586170 597884 586226
rect 597456 586046 597512 586102
rect 597580 586046 597636 586102
rect 597704 586046 597760 586102
rect 597828 586046 597884 586102
rect 597456 585922 597512 585978
rect 597580 585922 597636 585978
rect 597704 585922 597760 585978
rect 597828 585922 597884 585978
rect 597456 568294 597512 568350
rect 597580 568294 597636 568350
rect 597704 568294 597760 568350
rect 597828 568294 597884 568350
rect 597456 568170 597512 568226
rect 597580 568170 597636 568226
rect 597704 568170 597760 568226
rect 597828 568170 597884 568226
rect 597456 568046 597512 568102
rect 597580 568046 597636 568102
rect 597704 568046 597760 568102
rect 597828 568046 597884 568102
rect 597456 567922 597512 567978
rect 597580 567922 597636 567978
rect 597704 567922 597760 567978
rect 597828 567922 597884 567978
rect 597456 550294 597512 550350
rect 597580 550294 597636 550350
rect 597704 550294 597760 550350
rect 597828 550294 597884 550350
rect 597456 550170 597512 550226
rect 597580 550170 597636 550226
rect 597704 550170 597760 550226
rect 597828 550170 597884 550226
rect 597456 550046 597512 550102
rect 597580 550046 597636 550102
rect 597704 550046 597760 550102
rect 597828 550046 597884 550102
rect 597456 549922 597512 549978
rect 597580 549922 597636 549978
rect 597704 549922 597760 549978
rect 597828 549922 597884 549978
rect 597456 532294 597512 532350
rect 597580 532294 597636 532350
rect 597704 532294 597760 532350
rect 597828 532294 597884 532350
rect 597456 532170 597512 532226
rect 597580 532170 597636 532226
rect 597704 532170 597760 532226
rect 597828 532170 597884 532226
rect 597456 532046 597512 532102
rect 597580 532046 597636 532102
rect 597704 532046 597760 532102
rect 597828 532046 597884 532102
rect 597456 531922 597512 531978
rect 597580 531922 597636 531978
rect 597704 531922 597760 531978
rect 597828 531922 597884 531978
rect 597456 514294 597512 514350
rect 597580 514294 597636 514350
rect 597704 514294 597760 514350
rect 597828 514294 597884 514350
rect 597456 514170 597512 514226
rect 597580 514170 597636 514226
rect 597704 514170 597760 514226
rect 597828 514170 597884 514226
rect 597456 514046 597512 514102
rect 597580 514046 597636 514102
rect 597704 514046 597760 514102
rect 597828 514046 597884 514102
rect 597456 513922 597512 513978
rect 597580 513922 597636 513978
rect 597704 513922 597760 513978
rect 597828 513922 597884 513978
rect 597456 496294 597512 496350
rect 597580 496294 597636 496350
rect 597704 496294 597760 496350
rect 597828 496294 597884 496350
rect 597456 496170 597512 496226
rect 597580 496170 597636 496226
rect 597704 496170 597760 496226
rect 597828 496170 597884 496226
rect 597456 496046 597512 496102
rect 597580 496046 597636 496102
rect 597704 496046 597760 496102
rect 597828 496046 597884 496102
rect 597456 495922 597512 495978
rect 597580 495922 597636 495978
rect 597704 495922 597760 495978
rect 597828 495922 597884 495978
rect 597456 478294 597512 478350
rect 597580 478294 597636 478350
rect 597704 478294 597760 478350
rect 597828 478294 597884 478350
rect 597456 478170 597512 478226
rect 597580 478170 597636 478226
rect 597704 478170 597760 478226
rect 597828 478170 597884 478226
rect 597456 478046 597512 478102
rect 597580 478046 597636 478102
rect 597704 478046 597760 478102
rect 597828 478046 597884 478102
rect 597456 477922 597512 477978
rect 597580 477922 597636 477978
rect 597704 477922 597760 477978
rect 597828 477922 597884 477978
rect 597456 460294 597512 460350
rect 597580 460294 597636 460350
rect 597704 460294 597760 460350
rect 597828 460294 597884 460350
rect 597456 460170 597512 460226
rect 597580 460170 597636 460226
rect 597704 460170 597760 460226
rect 597828 460170 597884 460226
rect 597456 460046 597512 460102
rect 597580 460046 597636 460102
rect 597704 460046 597760 460102
rect 597828 460046 597884 460102
rect 597456 459922 597512 459978
rect 597580 459922 597636 459978
rect 597704 459922 597760 459978
rect 597828 459922 597884 459978
rect 597456 442294 597512 442350
rect 597580 442294 597636 442350
rect 597704 442294 597760 442350
rect 597828 442294 597884 442350
rect 597456 442170 597512 442226
rect 597580 442170 597636 442226
rect 597704 442170 597760 442226
rect 597828 442170 597884 442226
rect 597456 442046 597512 442102
rect 597580 442046 597636 442102
rect 597704 442046 597760 442102
rect 597828 442046 597884 442102
rect 597456 441922 597512 441978
rect 597580 441922 597636 441978
rect 597704 441922 597760 441978
rect 597828 441922 597884 441978
rect 597456 424294 597512 424350
rect 597580 424294 597636 424350
rect 597704 424294 597760 424350
rect 597828 424294 597884 424350
rect 597456 424170 597512 424226
rect 597580 424170 597636 424226
rect 597704 424170 597760 424226
rect 597828 424170 597884 424226
rect 597456 424046 597512 424102
rect 597580 424046 597636 424102
rect 597704 424046 597760 424102
rect 597828 424046 597884 424102
rect 597456 423922 597512 423978
rect 597580 423922 597636 423978
rect 597704 423922 597760 423978
rect 597828 423922 597884 423978
rect 597456 406294 597512 406350
rect 597580 406294 597636 406350
rect 597704 406294 597760 406350
rect 597828 406294 597884 406350
rect 597456 406170 597512 406226
rect 597580 406170 597636 406226
rect 597704 406170 597760 406226
rect 597828 406170 597884 406226
rect 597456 406046 597512 406102
rect 597580 406046 597636 406102
rect 597704 406046 597760 406102
rect 597828 406046 597884 406102
rect 597456 405922 597512 405978
rect 597580 405922 597636 405978
rect 597704 405922 597760 405978
rect 597828 405922 597884 405978
rect 597456 388294 597512 388350
rect 597580 388294 597636 388350
rect 597704 388294 597760 388350
rect 597828 388294 597884 388350
rect 597456 388170 597512 388226
rect 597580 388170 597636 388226
rect 597704 388170 597760 388226
rect 597828 388170 597884 388226
rect 597456 388046 597512 388102
rect 597580 388046 597636 388102
rect 597704 388046 597760 388102
rect 597828 388046 597884 388102
rect 597456 387922 597512 387978
rect 597580 387922 597636 387978
rect 597704 387922 597760 387978
rect 597828 387922 597884 387978
rect 597456 370294 597512 370350
rect 597580 370294 597636 370350
rect 597704 370294 597760 370350
rect 597828 370294 597884 370350
rect 597456 370170 597512 370226
rect 597580 370170 597636 370226
rect 597704 370170 597760 370226
rect 597828 370170 597884 370226
rect 597456 370046 597512 370102
rect 597580 370046 597636 370102
rect 597704 370046 597760 370102
rect 597828 370046 597884 370102
rect 597456 369922 597512 369978
rect 597580 369922 597636 369978
rect 597704 369922 597760 369978
rect 597828 369922 597884 369978
rect 597456 352294 597512 352350
rect 597580 352294 597636 352350
rect 597704 352294 597760 352350
rect 597828 352294 597884 352350
rect 597456 352170 597512 352226
rect 597580 352170 597636 352226
rect 597704 352170 597760 352226
rect 597828 352170 597884 352226
rect 597456 352046 597512 352102
rect 597580 352046 597636 352102
rect 597704 352046 597760 352102
rect 597828 352046 597884 352102
rect 597456 351922 597512 351978
rect 597580 351922 597636 351978
rect 597704 351922 597760 351978
rect 597828 351922 597884 351978
rect 597456 334294 597512 334350
rect 597580 334294 597636 334350
rect 597704 334294 597760 334350
rect 597828 334294 597884 334350
rect 597456 334170 597512 334226
rect 597580 334170 597636 334226
rect 597704 334170 597760 334226
rect 597828 334170 597884 334226
rect 597456 334046 597512 334102
rect 597580 334046 597636 334102
rect 597704 334046 597760 334102
rect 597828 334046 597884 334102
rect 597456 333922 597512 333978
rect 597580 333922 597636 333978
rect 597704 333922 597760 333978
rect 597828 333922 597884 333978
rect 597456 316294 597512 316350
rect 597580 316294 597636 316350
rect 597704 316294 597760 316350
rect 597828 316294 597884 316350
rect 597456 316170 597512 316226
rect 597580 316170 597636 316226
rect 597704 316170 597760 316226
rect 597828 316170 597884 316226
rect 597456 316046 597512 316102
rect 597580 316046 597636 316102
rect 597704 316046 597760 316102
rect 597828 316046 597884 316102
rect 597456 315922 597512 315978
rect 597580 315922 597636 315978
rect 597704 315922 597760 315978
rect 597828 315922 597884 315978
rect 597456 298294 597512 298350
rect 597580 298294 597636 298350
rect 597704 298294 597760 298350
rect 597828 298294 597884 298350
rect 597456 298170 597512 298226
rect 597580 298170 597636 298226
rect 597704 298170 597760 298226
rect 597828 298170 597884 298226
rect 597456 298046 597512 298102
rect 597580 298046 597636 298102
rect 597704 298046 597760 298102
rect 597828 298046 597884 298102
rect 597456 297922 597512 297978
rect 597580 297922 597636 297978
rect 597704 297922 597760 297978
rect 597828 297922 597884 297978
rect 597456 280294 597512 280350
rect 597580 280294 597636 280350
rect 597704 280294 597760 280350
rect 597828 280294 597884 280350
rect 597456 280170 597512 280226
rect 597580 280170 597636 280226
rect 597704 280170 597760 280226
rect 597828 280170 597884 280226
rect 597456 280046 597512 280102
rect 597580 280046 597636 280102
rect 597704 280046 597760 280102
rect 597828 280046 597884 280102
rect 597456 279922 597512 279978
rect 597580 279922 597636 279978
rect 597704 279922 597760 279978
rect 597828 279922 597884 279978
rect 597456 262294 597512 262350
rect 597580 262294 597636 262350
rect 597704 262294 597760 262350
rect 597828 262294 597884 262350
rect 597456 262170 597512 262226
rect 597580 262170 597636 262226
rect 597704 262170 597760 262226
rect 597828 262170 597884 262226
rect 597456 262046 597512 262102
rect 597580 262046 597636 262102
rect 597704 262046 597760 262102
rect 597828 262046 597884 262102
rect 597456 261922 597512 261978
rect 597580 261922 597636 261978
rect 597704 261922 597760 261978
rect 597828 261922 597884 261978
rect 597456 244294 597512 244350
rect 597580 244294 597636 244350
rect 597704 244294 597760 244350
rect 597828 244294 597884 244350
rect 597456 244170 597512 244226
rect 597580 244170 597636 244226
rect 597704 244170 597760 244226
rect 597828 244170 597884 244226
rect 597456 244046 597512 244102
rect 597580 244046 597636 244102
rect 597704 244046 597760 244102
rect 597828 244046 597884 244102
rect 597456 243922 597512 243978
rect 597580 243922 597636 243978
rect 597704 243922 597760 243978
rect 597828 243922 597884 243978
rect 597456 226294 597512 226350
rect 597580 226294 597636 226350
rect 597704 226294 597760 226350
rect 597828 226294 597884 226350
rect 597456 226170 597512 226226
rect 597580 226170 597636 226226
rect 597704 226170 597760 226226
rect 597828 226170 597884 226226
rect 597456 226046 597512 226102
rect 597580 226046 597636 226102
rect 597704 226046 597760 226102
rect 597828 226046 597884 226102
rect 597456 225922 597512 225978
rect 597580 225922 597636 225978
rect 597704 225922 597760 225978
rect 597828 225922 597884 225978
rect 597456 208294 597512 208350
rect 597580 208294 597636 208350
rect 597704 208294 597760 208350
rect 597828 208294 597884 208350
rect 597456 208170 597512 208226
rect 597580 208170 597636 208226
rect 597704 208170 597760 208226
rect 597828 208170 597884 208226
rect 597456 208046 597512 208102
rect 597580 208046 597636 208102
rect 597704 208046 597760 208102
rect 597828 208046 597884 208102
rect 597456 207922 597512 207978
rect 597580 207922 597636 207978
rect 597704 207922 597760 207978
rect 597828 207922 597884 207978
rect 597456 190294 597512 190350
rect 597580 190294 597636 190350
rect 597704 190294 597760 190350
rect 597828 190294 597884 190350
rect 597456 190170 597512 190226
rect 597580 190170 597636 190226
rect 597704 190170 597760 190226
rect 597828 190170 597884 190226
rect 597456 190046 597512 190102
rect 597580 190046 597636 190102
rect 597704 190046 597760 190102
rect 597828 190046 597884 190102
rect 597456 189922 597512 189978
rect 597580 189922 597636 189978
rect 597704 189922 597760 189978
rect 597828 189922 597884 189978
rect 597456 172294 597512 172350
rect 597580 172294 597636 172350
rect 597704 172294 597760 172350
rect 597828 172294 597884 172350
rect 597456 172170 597512 172226
rect 597580 172170 597636 172226
rect 597704 172170 597760 172226
rect 597828 172170 597884 172226
rect 597456 172046 597512 172102
rect 597580 172046 597636 172102
rect 597704 172046 597760 172102
rect 597828 172046 597884 172102
rect 597456 171922 597512 171978
rect 597580 171922 597636 171978
rect 597704 171922 597760 171978
rect 597828 171922 597884 171978
rect 597456 154294 597512 154350
rect 597580 154294 597636 154350
rect 597704 154294 597760 154350
rect 597828 154294 597884 154350
rect 597456 154170 597512 154226
rect 597580 154170 597636 154226
rect 597704 154170 597760 154226
rect 597828 154170 597884 154226
rect 597456 154046 597512 154102
rect 597580 154046 597636 154102
rect 597704 154046 597760 154102
rect 597828 154046 597884 154102
rect 597456 153922 597512 153978
rect 597580 153922 597636 153978
rect 597704 153922 597760 153978
rect 597828 153922 597884 153978
rect 597456 136294 597512 136350
rect 597580 136294 597636 136350
rect 597704 136294 597760 136350
rect 597828 136294 597884 136350
rect 597456 136170 597512 136226
rect 597580 136170 597636 136226
rect 597704 136170 597760 136226
rect 597828 136170 597884 136226
rect 597456 136046 597512 136102
rect 597580 136046 597636 136102
rect 597704 136046 597760 136102
rect 597828 136046 597884 136102
rect 597456 135922 597512 135978
rect 597580 135922 597636 135978
rect 597704 135922 597760 135978
rect 597828 135922 597884 135978
rect 597456 118294 597512 118350
rect 597580 118294 597636 118350
rect 597704 118294 597760 118350
rect 597828 118294 597884 118350
rect 597456 118170 597512 118226
rect 597580 118170 597636 118226
rect 597704 118170 597760 118226
rect 597828 118170 597884 118226
rect 597456 118046 597512 118102
rect 597580 118046 597636 118102
rect 597704 118046 597760 118102
rect 597828 118046 597884 118102
rect 597456 117922 597512 117978
rect 597580 117922 597636 117978
rect 597704 117922 597760 117978
rect 597828 117922 597884 117978
rect 597456 100294 597512 100350
rect 597580 100294 597636 100350
rect 597704 100294 597760 100350
rect 597828 100294 597884 100350
rect 597456 100170 597512 100226
rect 597580 100170 597636 100226
rect 597704 100170 597760 100226
rect 597828 100170 597884 100226
rect 597456 100046 597512 100102
rect 597580 100046 597636 100102
rect 597704 100046 597760 100102
rect 597828 100046 597884 100102
rect 597456 99922 597512 99978
rect 597580 99922 597636 99978
rect 597704 99922 597760 99978
rect 597828 99922 597884 99978
rect 597456 82294 597512 82350
rect 597580 82294 597636 82350
rect 597704 82294 597760 82350
rect 597828 82294 597884 82350
rect 597456 82170 597512 82226
rect 597580 82170 597636 82226
rect 597704 82170 597760 82226
rect 597828 82170 597884 82226
rect 597456 82046 597512 82102
rect 597580 82046 597636 82102
rect 597704 82046 597760 82102
rect 597828 82046 597884 82102
rect 597456 81922 597512 81978
rect 597580 81922 597636 81978
rect 597704 81922 597760 81978
rect 597828 81922 597884 81978
rect 597456 64294 597512 64350
rect 597580 64294 597636 64350
rect 597704 64294 597760 64350
rect 597828 64294 597884 64350
rect 597456 64170 597512 64226
rect 597580 64170 597636 64226
rect 597704 64170 597760 64226
rect 597828 64170 597884 64226
rect 597456 64046 597512 64102
rect 597580 64046 597636 64102
rect 597704 64046 597760 64102
rect 597828 64046 597884 64102
rect 597456 63922 597512 63978
rect 597580 63922 597636 63978
rect 597704 63922 597760 63978
rect 597828 63922 597884 63978
rect 597456 46294 597512 46350
rect 597580 46294 597636 46350
rect 597704 46294 597760 46350
rect 597828 46294 597884 46350
rect 597456 46170 597512 46226
rect 597580 46170 597636 46226
rect 597704 46170 597760 46226
rect 597828 46170 597884 46226
rect 597456 46046 597512 46102
rect 597580 46046 597636 46102
rect 597704 46046 597760 46102
rect 597828 46046 597884 46102
rect 597456 45922 597512 45978
rect 597580 45922 597636 45978
rect 597704 45922 597760 45978
rect 597828 45922 597884 45978
rect 597456 28294 597512 28350
rect 597580 28294 597636 28350
rect 597704 28294 597760 28350
rect 597828 28294 597884 28350
rect 597456 28170 597512 28226
rect 597580 28170 597636 28226
rect 597704 28170 597760 28226
rect 597828 28170 597884 28226
rect 597456 28046 597512 28102
rect 597580 28046 597636 28102
rect 597704 28046 597760 28102
rect 597828 28046 597884 28102
rect 597456 27922 597512 27978
rect 597580 27922 597636 27978
rect 597704 27922 597760 27978
rect 597828 27922 597884 27978
rect 597456 10294 597512 10350
rect 597580 10294 597636 10350
rect 597704 10294 597760 10350
rect 597828 10294 597884 10350
rect 597456 10170 597512 10226
rect 597580 10170 597636 10226
rect 597704 10170 597760 10226
rect 597828 10170 597884 10226
rect 597456 10046 597512 10102
rect 597580 10046 597636 10102
rect 597704 10046 597760 10102
rect 597828 10046 597884 10102
rect 597456 9922 597512 9978
rect 597580 9922 597636 9978
rect 597704 9922 597760 9978
rect 597828 9922 597884 9978
rect 592914 -1176 592970 -1120
rect 593038 -1176 593094 -1120
rect 593162 -1176 593218 -1120
rect 593286 -1176 593342 -1120
rect 592914 -1300 592970 -1244
rect 593038 -1300 593094 -1244
rect 593162 -1300 593218 -1244
rect 593286 -1300 593342 -1244
rect 592914 -1424 592970 -1368
rect 593038 -1424 593094 -1368
rect 593162 -1424 593218 -1368
rect 593286 -1424 593342 -1368
rect 592914 -1548 592970 -1492
rect 593038 -1548 593094 -1492
rect 593162 -1548 593218 -1492
rect 593286 -1548 593342 -1492
rect 597456 -1176 597512 -1120
rect 597580 -1176 597636 -1120
rect 597704 -1176 597760 -1120
rect 597828 -1176 597884 -1120
rect 597456 -1300 597512 -1244
rect 597580 -1300 597636 -1244
rect 597704 -1300 597760 -1244
rect 597828 -1300 597884 -1244
rect 597456 -1424 597512 -1368
rect 597580 -1424 597636 -1368
rect 597704 -1424 597760 -1368
rect 597828 -1424 597884 -1368
rect 597456 -1548 597512 -1492
rect 597580 -1548 597636 -1492
rect 597704 -1548 597760 -1492
rect 597828 -1548 597884 -1492
<< metal5 >>
rect -1916 598172 597980 598268
rect -1916 598116 -1820 598172
rect -1764 598116 -1696 598172
rect -1640 598116 -1572 598172
rect -1516 598116 -1448 598172
rect -1392 598116 9234 598172
rect 9290 598116 9358 598172
rect 9414 598116 9482 598172
rect 9538 598116 9606 598172
rect 9662 598116 39954 598172
rect 40010 598116 40078 598172
rect 40134 598116 40202 598172
rect 40258 598116 40326 598172
rect 40382 598116 70674 598172
rect 70730 598116 70798 598172
rect 70854 598116 70922 598172
rect 70978 598116 71046 598172
rect 71102 598116 101394 598172
rect 101450 598116 101518 598172
rect 101574 598116 101642 598172
rect 101698 598116 101766 598172
rect 101822 598116 132114 598172
rect 132170 598116 132238 598172
rect 132294 598116 132362 598172
rect 132418 598116 132486 598172
rect 132542 598116 162834 598172
rect 162890 598116 162958 598172
rect 163014 598116 163082 598172
rect 163138 598116 163206 598172
rect 163262 598116 193554 598172
rect 193610 598116 193678 598172
rect 193734 598116 193802 598172
rect 193858 598116 193926 598172
rect 193982 598116 224274 598172
rect 224330 598116 224398 598172
rect 224454 598116 224522 598172
rect 224578 598116 224646 598172
rect 224702 598116 254994 598172
rect 255050 598116 255118 598172
rect 255174 598116 255242 598172
rect 255298 598116 255366 598172
rect 255422 598116 285714 598172
rect 285770 598116 285838 598172
rect 285894 598116 285962 598172
rect 286018 598116 286086 598172
rect 286142 598116 316434 598172
rect 316490 598116 316558 598172
rect 316614 598116 316682 598172
rect 316738 598116 316806 598172
rect 316862 598116 347154 598172
rect 347210 598116 347278 598172
rect 347334 598116 347402 598172
rect 347458 598116 347526 598172
rect 347582 598116 377874 598172
rect 377930 598116 377998 598172
rect 378054 598116 378122 598172
rect 378178 598116 378246 598172
rect 378302 598116 408594 598172
rect 408650 598116 408718 598172
rect 408774 598116 408842 598172
rect 408898 598116 408966 598172
rect 409022 598116 439314 598172
rect 439370 598116 439438 598172
rect 439494 598116 439562 598172
rect 439618 598116 439686 598172
rect 439742 598116 470034 598172
rect 470090 598116 470158 598172
rect 470214 598116 470282 598172
rect 470338 598116 470406 598172
rect 470462 598116 500754 598172
rect 500810 598116 500878 598172
rect 500934 598116 501002 598172
rect 501058 598116 501126 598172
rect 501182 598116 531474 598172
rect 531530 598116 531598 598172
rect 531654 598116 531722 598172
rect 531778 598116 531846 598172
rect 531902 598116 562194 598172
rect 562250 598116 562318 598172
rect 562374 598116 562442 598172
rect 562498 598116 562566 598172
rect 562622 598116 592914 598172
rect 592970 598116 593038 598172
rect 593094 598116 593162 598172
rect 593218 598116 593286 598172
rect 593342 598116 597456 598172
rect 597512 598116 597580 598172
rect 597636 598116 597704 598172
rect 597760 598116 597828 598172
rect 597884 598116 597980 598172
rect -1916 598048 597980 598116
rect -1916 597992 -1820 598048
rect -1764 597992 -1696 598048
rect -1640 597992 -1572 598048
rect -1516 597992 -1448 598048
rect -1392 597992 9234 598048
rect 9290 597992 9358 598048
rect 9414 597992 9482 598048
rect 9538 597992 9606 598048
rect 9662 597992 39954 598048
rect 40010 597992 40078 598048
rect 40134 597992 40202 598048
rect 40258 597992 40326 598048
rect 40382 597992 70674 598048
rect 70730 597992 70798 598048
rect 70854 597992 70922 598048
rect 70978 597992 71046 598048
rect 71102 597992 101394 598048
rect 101450 597992 101518 598048
rect 101574 597992 101642 598048
rect 101698 597992 101766 598048
rect 101822 597992 132114 598048
rect 132170 597992 132238 598048
rect 132294 597992 132362 598048
rect 132418 597992 132486 598048
rect 132542 597992 162834 598048
rect 162890 597992 162958 598048
rect 163014 597992 163082 598048
rect 163138 597992 163206 598048
rect 163262 597992 193554 598048
rect 193610 597992 193678 598048
rect 193734 597992 193802 598048
rect 193858 597992 193926 598048
rect 193982 597992 224274 598048
rect 224330 597992 224398 598048
rect 224454 597992 224522 598048
rect 224578 597992 224646 598048
rect 224702 597992 254994 598048
rect 255050 597992 255118 598048
rect 255174 597992 255242 598048
rect 255298 597992 255366 598048
rect 255422 597992 285714 598048
rect 285770 597992 285838 598048
rect 285894 597992 285962 598048
rect 286018 597992 286086 598048
rect 286142 597992 316434 598048
rect 316490 597992 316558 598048
rect 316614 597992 316682 598048
rect 316738 597992 316806 598048
rect 316862 597992 347154 598048
rect 347210 597992 347278 598048
rect 347334 597992 347402 598048
rect 347458 597992 347526 598048
rect 347582 597992 377874 598048
rect 377930 597992 377998 598048
rect 378054 597992 378122 598048
rect 378178 597992 378246 598048
rect 378302 597992 408594 598048
rect 408650 597992 408718 598048
rect 408774 597992 408842 598048
rect 408898 597992 408966 598048
rect 409022 597992 439314 598048
rect 439370 597992 439438 598048
rect 439494 597992 439562 598048
rect 439618 597992 439686 598048
rect 439742 597992 470034 598048
rect 470090 597992 470158 598048
rect 470214 597992 470282 598048
rect 470338 597992 470406 598048
rect 470462 597992 500754 598048
rect 500810 597992 500878 598048
rect 500934 597992 501002 598048
rect 501058 597992 501126 598048
rect 501182 597992 531474 598048
rect 531530 597992 531598 598048
rect 531654 597992 531722 598048
rect 531778 597992 531846 598048
rect 531902 597992 562194 598048
rect 562250 597992 562318 598048
rect 562374 597992 562442 598048
rect 562498 597992 562566 598048
rect 562622 597992 592914 598048
rect 592970 597992 593038 598048
rect 593094 597992 593162 598048
rect 593218 597992 593286 598048
rect 593342 597992 597456 598048
rect 597512 597992 597580 598048
rect 597636 597992 597704 598048
rect 597760 597992 597828 598048
rect 597884 597992 597980 598048
rect -1916 597924 597980 597992
rect -1916 597868 -1820 597924
rect -1764 597868 -1696 597924
rect -1640 597868 -1572 597924
rect -1516 597868 -1448 597924
rect -1392 597868 9234 597924
rect 9290 597868 9358 597924
rect 9414 597868 9482 597924
rect 9538 597868 9606 597924
rect 9662 597868 39954 597924
rect 40010 597868 40078 597924
rect 40134 597868 40202 597924
rect 40258 597868 40326 597924
rect 40382 597868 70674 597924
rect 70730 597868 70798 597924
rect 70854 597868 70922 597924
rect 70978 597868 71046 597924
rect 71102 597868 101394 597924
rect 101450 597868 101518 597924
rect 101574 597868 101642 597924
rect 101698 597868 101766 597924
rect 101822 597868 132114 597924
rect 132170 597868 132238 597924
rect 132294 597868 132362 597924
rect 132418 597868 132486 597924
rect 132542 597868 162834 597924
rect 162890 597868 162958 597924
rect 163014 597868 163082 597924
rect 163138 597868 163206 597924
rect 163262 597868 193554 597924
rect 193610 597868 193678 597924
rect 193734 597868 193802 597924
rect 193858 597868 193926 597924
rect 193982 597868 224274 597924
rect 224330 597868 224398 597924
rect 224454 597868 224522 597924
rect 224578 597868 224646 597924
rect 224702 597868 254994 597924
rect 255050 597868 255118 597924
rect 255174 597868 255242 597924
rect 255298 597868 255366 597924
rect 255422 597868 285714 597924
rect 285770 597868 285838 597924
rect 285894 597868 285962 597924
rect 286018 597868 286086 597924
rect 286142 597868 316434 597924
rect 316490 597868 316558 597924
rect 316614 597868 316682 597924
rect 316738 597868 316806 597924
rect 316862 597868 347154 597924
rect 347210 597868 347278 597924
rect 347334 597868 347402 597924
rect 347458 597868 347526 597924
rect 347582 597868 377874 597924
rect 377930 597868 377998 597924
rect 378054 597868 378122 597924
rect 378178 597868 378246 597924
rect 378302 597868 408594 597924
rect 408650 597868 408718 597924
rect 408774 597868 408842 597924
rect 408898 597868 408966 597924
rect 409022 597868 439314 597924
rect 439370 597868 439438 597924
rect 439494 597868 439562 597924
rect 439618 597868 439686 597924
rect 439742 597868 470034 597924
rect 470090 597868 470158 597924
rect 470214 597868 470282 597924
rect 470338 597868 470406 597924
rect 470462 597868 500754 597924
rect 500810 597868 500878 597924
rect 500934 597868 501002 597924
rect 501058 597868 501126 597924
rect 501182 597868 531474 597924
rect 531530 597868 531598 597924
rect 531654 597868 531722 597924
rect 531778 597868 531846 597924
rect 531902 597868 562194 597924
rect 562250 597868 562318 597924
rect 562374 597868 562442 597924
rect 562498 597868 562566 597924
rect 562622 597868 592914 597924
rect 592970 597868 593038 597924
rect 593094 597868 593162 597924
rect 593218 597868 593286 597924
rect 593342 597868 597456 597924
rect 597512 597868 597580 597924
rect 597636 597868 597704 597924
rect 597760 597868 597828 597924
rect 597884 597868 597980 597924
rect -1916 597800 597980 597868
rect -1916 597744 -1820 597800
rect -1764 597744 -1696 597800
rect -1640 597744 -1572 597800
rect -1516 597744 -1448 597800
rect -1392 597744 9234 597800
rect 9290 597744 9358 597800
rect 9414 597744 9482 597800
rect 9538 597744 9606 597800
rect 9662 597744 39954 597800
rect 40010 597744 40078 597800
rect 40134 597744 40202 597800
rect 40258 597744 40326 597800
rect 40382 597744 70674 597800
rect 70730 597744 70798 597800
rect 70854 597744 70922 597800
rect 70978 597744 71046 597800
rect 71102 597744 101394 597800
rect 101450 597744 101518 597800
rect 101574 597744 101642 597800
rect 101698 597744 101766 597800
rect 101822 597744 132114 597800
rect 132170 597744 132238 597800
rect 132294 597744 132362 597800
rect 132418 597744 132486 597800
rect 132542 597744 162834 597800
rect 162890 597744 162958 597800
rect 163014 597744 163082 597800
rect 163138 597744 163206 597800
rect 163262 597744 193554 597800
rect 193610 597744 193678 597800
rect 193734 597744 193802 597800
rect 193858 597744 193926 597800
rect 193982 597744 224274 597800
rect 224330 597744 224398 597800
rect 224454 597744 224522 597800
rect 224578 597744 224646 597800
rect 224702 597744 254994 597800
rect 255050 597744 255118 597800
rect 255174 597744 255242 597800
rect 255298 597744 255366 597800
rect 255422 597744 285714 597800
rect 285770 597744 285838 597800
rect 285894 597744 285962 597800
rect 286018 597744 286086 597800
rect 286142 597744 316434 597800
rect 316490 597744 316558 597800
rect 316614 597744 316682 597800
rect 316738 597744 316806 597800
rect 316862 597744 347154 597800
rect 347210 597744 347278 597800
rect 347334 597744 347402 597800
rect 347458 597744 347526 597800
rect 347582 597744 377874 597800
rect 377930 597744 377998 597800
rect 378054 597744 378122 597800
rect 378178 597744 378246 597800
rect 378302 597744 408594 597800
rect 408650 597744 408718 597800
rect 408774 597744 408842 597800
rect 408898 597744 408966 597800
rect 409022 597744 439314 597800
rect 439370 597744 439438 597800
rect 439494 597744 439562 597800
rect 439618 597744 439686 597800
rect 439742 597744 470034 597800
rect 470090 597744 470158 597800
rect 470214 597744 470282 597800
rect 470338 597744 470406 597800
rect 470462 597744 500754 597800
rect 500810 597744 500878 597800
rect 500934 597744 501002 597800
rect 501058 597744 501126 597800
rect 501182 597744 531474 597800
rect 531530 597744 531598 597800
rect 531654 597744 531722 597800
rect 531778 597744 531846 597800
rect 531902 597744 562194 597800
rect 562250 597744 562318 597800
rect 562374 597744 562442 597800
rect 562498 597744 562566 597800
rect 562622 597744 592914 597800
rect 592970 597744 593038 597800
rect 593094 597744 593162 597800
rect 593218 597744 593286 597800
rect 593342 597744 597456 597800
rect 597512 597744 597580 597800
rect 597636 597744 597704 597800
rect 597760 597744 597828 597800
rect 597884 597744 597980 597800
rect -1916 597648 597980 597744
rect -956 597212 597020 597308
rect -956 597156 -860 597212
rect -804 597156 -736 597212
rect -680 597156 -612 597212
rect -556 597156 -488 597212
rect -432 597156 5514 597212
rect 5570 597156 5638 597212
rect 5694 597156 5762 597212
rect 5818 597156 5886 597212
rect 5942 597156 36234 597212
rect 36290 597156 36358 597212
rect 36414 597156 36482 597212
rect 36538 597156 36606 597212
rect 36662 597156 66954 597212
rect 67010 597156 67078 597212
rect 67134 597156 67202 597212
rect 67258 597156 67326 597212
rect 67382 597156 97674 597212
rect 97730 597156 97798 597212
rect 97854 597156 97922 597212
rect 97978 597156 98046 597212
rect 98102 597156 128394 597212
rect 128450 597156 128518 597212
rect 128574 597156 128642 597212
rect 128698 597156 128766 597212
rect 128822 597156 159114 597212
rect 159170 597156 159238 597212
rect 159294 597156 159362 597212
rect 159418 597156 159486 597212
rect 159542 597156 189834 597212
rect 189890 597156 189958 597212
rect 190014 597156 190082 597212
rect 190138 597156 190206 597212
rect 190262 597156 220554 597212
rect 220610 597156 220678 597212
rect 220734 597156 220802 597212
rect 220858 597156 220926 597212
rect 220982 597156 251274 597212
rect 251330 597156 251398 597212
rect 251454 597156 251522 597212
rect 251578 597156 251646 597212
rect 251702 597156 281994 597212
rect 282050 597156 282118 597212
rect 282174 597156 282242 597212
rect 282298 597156 282366 597212
rect 282422 597156 312714 597212
rect 312770 597156 312838 597212
rect 312894 597156 312962 597212
rect 313018 597156 313086 597212
rect 313142 597156 343434 597212
rect 343490 597156 343558 597212
rect 343614 597156 343682 597212
rect 343738 597156 343806 597212
rect 343862 597156 374154 597212
rect 374210 597156 374278 597212
rect 374334 597156 374402 597212
rect 374458 597156 374526 597212
rect 374582 597156 404874 597212
rect 404930 597156 404998 597212
rect 405054 597156 405122 597212
rect 405178 597156 405246 597212
rect 405302 597156 435594 597212
rect 435650 597156 435718 597212
rect 435774 597156 435842 597212
rect 435898 597156 435966 597212
rect 436022 597156 466314 597212
rect 466370 597156 466438 597212
rect 466494 597156 466562 597212
rect 466618 597156 466686 597212
rect 466742 597156 497034 597212
rect 497090 597156 497158 597212
rect 497214 597156 497282 597212
rect 497338 597156 497406 597212
rect 497462 597156 527754 597212
rect 527810 597156 527878 597212
rect 527934 597156 528002 597212
rect 528058 597156 528126 597212
rect 528182 597156 558474 597212
rect 558530 597156 558598 597212
rect 558654 597156 558722 597212
rect 558778 597156 558846 597212
rect 558902 597156 589194 597212
rect 589250 597156 589318 597212
rect 589374 597156 589442 597212
rect 589498 597156 589566 597212
rect 589622 597156 596496 597212
rect 596552 597156 596620 597212
rect 596676 597156 596744 597212
rect 596800 597156 596868 597212
rect 596924 597156 597020 597212
rect -956 597088 597020 597156
rect -956 597032 -860 597088
rect -804 597032 -736 597088
rect -680 597032 -612 597088
rect -556 597032 -488 597088
rect -432 597032 5514 597088
rect 5570 597032 5638 597088
rect 5694 597032 5762 597088
rect 5818 597032 5886 597088
rect 5942 597032 36234 597088
rect 36290 597032 36358 597088
rect 36414 597032 36482 597088
rect 36538 597032 36606 597088
rect 36662 597032 66954 597088
rect 67010 597032 67078 597088
rect 67134 597032 67202 597088
rect 67258 597032 67326 597088
rect 67382 597032 97674 597088
rect 97730 597032 97798 597088
rect 97854 597032 97922 597088
rect 97978 597032 98046 597088
rect 98102 597032 128394 597088
rect 128450 597032 128518 597088
rect 128574 597032 128642 597088
rect 128698 597032 128766 597088
rect 128822 597032 159114 597088
rect 159170 597032 159238 597088
rect 159294 597032 159362 597088
rect 159418 597032 159486 597088
rect 159542 597032 189834 597088
rect 189890 597032 189958 597088
rect 190014 597032 190082 597088
rect 190138 597032 190206 597088
rect 190262 597032 220554 597088
rect 220610 597032 220678 597088
rect 220734 597032 220802 597088
rect 220858 597032 220926 597088
rect 220982 597032 251274 597088
rect 251330 597032 251398 597088
rect 251454 597032 251522 597088
rect 251578 597032 251646 597088
rect 251702 597032 281994 597088
rect 282050 597032 282118 597088
rect 282174 597032 282242 597088
rect 282298 597032 282366 597088
rect 282422 597032 312714 597088
rect 312770 597032 312838 597088
rect 312894 597032 312962 597088
rect 313018 597032 313086 597088
rect 313142 597032 343434 597088
rect 343490 597032 343558 597088
rect 343614 597032 343682 597088
rect 343738 597032 343806 597088
rect 343862 597032 374154 597088
rect 374210 597032 374278 597088
rect 374334 597032 374402 597088
rect 374458 597032 374526 597088
rect 374582 597032 404874 597088
rect 404930 597032 404998 597088
rect 405054 597032 405122 597088
rect 405178 597032 405246 597088
rect 405302 597032 435594 597088
rect 435650 597032 435718 597088
rect 435774 597032 435842 597088
rect 435898 597032 435966 597088
rect 436022 597032 466314 597088
rect 466370 597032 466438 597088
rect 466494 597032 466562 597088
rect 466618 597032 466686 597088
rect 466742 597032 497034 597088
rect 497090 597032 497158 597088
rect 497214 597032 497282 597088
rect 497338 597032 497406 597088
rect 497462 597032 527754 597088
rect 527810 597032 527878 597088
rect 527934 597032 528002 597088
rect 528058 597032 528126 597088
rect 528182 597032 558474 597088
rect 558530 597032 558598 597088
rect 558654 597032 558722 597088
rect 558778 597032 558846 597088
rect 558902 597032 589194 597088
rect 589250 597032 589318 597088
rect 589374 597032 589442 597088
rect 589498 597032 589566 597088
rect 589622 597032 596496 597088
rect 596552 597032 596620 597088
rect 596676 597032 596744 597088
rect 596800 597032 596868 597088
rect 596924 597032 597020 597088
rect -956 596964 597020 597032
rect -956 596908 -860 596964
rect -804 596908 -736 596964
rect -680 596908 -612 596964
rect -556 596908 -488 596964
rect -432 596908 5514 596964
rect 5570 596908 5638 596964
rect 5694 596908 5762 596964
rect 5818 596908 5886 596964
rect 5942 596908 36234 596964
rect 36290 596908 36358 596964
rect 36414 596908 36482 596964
rect 36538 596908 36606 596964
rect 36662 596908 66954 596964
rect 67010 596908 67078 596964
rect 67134 596908 67202 596964
rect 67258 596908 67326 596964
rect 67382 596908 97674 596964
rect 97730 596908 97798 596964
rect 97854 596908 97922 596964
rect 97978 596908 98046 596964
rect 98102 596908 128394 596964
rect 128450 596908 128518 596964
rect 128574 596908 128642 596964
rect 128698 596908 128766 596964
rect 128822 596908 159114 596964
rect 159170 596908 159238 596964
rect 159294 596908 159362 596964
rect 159418 596908 159486 596964
rect 159542 596908 189834 596964
rect 189890 596908 189958 596964
rect 190014 596908 190082 596964
rect 190138 596908 190206 596964
rect 190262 596908 220554 596964
rect 220610 596908 220678 596964
rect 220734 596908 220802 596964
rect 220858 596908 220926 596964
rect 220982 596908 251274 596964
rect 251330 596908 251398 596964
rect 251454 596908 251522 596964
rect 251578 596908 251646 596964
rect 251702 596908 281994 596964
rect 282050 596908 282118 596964
rect 282174 596908 282242 596964
rect 282298 596908 282366 596964
rect 282422 596908 312714 596964
rect 312770 596908 312838 596964
rect 312894 596908 312962 596964
rect 313018 596908 313086 596964
rect 313142 596908 343434 596964
rect 343490 596908 343558 596964
rect 343614 596908 343682 596964
rect 343738 596908 343806 596964
rect 343862 596908 374154 596964
rect 374210 596908 374278 596964
rect 374334 596908 374402 596964
rect 374458 596908 374526 596964
rect 374582 596908 404874 596964
rect 404930 596908 404998 596964
rect 405054 596908 405122 596964
rect 405178 596908 405246 596964
rect 405302 596908 435594 596964
rect 435650 596908 435718 596964
rect 435774 596908 435842 596964
rect 435898 596908 435966 596964
rect 436022 596908 466314 596964
rect 466370 596908 466438 596964
rect 466494 596908 466562 596964
rect 466618 596908 466686 596964
rect 466742 596908 497034 596964
rect 497090 596908 497158 596964
rect 497214 596908 497282 596964
rect 497338 596908 497406 596964
rect 497462 596908 527754 596964
rect 527810 596908 527878 596964
rect 527934 596908 528002 596964
rect 528058 596908 528126 596964
rect 528182 596908 558474 596964
rect 558530 596908 558598 596964
rect 558654 596908 558722 596964
rect 558778 596908 558846 596964
rect 558902 596908 589194 596964
rect 589250 596908 589318 596964
rect 589374 596908 589442 596964
rect 589498 596908 589566 596964
rect 589622 596908 596496 596964
rect 596552 596908 596620 596964
rect 596676 596908 596744 596964
rect 596800 596908 596868 596964
rect 596924 596908 597020 596964
rect -956 596840 597020 596908
rect -956 596784 -860 596840
rect -804 596784 -736 596840
rect -680 596784 -612 596840
rect -556 596784 -488 596840
rect -432 596784 5514 596840
rect 5570 596784 5638 596840
rect 5694 596784 5762 596840
rect 5818 596784 5886 596840
rect 5942 596784 36234 596840
rect 36290 596784 36358 596840
rect 36414 596784 36482 596840
rect 36538 596784 36606 596840
rect 36662 596784 66954 596840
rect 67010 596784 67078 596840
rect 67134 596784 67202 596840
rect 67258 596784 67326 596840
rect 67382 596784 97674 596840
rect 97730 596784 97798 596840
rect 97854 596784 97922 596840
rect 97978 596784 98046 596840
rect 98102 596784 128394 596840
rect 128450 596784 128518 596840
rect 128574 596784 128642 596840
rect 128698 596784 128766 596840
rect 128822 596784 159114 596840
rect 159170 596784 159238 596840
rect 159294 596784 159362 596840
rect 159418 596784 159486 596840
rect 159542 596784 189834 596840
rect 189890 596784 189958 596840
rect 190014 596784 190082 596840
rect 190138 596784 190206 596840
rect 190262 596784 220554 596840
rect 220610 596784 220678 596840
rect 220734 596784 220802 596840
rect 220858 596784 220926 596840
rect 220982 596784 251274 596840
rect 251330 596784 251398 596840
rect 251454 596784 251522 596840
rect 251578 596784 251646 596840
rect 251702 596784 281994 596840
rect 282050 596784 282118 596840
rect 282174 596784 282242 596840
rect 282298 596784 282366 596840
rect 282422 596784 312714 596840
rect 312770 596784 312838 596840
rect 312894 596784 312962 596840
rect 313018 596784 313086 596840
rect 313142 596784 343434 596840
rect 343490 596784 343558 596840
rect 343614 596784 343682 596840
rect 343738 596784 343806 596840
rect 343862 596784 374154 596840
rect 374210 596784 374278 596840
rect 374334 596784 374402 596840
rect 374458 596784 374526 596840
rect 374582 596784 404874 596840
rect 404930 596784 404998 596840
rect 405054 596784 405122 596840
rect 405178 596784 405246 596840
rect 405302 596784 435594 596840
rect 435650 596784 435718 596840
rect 435774 596784 435842 596840
rect 435898 596784 435966 596840
rect 436022 596784 466314 596840
rect 466370 596784 466438 596840
rect 466494 596784 466562 596840
rect 466618 596784 466686 596840
rect 466742 596784 497034 596840
rect 497090 596784 497158 596840
rect 497214 596784 497282 596840
rect 497338 596784 497406 596840
rect 497462 596784 527754 596840
rect 527810 596784 527878 596840
rect 527934 596784 528002 596840
rect 528058 596784 528126 596840
rect 528182 596784 558474 596840
rect 558530 596784 558598 596840
rect 558654 596784 558722 596840
rect 558778 596784 558846 596840
rect 558902 596784 589194 596840
rect 589250 596784 589318 596840
rect 589374 596784 589442 596840
rect 589498 596784 589566 596840
rect 589622 596784 596496 596840
rect 596552 596784 596620 596840
rect 596676 596784 596744 596840
rect 596800 596784 596868 596840
rect 596924 596784 597020 596840
rect -956 596688 597020 596784
rect -1916 586350 597980 586446
rect -1916 586294 -1820 586350
rect -1764 586294 -1696 586350
rect -1640 586294 -1572 586350
rect -1516 586294 -1448 586350
rect -1392 586294 9234 586350
rect 9290 586294 9358 586350
rect 9414 586294 9482 586350
rect 9538 586294 9606 586350
rect 9662 586294 39954 586350
rect 40010 586294 40078 586350
rect 40134 586294 40202 586350
rect 40258 586294 40326 586350
rect 40382 586294 70674 586350
rect 70730 586294 70798 586350
rect 70854 586294 70922 586350
rect 70978 586294 71046 586350
rect 71102 586294 101394 586350
rect 101450 586294 101518 586350
rect 101574 586294 101642 586350
rect 101698 586294 101766 586350
rect 101822 586294 132114 586350
rect 132170 586294 132238 586350
rect 132294 586294 132362 586350
rect 132418 586294 132486 586350
rect 132542 586294 162834 586350
rect 162890 586294 162958 586350
rect 163014 586294 163082 586350
rect 163138 586294 163206 586350
rect 163262 586294 193554 586350
rect 193610 586294 193678 586350
rect 193734 586294 193802 586350
rect 193858 586294 193926 586350
rect 193982 586294 224274 586350
rect 224330 586294 224398 586350
rect 224454 586294 224522 586350
rect 224578 586294 224646 586350
rect 224702 586294 254994 586350
rect 255050 586294 255118 586350
rect 255174 586294 255242 586350
rect 255298 586294 255366 586350
rect 255422 586294 285714 586350
rect 285770 586294 285838 586350
rect 285894 586294 285962 586350
rect 286018 586294 286086 586350
rect 286142 586294 316434 586350
rect 316490 586294 316558 586350
rect 316614 586294 316682 586350
rect 316738 586294 316806 586350
rect 316862 586294 347154 586350
rect 347210 586294 347278 586350
rect 347334 586294 347402 586350
rect 347458 586294 347526 586350
rect 347582 586294 377874 586350
rect 377930 586294 377998 586350
rect 378054 586294 378122 586350
rect 378178 586294 378246 586350
rect 378302 586294 408594 586350
rect 408650 586294 408718 586350
rect 408774 586294 408842 586350
rect 408898 586294 408966 586350
rect 409022 586294 439314 586350
rect 439370 586294 439438 586350
rect 439494 586294 439562 586350
rect 439618 586294 439686 586350
rect 439742 586294 470034 586350
rect 470090 586294 470158 586350
rect 470214 586294 470282 586350
rect 470338 586294 470406 586350
rect 470462 586294 500754 586350
rect 500810 586294 500878 586350
rect 500934 586294 501002 586350
rect 501058 586294 501126 586350
rect 501182 586294 531474 586350
rect 531530 586294 531598 586350
rect 531654 586294 531722 586350
rect 531778 586294 531846 586350
rect 531902 586294 562194 586350
rect 562250 586294 562318 586350
rect 562374 586294 562442 586350
rect 562498 586294 562566 586350
rect 562622 586294 592914 586350
rect 592970 586294 593038 586350
rect 593094 586294 593162 586350
rect 593218 586294 593286 586350
rect 593342 586294 597456 586350
rect 597512 586294 597580 586350
rect 597636 586294 597704 586350
rect 597760 586294 597828 586350
rect 597884 586294 597980 586350
rect -1916 586226 597980 586294
rect -1916 586170 -1820 586226
rect -1764 586170 -1696 586226
rect -1640 586170 -1572 586226
rect -1516 586170 -1448 586226
rect -1392 586170 9234 586226
rect 9290 586170 9358 586226
rect 9414 586170 9482 586226
rect 9538 586170 9606 586226
rect 9662 586170 39954 586226
rect 40010 586170 40078 586226
rect 40134 586170 40202 586226
rect 40258 586170 40326 586226
rect 40382 586170 70674 586226
rect 70730 586170 70798 586226
rect 70854 586170 70922 586226
rect 70978 586170 71046 586226
rect 71102 586170 101394 586226
rect 101450 586170 101518 586226
rect 101574 586170 101642 586226
rect 101698 586170 101766 586226
rect 101822 586170 132114 586226
rect 132170 586170 132238 586226
rect 132294 586170 132362 586226
rect 132418 586170 132486 586226
rect 132542 586170 162834 586226
rect 162890 586170 162958 586226
rect 163014 586170 163082 586226
rect 163138 586170 163206 586226
rect 163262 586170 193554 586226
rect 193610 586170 193678 586226
rect 193734 586170 193802 586226
rect 193858 586170 193926 586226
rect 193982 586170 224274 586226
rect 224330 586170 224398 586226
rect 224454 586170 224522 586226
rect 224578 586170 224646 586226
rect 224702 586170 254994 586226
rect 255050 586170 255118 586226
rect 255174 586170 255242 586226
rect 255298 586170 255366 586226
rect 255422 586170 285714 586226
rect 285770 586170 285838 586226
rect 285894 586170 285962 586226
rect 286018 586170 286086 586226
rect 286142 586170 316434 586226
rect 316490 586170 316558 586226
rect 316614 586170 316682 586226
rect 316738 586170 316806 586226
rect 316862 586170 347154 586226
rect 347210 586170 347278 586226
rect 347334 586170 347402 586226
rect 347458 586170 347526 586226
rect 347582 586170 377874 586226
rect 377930 586170 377998 586226
rect 378054 586170 378122 586226
rect 378178 586170 378246 586226
rect 378302 586170 408594 586226
rect 408650 586170 408718 586226
rect 408774 586170 408842 586226
rect 408898 586170 408966 586226
rect 409022 586170 439314 586226
rect 439370 586170 439438 586226
rect 439494 586170 439562 586226
rect 439618 586170 439686 586226
rect 439742 586170 470034 586226
rect 470090 586170 470158 586226
rect 470214 586170 470282 586226
rect 470338 586170 470406 586226
rect 470462 586170 500754 586226
rect 500810 586170 500878 586226
rect 500934 586170 501002 586226
rect 501058 586170 501126 586226
rect 501182 586170 531474 586226
rect 531530 586170 531598 586226
rect 531654 586170 531722 586226
rect 531778 586170 531846 586226
rect 531902 586170 562194 586226
rect 562250 586170 562318 586226
rect 562374 586170 562442 586226
rect 562498 586170 562566 586226
rect 562622 586170 592914 586226
rect 592970 586170 593038 586226
rect 593094 586170 593162 586226
rect 593218 586170 593286 586226
rect 593342 586170 597456 586226
rect 597512 586170 597580 586226
rect 597636 586170 597704 586226
rect 597760 586170 597828 586226
rect 597884 586170 597980 586226
rect -1916 586102 597980 586170
rect -1916 586046 -1820 586102
rect -1764 586046 -1696 586102
rect -1640 586046 -1572 586102
rect -1516 586046 -1448 586102
rect -1392 586046 9234 586102
rect 9290 586046 9358 586102
rect 9414 586046 9482 586102
rect 9538 586046 9606 586102
rect 9662 586046 39954 586102
rect 40010 586046 40078 586102
rect 40134 586046 40202 586102
rect 40258 586046 40326 586102
rect 40382 586046 70674 586102
rect 70730 586046 70798 586102
rect 70854 586046 70922 586102
rect 70978 586046 71046 586102
rect 71102 586046 101394 586102
rect 101450 586046 101518 586102
rect 101574 586046 101642 586102
rect 101698 586046 101766 586102
rect 101822 586046 132114 586102
rect 132170 586046 132238 586102
rect 132294 586046 132362 586102
rect 132418 586046 132486 586102
rect 132542 586046 162834 586102
rect 162890 586046 162958 586102
rect 163014 586046 163082 586102
rect 163138 586046 163206 586102
rect 163262 586046 193554 586102
rect 193610 586046 193678 586102
rect 193734 586046 193802 586102
rect 193858 586046 193926 586102
rect 193982 586046 224274 586102
rect 224330 586046 224398 586102
rect 224454 586046 224522 586102
rect 224578 586046 224646 586102
rect 224702 586046 254994 586102
rect 255050 586046 255118 586102
rect 255174 586046 255242 586102
rect 255298 586046 255366 586102
rect 255422 586046 285714 586102
rect 285770 586046 285838 586102
rect 285894 586046 285962 586102
rect 286018 586046 286086 586102
rect 286142 586046 316434 586102
rect 316490 586046 316558 586102
rect 316614 586046 316682 586102
rect 316738 586046 316806 586102
rect 316862 586046 347154 586102
rect 347210 586046 347278 586102
rect 347334 586046 347402 586102
rect 347458 586046 347526 586102
rect 347582 586046 377874 586102
rect 377930 586046 377998 586102
rect 378054 586046 378122 586102
rect 378178 586046 378246 586102
rect 378302 586046 408594 586102
rect 408650 586046 408718 586102
rect 408774 586046 408842 586102
rect 408898 586046 408966 586102
rect 409022 586046 439314 586102
rect 439370 586046 439438 586102
rect 439494 586046 439562 586102
rect 439618 586046 439686 586102
rect 439742 586046 470034 586102
rect 470090 586046 470158 586102
rect 470214 586046 470282 586102
rect 470338 586046 470406 586102
rect 470462 586046 500754 586102
rect 500810 586046 500878 586102
rect 500934 586046 501002 586102
rect 501058 586046 501126 586102
rect 501182 586046 531474 586102
rect 531530 586046 531598 586102
rect 531654 586046 531722 586102
rect 531778 586046 531846 586102
rect 531902 586046 562194 586102
rect 562250 586046 562318 586102
rect 562374 586046 562442 586102
rect 562498 586046 562566 586102
rect 562622 586046 592914 586102
rect 592970 586046 593038 586102
rect 593094 586046 593162 586102
rect 593218 586046 593286 586102
rect 593342 586046 597456 586102
rect 597512 586046 597580 586102
rect 597636 586046 597704 586102
rect 597760 586046 597828 586102
rect 597884 586046 597980 586102
rect -1916 585978 597980 586046
rect -1916 585922 -1820 585978
rect -1764 585922 -1696 585978
rect -1640 585922 -1572 585978
rect -1516 585922 -1448 585978
rect -1392 585922 9234 585978
rect 9290 585922 9358 585978
rect 9414 585922 9482 585978
rect 9538 585922 9606 585978
rect 9662 585922 39954 585978
rect 40010 585922 40078 585978
rect 40134 585922 40202 585978
rect 40258 585922 40326 585978
rect 40382 585922 70674 585978
rect 70730 585922 70798 585978
rect 70854 585922 70922 585978
rect 70978 585922 71046 585978
rect 71102 585922 101394 585978
rect 101450 585922 101518 585978
rect 101574 585922 101642 585978
rect 101698 585922 101766 585978
rect 101822 585922 132114 585978
rect 132170 585922 132238 585978
rect 132294 585922 132362 585978
rect 132418 585922 132486 585978
rect 132542 585922 162834 585978
rect 162890 585922 162958 585978
rect 163014 585922 163082 585978
rect 163138 585922 163206 585978
rect 163262 585922 193554 585978
rect 193610 585922 193678 585978
rect 193734 585922 193802 585978
rect 193858 585922 193926 585978
rect 193982 585922 224274 585978
rect 224330 585922 224398 585978
rect 224454 585922 224522 585978
rect 224578 585922 224646 585978
rect 224702 585922 254994 585978
rect 255050 585922 255118 585978
rect 255174 585922 255242 585978
rect 255298 585922 255366 585978
rect 255422 585922 285714 585978
rect 285770 585922 285838 585978
rect 285894 585922 285962 585978
rect 286018 585922 286086 585978
rect 286142 585922 316434 585978
rect 316490 585922 316558 585978
rect 316614 585922 316682 585978
rect 316738 585922 316806 585978
rect 316862 585922 347154 585978
rect 347210 585922 347278 585978
rect 347334 585922 347402 585978
rect 347458 585922 347526 585978
rect 347582 585922 377874 585978
rect 377930 585922 377998 585978
rect 378054 585922 378122 585978
rect 378178 585922 378246 585978
rect 378302 585922 408594 585978
rect 408650 585922 408718 585978
rect 408774 585922 408842 585978
rect 408898 585922 408966 585978
rect 409022 585922 439314 585978
rect 439370 585922 439438 585978
rect 439494 585922 439562 585978
rect 439618 585922 439686 585978
rect 439742 585922 470034 585978
rect 470090 585922 470158 585978
rect 470214 585922 470282 585978
rect 470338 585922 470406 585978
rect 470462 585922 500754 585978
rect 500810 585922 500878 585978
rect 500934 585922 501002 585978
rect 501058 585922 501126 585978
rect 501182 585922 531474 585978
rect 531530 585922 531598 585978
rect 531654 585922 531722 585978
rect 531778 585922 531846 585978
rect 531902 585922 562194 585978
rect 562250 585922 562318 585978
rect 562374 585922 562442 585978
rect 562498 585922 562566 585978
rect 562622 585922 592914 585978
rect 592970 585922 593038 585978
rect 593094 585922 593162 585978
rect 593218 585922 593286 585978
rect 593342 585922 597456 585978
rect 597512 585922 597580 585978
rect 597636 585922 597704 585978
rect 597760 585922 597828 585978
rect 597884 585922 597980 585978
rect -1916 585826 597980 585922
rect -1916 580350 597980 580446
rect -1916 580294 -860 580350
rect -804 580294 -736 580350
rect -680 580294 -612 580350
rect -556 580294 -488 580350
rect -432 580294 5514 580350
rect 5570 580294 5638 580350
rect 5694 580294 5762 580350
rect 5818 580294 5886 580350
rect 5942 580294 36234 580350
rect 36290 580294 36358 580350
rect 36414 580294 36482 580350
rect 36538 580294 36606 580350
rect 36662 580294 66954 580350
rect 67010 580294 67078 580350
rect 67134 580294 67202 580350
rect 67258 580294 67326 580350
rect 67382 580294 97674 580350
rect 97730 580294 97798 580350
rect 97854 580294 97922 580350
rect 97978 580294 98046 580350
rect 98102 580294 128394 580350
rect 128450 580294 128518 580350
rect 128574 580294 128642 580350
rect 128698 580294 128766 580350
rect 128822 580294 159114 580350
rect 159170 580294 159238 580350
rect 159294 580294 159362 580350
rect 159418 580294 159486 580350
rect 159542 580294 189834 580350
rect 189890 580294 189958 580350
rect 190014 580294 190082 580350
rect 190138 580294 190206 580350
rect 190262 580294 220554 580350
rect 220610 580294 220678 580350
rect 220734 580294 220802 580350
rect 220858 580294 220926 580350
rect 220982 580294 251274 580350
rect 251330 580294 251398 580350
rect 251454 580294 251522 580350
rect 251578 580294 251646 580350
rect 251702 580294 281994 580350
rect 282050 580294 282118 580350
rect 282174 580294 282242 580350
rect 282298 580294 282366 580350
rect 282422 580294 312714 580350
rect 312770 580294 312838 580350
rect 312894 580294 312962 580350
rect 313018 580294 313086 580350
rect 313142 580294 343434 580350
rect 343490 580294 343558 580350
rect 343614 580294 343682 580350
rect 343738 580294 343806 580350
rect 343862 580294 374154 580350
rect 374210 580294 374278 580350
rect 374334 580294 374402 580350
rect 374458 580294 374526 580350
rect 374582 580294 404874 580350
rect 404930 580294 404998 580350
rect 405054 580294 405122 580350
rect 405178 580294 405246 580350
rect 405302 580294 435594 580350
rect 435650 580294 435718 580350
rect 435774 580294 435842 580350
rect 435898 580294 435966 580350
rect 436022 580294 466314 580350
rect 466370 580294 466438 580350
rect 466494 580294 466562 580350
rect 466618 580294 466686 580350
rect 466742 580294 497034 580350
rect 497090 580294 497158 580350
rect 497214 580294 497282 580350
rect 497338 580294 497406 580350
rect 497462 580294 527754 580350
rect 527810 580294 527878 580350
rect 527934 580294 528002 580350
rect 528058 580294 528126 580350
rect 528182 580294 558474 580350
rect 558530 580294 558598 580350
rect 558654 580294 558722 580350
rect 558778 580294 558846 580350
rect 558902 580294 589194 580350
rect 589250 580294 589318 580350
rect 589374 580294 589442 580350
rect 589498 580294 589566 580350
rect 589622 580294 596496 580350
rect 596552 580294 596620 580350
rect 596676 580294 596744 580350
rect 596800 580294 596868 580350
rect 596924 580294 597980 580350
rect -1916 580226 597980 580294
rect -1916 580170 -860 580226
rect -804 580170 -736 580226
rect -680 580170 -612 580226
rect -556 580170 -488 580226
rect -432 580170 5514 580226
rect 5570 580170 5638 580226
rect 5694 580170 5762 580226
rect 5818 580170 5886 580226
rect 5942 580170 36234 580226
rect 36290 580170 36358 580226
rect 36414 580170 36482 580226
rect 36538 580170 36606 580226
rect 36662 580170 66954 580226
rect 67010 580170 67078 580226
rect 67134 580170 67202 580226
rect 67258 580170 67326 580226
rect 67382 580170 97674 580226
rect 97730 580170 97798 580226
rect 97854 580170 97922 580226
rect 97978 580170 98046 580226
rect 98102 580170 128394 580226
rect 128450 580170 128518 580226
rect 128574 580170 128642 580226
rect 128698 580170 128766 580226
rect 128822 580170 159114 580226
rect 159170 580170 159238 580226
rect 159294 580170 159362 580226
rect 159418 580170 159486 580226
rect 159542 580170 189834 580226
rect 189890 580170 189958 580226
rect 190014 580170 190082 580226
rect 190138 580170 190206 580226
rect 190262 580170 220554 580226
rect 220610 580170 220678 580226
rect 220734 580170 220802 580226
rect 220858 580170 220926 580226
rect 220982 580170 251274 580226
rect 251330 580170 251398 580226
rect 251454 580170 251522 580226
rect 251578 580170 251646 580226
rect 251702 580170 281994 580226
rect 282050 580170 282118 580226
rect 282174 580170 282242 580226
rect 282298 580170 282366 580226
rect 282422 580170 312714 580226
rect 312770 580170 312838 580226
rect 312894 580170 312962 580226
rect 313018 580170 313086 580226
rect 313142 580170 343434 580226
rect 343490 580170 343558 580226
rect 343614 580170 343682 580226
rect 343738 580170 343806 580226
rect 343862 580170 374154 580226
rect 374210 580170 374278 580226
rect 374334 580170 374402 580226
rect 374458 580170 374526 580226
rect 374582 580170 404874 580226
rect 404930 580170 404998 580226
rect 405054 580170 405122 580226
rect 405178 580170 405246 580226
rect 405302 580170 435594 580226
rect 435650 580170 435718 580226
rect 435774 580170 435842 580226
rect 435898 580170 435966 580226
rect 436022 580170 466314 580226
rect 466370 580170 466438 580226
rect 466494 580170 466562 580226
rect 466618 580170 466686 580226
rect 466742 580170 497034 580226
rect 497090 580170 497158 580226
rect 497214 580170 497282 580226
rect 497338 580170 497406 580226
rect 497462 580170 527754 580226
rect 527810 580170 527878 580226
rect 527934 580170 528002 580226
rect 528058 580170 528126 580226
rect 528182 580170 558474 580226
rect 558530 580170 558598 580226
rect 558654 580170 558722 580226
rect 558778 580170 558846 580226
rect 558902 580170 589194 580226
rect 589250 580170 589318 580226
rect 589374 580170 589442 580226
rect 589498 580170 589566 580226
rect 589622 580170 596496 580226
rect 596552 580170 596620 580226
rect 596676 580170 596744 580226
rect 596800 580170 596868 580226
rect 596924 580170 597980 580226
rect -1916 580102 597980 580170
rect -1916 580046 -860 580102
rect -804 580046 -736 580102
rect -680 580046 -612 580102
rect -556 580046 -488 580102
rect -432 580046 5514 580102
rect 5570 580046 5638 580102
rect 5694 580046 5762 580102
rect 5818 580046 5886 580102
rect 5942 580046 36234 580102
rect 36290 580046 36358 580102
rect 36414 580046 36482 580102
rect 36538 580046 36606 580102
rect 36662 580046 66954 580102
rect 67010 580046 67078 580102
rect 67134 580046 67202 580102
rect 67258 580046 67326 580102
rect 67382 580046 97674 580102
rect 97730 580046 97798 580102
rect 97854 580046 97922 580102
rect 97978 580046 98046 580102
rect 98102 580046 128394 580102
rect 128450 580046 128518 580102
rect 128574 580046 128642 580102
rect 128698 580046 128766 580102
rect 128822 580046 159114 580102
rect 159170 580046 159238 580102
rect 159294 580046 159362 580102
rect 159418 580046 159486 580102
rect 159542 580046 189834 580102
rect 189890 580046 189958 580102
rect 190014 580046 190082 580102
rect 190138 580046 190206 580102
rect 190262 580046 220554 580102
rect 220610 580046 220678 580102
rect 220734 580046 220802 580102
rect 220858 580046 220926 580102
rect 220982 580046 251274 580102
rect 251330 580046 251398 580102
rect 251454 580046 251522 580102
rect 251578 580046 251646 580102
rect 251702 580046 281994 580102
rect 282050 580046 282118 580102
rect 282174 580046 282242 580102
rect 282298 580046 282366 580102
rect 282422 580046 312714 580102
rect 312770 580046 312838 580102
rect 312894 580046 312962 580102
rect 313018 580046 313086 580102
rect 313142 580046 343434 580102
rect 343490 580046 343558 580102
rect 343614 580046 343682 580102
rect 343738 580046 343806 580102
rect 343862 580046 374154 580102
rect 374210 580046 374278 580102
rect 374334 580046 374402 580102
rect 374458 580046 374526 580102
rect 374582 580046 404874 580102
rect 404930 580046 404998 580102
rect 405054 580046 405122 580102
rect 405178 580046 405246 580102
rect 405302 580046 435594 580102
rect 435650 580046 435718 580102
rect 435774 580046 435842 580102
rect 435898 580046 435966 580102
rect 436022 580046 466314 580102
rect 466370 580046 466438 580102
rect 466494 580046 466562 580102
rect 466618 580046 466686 580102
rect 466742 580046 497034 580102
rect 497090 580046 497158 580102
rect 497214 580046 497282 580102
rect 497338 580046 497406 580102
rect 497462 580046 527754 580102
rect 527810 580046 527878 580102
rect 527934 580046 528002 580102
rect 528058 580046 528126 580102
rect 528182 580046 558474 580102
rect 558530 580046 558598 580102
rect 558654 580046 558722 580102
rect 558778 580046 558846 580102
rect 558902 580046 589194 580102
rect 589250 580046 589318 580102
rect 589374 580046 589442 580102
rect 589498 580046 589566 580102
rect 589622 580046 596496 580102
rect 596552 580046 596620 580102
rect 596676 580046 596744 580102
rect 596800 580046 596868 580102
rect 596924 580046 597980 580102
rect -1916 579978 597980 580046
rect -1916 579922 -860 579978
rect -804 579922 -736 579978
rect -680 579922 -612 579978
rect -556 579922 -488 579978
rect -432 579922 5514 579978
rect 5570 579922 5638 579978
rect 5694 579922 5762 579978
rect 5818 579922 5886 579978
rect 5942 579922 36234 579978
rect 36290 579922 36358 579978
rect 36414 579922 36482 579978
rect 36538 579922 36606 579978
rect 36662 579922 66954 579978
rect 67010 579922 67078 579978
rect 67134 579922 67202 579978
rect 67258 579922 67326 579978
rect 67382 579922 97674 579978
rect 97730 579922 97798 579978
rect 97854 579922 97922 579978
rect 97978 579922 98046 579978
rect 98102 579922 128394 579978
rect 128450 579922 128518 579978
rect 128574 579922 128642 579978
rect 128698 579922 128766 579978
rect 128822 579922 159114 579978
rect 159170 579922 159238 579978
rect 159294 579922 159362 579978
rect 159418 579922 159486 579978
rect 159542 579922 189834 579978
rect 189890 579922 189958 579978
rect 190014 579922 190082 579978
rect 190138 579922 190206 579978
rect 190262 579922 220554 579978
rect 220610 579922 220678 579978
rect 220734 579922 220802 579978
rect 220858 579922 220926 579978
rect 220982 579922 251274 579978
rect 251330 579922 251398 579978
rect 251454 579922 251522 579978
rect 251578 579922 251646 579978
rect 251702 579922 281994 579978
rect 282050 579922 282118 579978
rect 282174 579922 282242 579978
rect 282298 579922 282366 579978
rect 282422 579922 312714 579978
rect 312770 579922 312838 579978
rect 312894 579922 312962 579978
rect 313018 579922 313086 579978
rect 313142 579922 343434 579978
rect 343490 579922 343558 579978
rect 343614 579922 343682 579978
rect 343738 579922 343806 579978
rect 343862 579922 374154 579978
rect 374210 579922 374278 579978
rect 374334 579922 374402 579978
rect 374458 579922 374526 579978
rect 374582 579922 404874 579978
rect 404930 579922 404998 579978
rect 405054 579922 405122 579978
rect 405178 579922 405246 579978
rect 405302 579922 435594 579978
rect 435650 579922 435718 579978
rect 435774 579922 435842 579978
rect 435898 579922 435966 579978
rect 436022 579922 466314 579978
rect 466370 579922 466438 579978
rect 466494 579922 466562 579978
rect 466618 579922 466686 579978
rect 466742 579922 497034 579978
rect 497090 579922 497158 579978
rect 497214 579922 497282 579978
rect 497338 579922 497406 579978
rect 497462 579922 527754 579978
rect 527810 579922 527878 579978
rect 527934 579922 528002 579978
rect 528058 579922 528126 579978
rect 528182 579922 558474 579978
rect 558530 579922 558598 579978
rect 558654 579922 558722 579978
rect 558778 579922 558846 579978
rect 558902 579922 589194 579978
rect 589250 579922 589318 579978
rect 589374 579922 589442 579978
rect 589498 579922 589566 579978
rect 589622 579922 596496 579978
rect 596552 579922 596620 579978
rect 596676 579922 596744 579978
rect 596800 579922 596868 579978
rect 596924 579922 597980 579978
rect -1916 579826 597980 579922
rect -1916 568350 597980 568446
rect -1916 568294 -1820 568350
rect -1764 568294 -1696 568350
rect -1640 568294 -1572 568350
rect -1516 568294 -1448 568350
rect -1392 568294 9234 568350
rect 9290 568294 9358 568350
rect 9414 568294 9482 568350
rect 9538 568294 9606 568350
rect 9662 568294 39954 568350
rect 40010 568294 40078 568350
rect 40134 568294 40202 568350
rect 40258 568294 40326 568350
rect 40382 568294 70674 568350
rect 70730 568294 70798 568350
rect 70854 568294 70922 568350
rect 70978 568294 71046 568350
rect 71102 568294 101394 568350
rect 101450 568294 101518 568350
rect 101574 568294 101642 568350
rect 101698 568294 101766 568350
rect 101822 568294 132114 568350
rect 132170 568294 132238 568350
rect 132294 568294 132362 568350
rect 132418 568294 132486 568350
rect 132542 568294 162834 568350
rect 162890 568294 162958 568350
rect 163014 568294 163082 568350
rect 163138 568294 163206 568350
rect 163262 568294 193554 568350
rect 193610 568294 193678 568350
rect 193734 568294 193802 568350
rect 193858 568294 193926 568350
rect 193982 568294 224274 568350
rect 224330 568294 224398 568350
rect 224454 568294 224522 568350
rect 224578 568294 224646 568350
rect 224702 568294 254994 568350
rect 255050 568294 255118 568350
rect 255174 568294 255242 568350
rect 255298 568294 255366 568350
rect 255422 568294 285714 568350
rect 285770 568294 285838 568350
rect 285894 568294 285962 568350
rect 286018 568294 286086 568350
rect 286142 568294 316434 568350
rect 316490 568294 316558 568350
rect 316614 568294 316682 568350
rect 316738 568294 316806 568350
rect 316862 568294 347154 568350
rect 347210 568294 347278 568350
rect 347334 568294 347402 568350
rect 347458 568294 347526 568350
rect 347582 568294 377874 568350
rect 377930 568294 377998 568350
rect 378054 568294 378122 568350
rect 378178 568294 378246 568350
rect 378302 568294 408594 568350
rect 408650 568294 408718 568350
rect 408774 568294 408842 568350
rect 408898 568294 408966 568350
rect 409022 568294 439314 568350
rect 439370 568294 439438 568350
rect 439494 568294 439562 568350
rect 439618 568294 439686 568350
rect 439742 568294 470034 568350
rect 470090 568294 470158 568350
rect 470214 568294 470282 568350
rect 470338 568294 470406 568350
rect 470462 568294 500754 568350
rect 500810 568294 500878 568350
rect 500934 568294 501002 568350
rect 501058 568294 501126 568350
rect 501182 568294 531474 568350
rect 531530 568294 531598 568350
rect 531654 568294 531722 568350
rect 531778 568294 531846 568350
rect 531902 568294 562194 568350
rect 562250 568294 562318 568350
rect 562374 568294 562442 568350
rect 562498 568294 562566 568350
rect 562622 568294 592914 568350
rect 592970 568294 593038 568350
rect 593094 568294 593162 568350
rect 593218 568294 593286 568350
rect 593342 568294 597456 568350
rect 597512 568294 597580 568350
rect 597636 568294 597704 568350
rect 597760 568294 597828 568350
rect 597884 568294 597980 568350
rect -1916 568226 597980 568294
rect -1916 568170 -1820 568226
rect -1764 568170 -1696 568226
rect -1640 568170 -1572 568226
rect -1516 568170 -1448 568226
rect -1392 568170 9234 568226
rect 9290 568170 9358 568226
rect 9414 568170 9482 568226
rect 9538 568170 9606 568226
rect 9662 568170 39954 568226
rect 40010 568170 40078 568226
rect 40134 568170 40202 568226
rect 40258 568170 40326 568226
rect 40382 568170 70674 568226
rect 70730 568170 70798 568226
rect 70854 568170 70922 568226
rect 70978 568170 71046 568226
rect 71102 568170 101394 568226
rect 101450 568170 101518 568226
rect 101574 568170 101642 568226
rect 101698 568170 101766 568226
rect 101822 568170 132114 568226
rect 132170 568170 132238 568226
rect 132294 568170 132362 568226
rect 132418 568170 132486 568226
rect 132542 568170 162834 568226
rect 162890 568170 162958 568226
rect 163014 568170 163082 568226
rect 163138 568170 163206 568226
rect 163262 568170 193554 568226
rect 193610 568170 193678 568226
rect 193734 568170 193802 568226
rect 193858 568170 193926 568226
rect 193982 568170 224274 568226
rect 224330 568170 224398 568226
rect 224454 568170 224522 568226
rect 224578 568170 224646 568226
rect 224702 568170 254994 568226
rect 255050 568170 255118 568226
rect 255174 568170 255242 568226
rect 255298 568170 255366 568226
rect 255422 568170 285714 568226
rect 285770 568170 285838 568226
rect 285894 568170 285962 568226
rect 286018 568170 286086 568226
rect 286142 568170 316434 568226
rect 316490 568170 316558 568226
rect 316614 568170 316682 568226
rect 316738 568170 316806 568226
rect 316862 568170 347154 568226
rect 347210 568170 347278 568226
rect 347334 568170 347402 568226
rect 347458 568170 347526 568226
rect 347582 568170 377874 568226
rect 377930 568170 377998 568226
rect 378054 568170 378122 568226
rect 378178 568170 378246 568226
rect 378302 568170 408594 568226
rect 408650 568170 408718 568226
rect 408774 568170 408842 568226
rect 408898 568170 408966 568226
rect 409022 568170 439314 568226
rect 439370 568170 439438 568226
rect 439494 568170 439562 568226
rect 439618 568170 439686 568226
rect 439742 568170 470034 568226
rect 470090 568170 470158 568226
rect 470214 568170 470282 568226
rect 470338 568170 470406 568226
rect 470462 568170 500754 568226
rect 500810 568170 500878 568226
rect 500934 568170 501002 568226
rect 501058 568170 501126 568226
rect 501182 568170 531474 568226
rect 531530 568170 531598 568226
rect 531654 568170 531722 568226
rect 531778 568170 531846 568226
rect 531902 568170 562194 568226
rect 562250 568170 562318 568226
rect 562374 568170 562442 568226
rect 562498 568170 562566 568226
rect 562622 568170 592914 568226
rect 592970 568170 593038 568226
rect 593094 568170 593162 568226
rect 593218 568170 593286 568226
rect 593342 568170 597456 568226
rect 597512 568170 597580 568226
rect 597636 568170 597704 568226
rect 597760 568170 597828 568226
rect 597884 568170 597980 568226
rect -1916 568102 597980 568170
rect -1916 568046 -1820 568102
rect -1764 568046 -1696 568102
rect -1640 568046 -1572 568102
rect -1516 568046 -1448 568102
rect -1392 568046 9234 568102
rect 9290 568046 9358 568102
rect 9414 568046 9482 568102
rect 9538 568046 9606 568102
rect 9662 568046 39954 568102
rect 40010 568046 40078 568102
rect 40134 568046 40202 568102
rect 40258 568046 40326 568102
rect 40382 568046 70674 568102
rect 70730 568046 70798 568102
rect 70854 568046 70922 568102
rect 70978 568046 71046 568102
rect 71102 568046 101394 568102
rect 101450 568046 101518 568102
rect 101574 568046 101642 568102
rect 101698 568046 101766 568102
rect 101822 568046 132114 568102
rect 132170 568046 132238 568102
rect 132294 568046 132362 568102
rect 132418 568046 132486 568102
rect 132542 568046 162834 568102
rect 162890 568046 162958 568102
rect 163014 568046 163082 568102
rect 163138 568046 163206 568102
rect 163262 568046 193554 568102
rect 193610 568046 193678 568102
rect 193734 568046 193802 568102
rect 193858 568046 193926 568102
rect 193982 568046 224274 568102
rect 224330 568046 224398 568102
rect 224454 568046 224522 568102
rect 224578 568046 224646 568102
rect 224702 568046 254994 568102
rect 255050 568046 255118 568102
rect 255174 568046 255242 568102
rect 255298 568046 255366 568102
rect 255422 568046 285714 568102
rect 285770 568046 285838 568102
rect 285894 568046 285962 568102
rect 286018 568046 286086 568102
rect 286142 568046 316434 568102
rect 316490 568046 316558 568102
rect 316614 568046 316682 568102
rect 316738 568046 316806 568102
rect 316862 568046 347154 568102
rect 347210 568046 347278 568102
rect 347334 568046 347402 568102
rect 347458 568046 347526 568102
rect 347582 568046 377874 568102
rect 377930 568046 377998 568102
rect 378054 568046 378122 568102
rect 378178 568046 378246 568102
rect 378302 568046 408594 568102
rect 408650 568046 408718 568102
rect 408774 568046 408842 568102
rect 408898 568046 408966 568102
rect 409022 568046 439314 568102
rect 439370 568046 439438 568102
rect 439494 568046 439562 568102
rect 439618 568046 439686 568102
rect 439742 568046 470034 568102
rect 470090 568046 470158 568102
rect 470214 568046 470282 568102
rect 470338 568046 470406 568102
rect 470462 568046 500754 568102
rect 500810 568046 500878 568102
rect 500934 568046 501002 568102
rect 501058 568046 501126 568102
rect 501182 568046 531474 568102
rect 531530 568046 531598 568102
rect 531654 568046 531722 568102
rect 531778 568046 531846 568102
rect 531902 568046 562194 568102
rect 562250 568046 562318 568102
rect 562374 568046 562442 568102
rect 562498 568046 562566 568102
rect 562622 568046 592914 568102
rect 592970 568046 593038 568102
rect 593094 568046 593162 568102
rect 593218 568046 593286 568102
rect 593342 568046 597456 568102
rect 597512 568046 597580 568102
rect 597636 568046 597704 568102
rect 597760 568046 597828 568102
rect 597884 568046 597980 568102
rect -1916 567978 597980 568046
rect -1916 567922 -1820 567978
rect -1764 567922 -1696 567978
rect -1640 567922 -1572 567978
rect -1516 567922 -1448 567978
rect -1392 567922 9234 567978
rect 9290 567922 9358 567978
rect 9414 567922 9482 567978
rect 9538 567922 9606 567978
rect 9662 567922 39954 567978
rect 40010 567922 40078 567978
rect 40134 567922 40202 567978
rect 40258 567922 40326 567978
rect 40382 567922 70674 567978
rect 70730 567922 70798 567978
rect 70854 567922 70922 567978
rect 70978 567922 71046 567978
rect 71102 567922 101394 567978
rect 101450 567922 101518 567978
rect 101574 567922 101642 567978
rect 101698 567922 101766 567978
rect 101822 567922 132114 567978
rect 132170 567922 132238 567978
rect 132294 567922 132362 567978
rect 132418 567922 132486 567978
rect 132542 567922 162834 567978
rect 162890 567922 162958 567978
rect 163014 567922 163082 567978
rect 163138 567922 163206 567978
rect 163262 567922 193554 567978
rect 193610 567922 193678 567978
rect 193734 567922 193802 567978
rect 193858 567922 193926 567978
rect 193982 567922 224274 567978
rect 224330 567922 224398 567978
rect 224454 567922 224522 567978
rect 224578 567922 224646 567978
rect 224702 567922 254994 567978
rect 255050 567922 255118 567978
rect 255174 567922 255242 567978
rect 255298 567922 255366 567978
rect 255422 567922 285714 567978
rect 285770 567922 285838 567978
rect 285894 567922 285962 567978
rect 286018 567922 286086 567978
rect 286142 567922 316434 567978
rect 316490 567922 316558 567978
rect 316614 567922 316682 567978
rect 316738 567922 316806 567978
rect 316862 567922 347154 567978
rect 347210 567922 347278 567978
rect 347334 567922 347402 567978
rect 347458 567922 347526 567978
rect 347582 567922 377874 567978
rect 377930 567922 377998 567978
rect 378054 567922 378122 567978
rect 378178 567922 378246 567978
rect 378302 567922 408594 567978
rect 408650 567922 408718 567978
rect 408774 567922 408842 567978
rect 408898 567922 408966 567978
rect 409022 567922 439314 567978
rect 439370 567922 439438 567978
rect 439494 567922 439562 567978
rect 439618 567922 439686 567978
rect 439742 567922 470034 567978
rect 470090 567922 470158 567978
rect 470214 567922 470282 567978
rect 470338 567922 470406 567978
rect 470462 567922 500754 567978
rect 500810 567922 500878 567978
rect 500934 567922 501002 567978
rect 501058 567922 501126 567978
rect 501182 567922 531474 567978
rect 531530 567922 531598 567978
rect 531654 567922 531722 567978
rect 531778 567922 531846 567978
rect 531902 567922 562194 567978
rect 562250 567922 562318 567978
rect 562374 567922 562442 567978
rect 562498 567922 562566 567978
rect 562622 567922 592914 567978
rect 592970 567922 593038 567978
rect 593094 567922 593162 567978
rect 593218 567922 593286 567978
rect 593342 567922 597456 567978
rect 597512 567922 597580 567978
rect 597636 567922 597704 567978
rect 597760 567922 597828 567978
rect 597884 567922 597980 567978
rect -1916 567826 597980 567922
rect -1916 562350 597980 562446
rect -1916 562294 -860 562350
rect -804 562294 -736 562350
rect -680 562294 -612 562350
rect -556 562294 -488 562350
rect -432 562294 5514 562350
rect 5570 562294 5638 562350
rect 5694 562294 5762 562350
rect 5818 562294 5886 562350
rect 5942 562294 36234 562350
rect 36290 562294 36358 562350
rect 36414 562294 36482 562350
rect 36538 562294 36606 562350
rect 36662 562294 66954 562350
rect 67010 562294 67078 562350
rect 67134 562294 67202 562350
rect 67258 562294 67326 562350
rect 67382 562294 97674 562350
rect 97730 562294 97798 562350
rect 97854 562294 97922 562350
rect 97978 562294 98046 562350
rect 98102 562294 128394 562350
rect 128450 562294 128518 562350
rect 128574 562294 128642 562350
rect 128698 562294 128766 562350
rect 128822 562294 159114 562350
rect 159170 562294 159238 562350
rect 159294 562294 159362 562350
rect 159418 562294 159486 562350
rect 159542 562294 189834 562350
rect 189890 562294 189958 562350
rect 190014 562294 190082 562350
rect 190138 562294 190206 562350
rect 190262 562294 220554 562350
rect 220610 562294 220678 562350
rect 220734 562294 220802 562350
rect 220858 562294 220926 562350
rect 220982 562294 251274 562350
rect 251330 562294 251398 562350
rect 251454 562294 251522 562350
rect 251578 562294 251646 562350
rect 251702 562294 281994 562350
rect 282050 562294 282118 562350
rect 282174 562294 282242 562350
rect 282298 562294 282366 562350
rect 282422 562294 312714 562350
rect 312770 562294 312838 562350
rect 312894 562294 312962 562350
rect 313018 562294 313086 562350
rect 313142 562294 343434 562350
rect 343490 562294 343558 562350
rect 343614 562294 343682 562350
rect 343738 562294 343806 562350
rect 343862 562294 374154 562350
rect 374210 562294 374278 562350
rect 374334 562294 374402 562350
rect 374458 562294 374526 562350
rect 374582 562294 404874 562350
rect 404930 562294 404998 562350
rect 405054 562294 405122 562350
rect 405178 562294 405246 562350
rect 405302 562294 435594 562350
rect 435650 562294 435718 562350
rect 435774 562294 435842 562350
rect 435898 562294 435966 562350
rect 436022 562294 466314 562350
rect 466370 562294 466438 562350
rect 466494 562294 466562 562350
rect 466618 562294 466686 562350
rect 466742 562294 497034 562350
rect 497090 562294 497158 562350
rect 497214 562294 497282 562350
rect 497338 562294 497406 562350
rect 497462 562294 527754 562350
rect 527810 562294 527878 562350
rect 527934 562294 528002 562350
rect 528058 562294 528126 562350
rect 528182 562294 558474 562350
rect 558530 562294 558598 562350
rect 558654 562294 558722 562350
rect 558778 562294 558846 562350
rect 558902 562294 589194 562350
rect 589250 562294 589318 562350
rect 589374 562294 589442 562350
rect 589498 562294 589566 562350
rect 589622 562294 596496 562350
rect 596552 562294 596620 562350
rect 596676 562294 596744 562350
rect 596800 562294 596868 562350
rect 596924 562294 597980 562350
rect -1916 562226 597980 562294
rect -1916 562170 -860 562226
rect -804 562170 -736 562226
rect -680 562170 -612 562226
rect -556 562170 -488 562226
rect -432 562170 5514 562226
rect 5570 562170 5638 562226
rect 5694 562170 5762 562226
rect 5818 562170 5886 562226
rect 5942 562170 36234 562226
rect 36290 562170 36358 562226
rect 36414 562170 36482 562226
rect 36538 562170 36606 562226
rect 36662 562170 66954 562226
rect 67010 562170 67078 562226
rect 67134 562170 67202 562226
rect 67258 562170 67326 562226
rect 67382 562170 97674 562226
rect 97730 562170 97798 562226
rect 97854 562170 97922 562226
rect 97978 562170 98046 562226
rect 98102 562170 128394 562226
rect 128450 562170 128518 562226
rect 128574 562170 128642 562226
rect 128698 562170 128766 562226
rect 128822 562170 159114 562226
rect 159170 562170 159238 562226
rect 159294 562170 159362 562226
rect 159418 562170 159486 562226
rect 159542 562170 189834 562226
rect 189890 562170 189958 562226
rect 190014 562170 190082 562226
rect 190138 562170 190206 562226
rect 190262 562170 220554 562226
rect 220610 562170 220678 562226
rect 220734 562170 220802 562226
rect 220858 562170 220926 562226
rect 220982 562170 251274 562226
rect 251330 562170 251398 562226
rect 251454 562170 251522 562226
rect 251578 562170 251646 562226
rect 251702 562170 281994 562226
rect 282050 562170 282118 562226
rect 282174 562170 282242 562226
rect 282298 562170 282366 562226
rect 282422 562170 312714 562226
rect 312770 562170 312838 562226
rect 312894 562170 312962 562226
rect 313018 562170 313086 562226
rect 313142 562170 343434 562226
rect 343490 562170 343558 562226
rect 343614 562170 343682 562226
rect 343738 562170 343806 562226
rect 343862 562170 374154 562226
rect 374210 562170 374278 562226
rect 374334 562170 374402 562226
rect 374458 562170 374526 562226
rect 374582 562170 404874 562226
rect 404930 562170 404998 562226
rect 405054 562170 405122 562226
rect 405178 562170 405246 562226
rect 405302 562170 435594 562226
rect 435650 562170 435718 562226
rect 435774 562170 435842 562226
rect 435898 562170 435966 562226
rect 436022 562170 466314 562226
rect 466370 562170 466438 562226
rect 466494 562170 466562 562226
rect 466618 562170 466686 562226
rect 466742 562170 497034 562226
rect 497090 562170 497158 562226
rect 497214 562170 497282 562226
rect 497338 562170 497406 562226
rect 497462 562170 527754 562226
rect 527810 562170 527878 562226
rect 527934 562170 528002 562226
rect 528058 562170 528126 562226
rect 528182 562170 558474 562226
rect 558530 562170 558598 562226
rect 558654 562170 558722 562226
rect 558778 562170 558846 562226
rect 558902 562170 589194 562226
rect 589250 562170 589318 562226
rect 589374 562170 589442 562226
rect 589498 562170 589566 562226
rect 589622 562170 596496 562226
rect 596552 562170 596620 562226
rect 596676 562170 596744 562226
rect 596800 562170 596868 562226
rect 596924 562170 597980 562226
rect -1916 562102 597980 562170
rect -1916 562046 -860 562102
rect -804 562046 -736 562102
rect -680 562046 -612 562102
rect -556 562046 -488 562102
rect -432 562046 5514 562102
rect 5570 562046 5638 562102
rect 5694 562046 5762 562102
rect 5818 562046 5886 562102
rect 5942 562046 36234 562102
rect 36290 562046 36358 562102
rect 36414 562046 36482 562102
rect 36538 562046 36606 562102
rect 36662 562046 66954 562102
rect 67010 562046 67078 562102
rect 67134 562046 67202 562102
rect 67258 562046 67326 562102
rect 67382 562046 97674 562102
rect 97730 562046 97798 562102
rect 97854 562046 97922 562102
rect 97978 562046 98046 562102
rect 98102 562046 128394 562102
rect 128450 562046 128518 562102
rect 128574 562046 128642 562102
rect 128698 562046 128766 562102
rect 128822 562046 159114 562102
rect 159170 562046 159238 562102
rect 159294 562046 159362 562102
rect 159418 562046 159486 562102
rect 159542 562046 189834 562102
rect 189890 562046 189958 562102
rect 190014 562046 190082 562102
rect 190138 562046 190206 562102
rect 190262 562046 220554 562102
rect 220610 562046 220678 562102
rect 220734 562046 220802 562102
rect 220858 562046 220926 562102
rect 220982 562046 251274 562102
rect 251330 562046 251398 562102
rect 251454 562046 251522 562102
rect 251578 562046 251646 562102
rect 251702 562046 281994 562102
rect 282050 562046 282118 562102
rect 282174 562046 282242 562102
rect 282298 562046 282366 562102
rect 282422 562046 312714 562102
rect 312770 562046 312838 562102
rect 312894 562046 312962 562102
rect 313018 562046 313086 562102
rect 313142 562046 343434 562102
rect 343490 562046 343558 562102
rect 343614 562046 343682 562102
rect 343738 562046 343806 562102
rect 343862 562046 374154 562102
rect 374210 562046 374278 562102
rect 374334 562046 374402 562102
rect 374458 562046 374526 562102
rect 374582 562046 404874 562102
rect 404930 562046 404998 562102
rect 405054 562046 405122 562102
rect 405178 562046 405246 562102
rect 405302 562046 435594 562102
rect 435650 562046 435718 562102
rect 435774 562046 435842 562102
rect 435898 562046 435966 562102
rect 436022 562046 466314 562102
rect 466370 562046 466438 562102
rect 466494 562046 466562 562102
rect 466618 562046 466686 562102
rect 466742 562046 497034 562102
rect 497090 562046 497158 562102
rect 497214 562046 497282 562102
rect 497338 562046 497406 562102
rect 497462 562046 527754 562102
rect 527810 562046 527878 562102
rect 527934 562046 528002 562102
rect 528058 562046 528126 562102
rect 528182 562046 558474 562102
rect 558530 562046 558598 562102
rect 558654 562046 558722 562102
rect 558778 562046 558846 562102
rect 558902 562046 589194 562102
rect 589250 562046 589318 562102
rect 589374 562046 589442 562102
rect 589498 562046 589566 562102
rect 589622 562046 596496 562102
rect 596552 562046 596620 562102
rect 596676 562046 596744 562102
rect 596800 562046 596868 562102
rect 596924 562046 597980 562102
rect -1916 561978 597980 562046
rect -1916 561922 -860 561978
rect -804 561922 -736 561978
rect -680 561922 -612 561978
rect -556 561922 -488 561978
rect -432 561922 5514 561978
rect 5570 561922 5638 561978
rect 5694 561922 5762 561978
rect 5818 561922 5886 561978
rect 5942 561922 36234 561978
rect 36290 561922 36358 561978
rect 36414 561922 36482 561978
rect 36538 561922 36606 561978
rect 36662 561922 66954 561978
rect 67010 561922 67078 561978
rect 67134 561922 67202 561978
rect 67258 561922 67326 561978
rect 67382 561922 97674 561978
rect 97730 561922 97798 561978
rect 97854 561922 97922 561978
rect 97978 561922 98046 561978
rect 98102 561922 128394 561978
rect 128450 561922 128518 561978
rect 128574 561922 128642 561978
rect 128698 561922 128766 561978
rect 128822 561922 159114 561978
rect 159170 561922 159238 561978
rect 159294 561922 159362 561978
rect 159418 561922 159486 561978
rect 159542 561922 189834 561978
rect 189890 561922 189958 561978
rect 190014 561922 190082 561978
rect 190138 561922 190206 561978
rect 190262 561922 220554 561978
rect 220610 561922 220678 561978
rect 220734 561922 220802 561978
rect 220858 561922 220926 561978
rect 220982 561922 251274 561978
rect 251330 561922 251398 561978
rect 251454 561922 251522 561978
rect 251578 561922 251646 561978
rect 251702 561922 281994 561978
rect 282050 561922 282118 561978
rect 282174 561922 282242 561978
rect 282298 561922 282366 561978
rect 282422 561922 312714 561978
rect 312770 561922 312838 561978
rect 312894 561922 312962 561978
rect 313018 561922 313086 561978
rect 313142 561922 343434 561978
rect 343490 561922 343558 561978
rect 343614 561922 343682 561978
rect 343738 561922 343806 561978
rect 343862 561922 374154 561978
rect 374210 561922 374278 561978
rect 374334 561922 374402 561978
rect 374458 561922 374526 561978
rect 374582 561922 404874 561978
rect 404930 561922 404998 561978
rect 405054 561922 405122 561978
rect 405178 561922 405246 561978
rect 405302 561922 435594 561978
rect 435650 561922 435718 561978
rect 435774 561922 435842 561978
rect 435898 561922 435966 561978
rect 436022 561922 466314 561978
rect 466370 561922 466438 561978
rect 466494 561922 466562 561978
rect 466618 561922 466686 561978
rect 466742 561922 497034 561978
rect 497090 561922 497158 561978
rect 497214 561922 497282 561978
rect 497338 561922 497406 561978
rect 497462 561922 527754 561978
rect 527810 561922 527878 561978
rect 527934 561922 528002 561978
rect 528058 561922 528126 561978
rect 528182 561922 558474 561978
rect 558530 561922 558598 561978
rect 558654 561922 558722 561978
rect 558778 561922 558846 561978
rect 558902 561922 589194 561978
rect 589250 561922 589318 561978
rect 589374 561922 589442 561978
rect 589498 561922 589566 561978
rect 589622 561922 596496 561978
rect 596552 561922 596620 561978
rect 596676 561922 596744 561978
rect 596800 561922 596868 561978
rect 596924 561922 597980 561978
rect -1916 561826 597980 561922
rect -1916 550350 597980 550446
rect -1916 550294 -1820 550350
rect -1764 550294 -1696 550350
rect -1640 550294 -1572 550350
rect -1516 550294 -1448 550350
rect -1392 550294 9234 550350
rect 9290 550294 9358 550350
rect 9414 550294 9482 550350
rect 9538 550294 9606 550350
rect 9662 550294 39954 550350
rect 40010 550294 40078 550350
rect 40134 550294 40202 550350
rect 40258 550294 40326 550350
rect 40382 550294 70674 550350
rect 70730 550294 70798 550350
rect 70854 550294 70922 550350
rect 70978 550294 71046 550350
rect 71102 550294 101394 550350
rect 101450 550294 101518 550350
rect 101574 550294 101642 550350
rect 101698 550294 101766 550350
rect 101822 550294 132114 550350
rect 132170 550294 132238 550350
rect 132294 550294 132362 550350
rect 132418 550294 132486 550350
rect 132542 550294 162834 550350
rect 162890 550294 162958 550350
rect 163014 550294 163082 550350
rect 163138 550294 163206 550350
rect 163262 550294 193554 550350
rect 193610 550294 193678 550350
rect 193734 550294 193802 550350
rect 193858 550294 193926 550350
rect 193982 550294 224274 550350
rect 224330 550294 224398 550350
rect 224454 550294 224522 550350
rect 224578 550294 224646 550350
rect 224702 550294 254994 550350
rect 255050 550294 255118 550350
rect 255174 550294 255242 550350
rect 255298 550294 255366 550350
rect 255422 550294 285714 550350
rect 285770 550294 285838 550350
rect 285894 550294 285962 550350
rect 286018 550294 286086 550350
rect 286142 550294 316434 550350
rect 316490 550294 316558 550350
rect 316614 550294 316682 550350
rect 316738 550294 316806 550350
rect 316862 550294 347154 550350
rect 347210 550294 347278 550350
rect 347334 550294 347402 550350
rect 347458 550294 347526 550350
rect 347582 550294 377874 550350
rect 377930 550294 377998 550350
rect 378054 550294 378122 550350
rect 378178 550294 378246 550350
rect 378302 550294 408594 550350
rect 408650 550294 408718 550350
rect 408774 550294 408842 550350
rect 408898 550294 408966 550350
rect 409022 550294 439314 550350
rect 439370 550294 439438 550350
rect 439494 550294 439562 550350
rect 439618 550294 439686 550350
rect 439742 550294 470034 550350
rect 470090 550294 470158 550350
rect 470214 550294 470282 550350
rect 470338 550294 470406 550350
rect 470462 550294 500754 550350
rect 500810 550294 500878 550350
rect 500934 550294 501002 550350
rect 501058 550294 501126 550350
rect 501182 550294 531474 550350
rect 531530 550294 531598 550350
rect 531654 550294 531722 550350
rect 531778 550294 531846 550350
rect 531902 550294 562194 550350
rect 562250 550294 562318 550350
rect 562374 550294 562442 550350
rect 562498 550294 562566 550350
rect 562622 550294 592914 550350
rect 592970 550294 593038 550350
rect 593094 550294 593162 550350
rect 593218 550294 593286 550350
rect 593342 550294 597456 550350
rect 597512 550294 597580 550350
rect 597636 550294 597704 550350
rect 597760 550294 597828 550350
rect 597884 550294 597980 550350
rect -1916 550226 597980 550294
rect -1916 550170 -1820 550226
rect -1764 550170 -1696 550226
rect -1640 550170 -1572 550226
rect -1516 550170 -1448 550226
rect -1392 550170 9234 550226
rect 9290 550170 9358 550226
rect 9414 550170 9482 550226
rect 9538 550170 9606 550226
rect 9662 550170 39954 550226
rect 40010 550170 40078 550226
rect 40134 550170 40202 550226
rect 40258 550170 40326 550226
rect 40382 550170 70674 550226
rect 70730 550170 70798 550226
rect 70854 550170 70922 550226
rect 70978 550170 71046 550226
rect 71102 550170 101394 550226
rect 101450 550170 101518 550226
rect 101574 550170 101642 550226
rect 101698 550170 101766 550226
rect 101822 550170 132114 550226
rect 132170 550170 132238 550226
rect 132294 550170 132362 550226
rect 132418 550170 132486 550226
rect 132542 550170 162834 550226
rect 162890 550170 162958 550226
rect 163014 550170 163082 550226
rect 163138 550170 163206 550226
rect 163262 550170 193554 550226
rect 193610 550170 193678 550226
rect 193734 550170 193802 550226
rect 193858 550170 193926 550226
rect 193982 550170 224274 550226
rect 224330 550170 224398 550226
rect 224454 550170 224522 550226
rect 224578 550170 224646 550226
rect 224702 550170 254994 550226
rect 255050 550170 255118 550226
rect 255174 550170 255242 550226
rect 255298 550170 255366 550226
rect 255422 550170 285714 550226
rect 285770 550170 285838 550226
rect 285894 550170 285962 550226
rect 286018 550170 286086 550226
rect 286142 550170 316434 550226
rect 316490 550170 316558 550226
rect 316614 550170 316682 550226
rect 316738 550170 316806 550226
rect 316862 550170 347154 550226
rect 347210 550170 347278 550226
rect 347334 550170 347402 550226
rect 347458 550170 347526 550226
rect 347582 550170 377874 550226
rect 377930 550170 377998 550226
rect 378054 550170 378122 550226
rect 378178 550170 378246 550226
rect 378302 550170 408594 550226
rect 408650 550170 408718 550226
rect 408774 550170 408842 550226
rect 408898 550170 408966 550226
rect 409022 550170 439314 550226
rect 439370 550170 439438 550226
rect 439494 550170 439562 550226
rect 439618 550170 439686 550226
rect 439742 550170 470034 550226
rect 470090 550170 470158 550226
rect 470214 550170 470282 550226
rect 470338 550170 470406 550226
rect 470462 550170 500754 550226
rect 500810 550170 500878 550226
rect 500934 550170 501002 550226
rect 501058 550170 501126 550226
rect 501182 550170 531474 550226
rect 531530 550170 531598 550226
rect 531654 550170 531722 550226
rect 531778 550170 531846 550226
rect 531902 550170 562194 550226
rect 562250 550170 562318 550226
rect 562374 550170 562442 550226
rect 562498 550170 562566 550226
rect 562622 550170 592914 550226
rect 592970 550170 593038 550226
rect 593094 550170 593162 550226
rect 593218 550170 593286 550226
rect 593342 550170 597456 550226
rect 597512 550170 597580 550226
rect 597636 550170 597704 550226
rect 597760 550170 597828 550226
rect 597884 550170 597980 550226
rect -1916 550102 597980 550170
rect -1916 550046 -1820 550102
rect -1764 550046 -1696 550102
rect -1640 550046 -1572 550102
rect -1516 550046 -1448 550102
rect -1392 550046 9234 550102
rect 9290 550046 9358 550102
rect 9414 550046 9482 550102
rect 9538 550046 9606 550102
rect 9662 550046 39954 550102
rect 40010 550046 40078 550102
rect 40134 550046 40202 550102
rect 40258 550046 40326 550102
rect 40382 550046 70674 550102
rect 70730 550046 70798 550102
rect 70854 550046 70922 550102
rect 70978 550046 71046 550102
rect 71102 550046 101394 550102
rect 101450 550046 101518 550102
rect 101574 550046 101642 550102
rect 101698 550046 101766 550102
rect 101822 550046 132114 550102
rect 132170 550046 132238 550102
rect 132294 550046 132362 550102
rect 132418 550046 132486 550102
rect 132542 550046 162834 550102
rect 162890 550046 162958 550102
rect 163014 550046 163082 550102
rect 163138 550046 163206 550102
rect 163262 550046 193554 550102
rect 193610 550046 193678 550102
rect 193734 550046 193802 550102
rect 193858 550046 193926 550102
rect 193982 550046 224274 550102
rect 224330 550046 224398 550102
rect 224454 550046 224522 550102
rect 224578 550046 224646 550102
rect 224702 550046 254994 550102
rect 255050 550046 255118 550102
rect 255174 550046 255242 550102
rect 255298 550046 255366 550102
rect 255422 550046 285714 550102
rect 285770 550046 285838 550102
rect 285894 550046 285962 550102
rect 286018 550046 286086 550102
rect 286142 550046 316434 550102
rect 316490 550046 316558 550102
rect 316614 550046 316682 550102
rect 316738 550046 316806 550102
rect 316862 550046 347154 550102
rect 347210 550046 347278 550102
rect 347334 550046 347402 550102
rect 347458 550046 347526 550102
rect 347582 550046 377874 550102
rect 377930 550046 377998 550102
rect 378054 550046 378122 550102
rect 378178 550046 378246 550102
rect 378302 550046 408594 550102
rect 408650 550046 408718 550102
rect 408774 550046 408842 550102
rect 408898 550046 408966 550102
rect 409022 550046 439314 550102
rect 439370 550046 439438 550102
rect 439494 550046 439562 550102
rect 439618 550046 439686 550102
rect 439742 550046 470034 550102
rect 470090 550046 470158 550102
rect 470214 550046 470282 550102
rect 470338 550046 470406 550102
rect 470462 550046 500754 550102
rect 500810 550046 500878 550102
rect 500934 550046 501002 550102
rect 501058 550046 501126 550102
rect 501182 550046 531474 550102
rect 531530 550046 531598 550102
rect 531654 550046 531722 550102
rect 531778 550046 531846 550102
rect 531902 550046 562194 550102
rect 562250 550046 562318 550102
rect 562374 550046 562442 550102
rect 562498 550046 562566 550102
rect 562622 550046 592914 550102
rect 592970 550046 593038 550102
rect 593094 550046 593162 550102
rect 593218 550046 593286 550102
rect 593342 550046 597456 550102
rect 597512 550046 597580 550102
rect 597636 550046 597704 550102
rect 597760 550046 597828 550102
rect 597884 550046 597980 550102
rect -1916 549978 597980 550046
rect -1916 549922 -1820 549978
rect -1764 549922 -1696 549978
rect -1640 549922 -1572 549978
rect -1516 549922 -1448 549978
rect -1392 549922 9234 549978
rect 9290 549922 9358 549978
rect 9414 549922 9482 549978
rect 9538 549922 9606 549978
rect 9662 549922 39954 549978
rect 40010 549922 40078 549978
rect 40134 549922 40202 549978
rect 40258 549922 40326 549978
rect 40382 549922 70674 549978
rect 70730 549922 70798 549978
rect 70854 549922 70922 549978
rect 70978 549922 71046 549978
rect 71102 549922 101394 549978
rect 101450 549922 101518 549978
rect 101574 549922 101642 549978
rect 101698 549922 101766 549978
rect 101822 549922 132114 549978
rect 132170 549922 132238 549978
rect 132294 549922 132362 549978
rect 132418 549922 132486 549978
rect 132542 549922 162834 549978
rect 162890 549922 162958 549978
rect 163014 549922 163082 549978
rect 163138 549922 163206 549978
rect 163262 549922 193554 549978
rect 193610 549922 193678 549978
rect 193734 549922 193802 549978
rect 193858 549922 193926 549978
rect 193982 549922 224274 549978
rect 224330 549922 224398 549978
rect 224454 549922 224522 549978
rect 224578 549922 224646 549978
rect 224702 549922 254994 549978
rect 255050 549922 255118 549978
rect 255174 549922 255242 549978
rect 255298 549922 255366 549978
rect 255422 549922 285714 549978
rect 285770 549922 285838 549978
rect 285894 549922 285962 549978
rect 286018 549922 286086 549978
rect 286142 549922 316434 549978
rect 316490 549922 316558 549978
rect 316614 549922 316682 549978
rect 316738 549922 316806 549978
rect 316862 549922 347154 549978
rect 347210 549922 347278 549978
rect 347334 549922 347402 549978
rect 347458 549922 347526 549978
rect 347582 549922 377874 549978
rect 377930 549922 377998 549978
rect 378054 549922 378122 549978
rect 378178 549922 378246 549978
rect 378302 549922 408594 549978
rect 408650 549922 408718 549978
rect 408774 549922 408842 549978
rect 408898 549922 408966 549978
rect 409022 549922 439314 549978
rect 439370 549922 439438 549978
rect 439494 549922 439562 549978
rect 439618 549922 439686 549978
rect 439742 549922 470034 549978
rect 470090 549922 470158 549978
rect 470214 549922 470282 549978
rect 470338 549922 470406 549978
rect 470462 549922 500754 549978
rect 500810 549922 500878 549978
rect 500934 549922 501002 549978
rect 501058 549922 501126 549978
rect 501182 549922 531474 549978
rect 531530 549922 531598 549978
rect 531654 549922 531722 549978
rect 531778 549922 531846 549978
rect 531902 549922 562194 549978
rect 562250 549922 562318 549978
rect 562374 549922 562442 549978
rect 562498 549922 562566 549978
rect 562622 549922 592914 549978
rect 592970 549922 593038 549978
rect 593094 549922 593162 549978
rect 593218 549922 593286 549978
rect 593342 549922 597456 549978
rect 597512 549922 597580 549978
rect 597636 549922 597704 549978
rect 597760 549922 597828 549978
rect 597884 549922 597980 549978
rect -1916 549826 597980 549922
rect -1916 544350 597980 544446
rect -1916 544294 -860 544350
rect -804 544294 -736 544350
rect -680 544294 -612 544350
rect -556 544294 -488 544350
rect -432 544294 5514 544350
rect 5570 544294 5638 544350
rect 5694 544294 5762 544350
rect 5818 544294 5886 544350
rect 5942 544294 36234 544350
rect 36290 544294 36358 544350
rect 36414 544294 36482 544350
rect 36538 544294 36606 544350
rect 36662 544294 66954 544350
rect 67010 544294 67078 544350
rect 67134 544294 67202 544350
rect 67258 544294 67326 544350
rect 67382 544294 97674 544350
rect 97730 544294 97798 544350
rect 97854 544294 97922 544350
rect 97978 544294 98046 544350
rect 98102 544294 128394 544350
rect 128450 544294 128518 544350
rect 128574 544294 128642 544350
rect 128698 544294 128766 544350
rect 128822 544294 159114 544350
rect 159170 544294 159238 544350
rect 159294 544294 159362 544350
rect 159418 544294 159486 544350
rect 159542 544294 189834 544350
rect 189890 544294 189958 544350
rect 190014 544294 190082 544350
rect 190138 544294 190206 544350
rect 190262 544294 220554 544350
rect 220610 544294 220678 544350
rect 220734 544294 220802 544350
rect 220858 544294 220926 544350
rect 220982 544294 251274 544350
rect 251330 544294 251398 544350
rect 251454 544294 251522 544350
rect 251578 544294 251646 544350
rect 251702 544294 281994 544350
rect 282050 544294 282118 544350
rect 282174 544294 282242 544350
rect 282298 544294 282366 544350
rect 282422 544294 312714 544350
rect 312770 544294 312838 544350
rect 312894 544294 312962 544350
rect 313018 544294 313086 544350
rect 313142 544294 343434 544350
rect 343490 544294 343558 544350
rect 343614 544294 343682 544350
rect 343738 544294 343806 544350
rect 343862 544294 374154 544350
rect 374210 544294 374278 544350
rect 374334 544294 374402 544350
rect 374458 544294 374526 544350
rect 374582 544294 404874 544350
rect 404930 544294 404998 544350
rect 405054 544294 405122 544350
rect 405178 544294 405246 544350
rect 405302 544294 435594 544350
rect 435650 544294 435718 544350
rect 435774 544294 435842 544350
rect 435898 544294 435966 544350
rect 436022 544294 466314 544350
rect 466370 544294 466438 544350
rect 466494 544294 466562 544350
rect 466618 544294 466686 544350
rect 466742 544294 497034 544350
rect 497090 544294 497158 544350
rect 497214 544294 497282 544350
rect 497338 544294 497406 544350
rect 497462 544294 527754 544350
rect 527810 544294 527878 544350
rect 527934 544294 528002 544350
rect 528058 544294 528126 544350
rect 528182 544294 558474 544350
rect 558530 544294 558598 544350
rect 558654 544294 558722 544350
rect 558778 544294 558846 544350
rect 558902 544294 589194 544350
rect 589250 544294 589318 544350
rect 589374 544294 589442 544350
rect 589498 544294 589566 544350
rect 589622 544294 596496 544350
rect 596552 544294 596620 544350
rect 596676 544294 596744 544350
rect 596800 544294 596868 544350
rect 596924 544294 597980 544350
rect -1916 544226 597980 544294
rect -1916 544170 -860 544226
rect -804 544170 -736 544226
rect -680 544170 -612 544226
rect -556 544170 -488 544226
rect -432 544170 5514 544226
rect 5570 544170 5638 544226
rect 5694 544170 5762 544226
rect 5818 544170 5886 544226
rect 5942 544170 36234 544226
rect 36290 544170 36358 544226
rect 36414 544170 36482 544226
rect 36538 544170 36606 544226
rect 36662 544170 66954 544226
rect 67010 544170 67078 544226
rect 67134 544170 67202 544226
rect 67258 544170 67326 544226
rect 67382 544170 97674 544226
rect 97730 544170 97798 544226
rect 97854 544170 97922 544226
rect 97978 544170 98046 544226
rect 98102 544170 128394 544226
rect 128450 544170 128518 544226
rect 128574 544170 128642 544226
rect 128698 544170 128766 544226
rect 128822 544170 159114 544226
rect 159170 544170 159238 544226
rect 159294 544170 159362 544226
rect 159418 544170 159486 544226
rect 159542 544170 189834 544226
rect 189890 544170 189958 544226
rect 190014 544170 190082 544226
rect 190138 544170 190206 544226
rect 190262 544170 220554 544226
rect 220610 544170 220678 544226
rect 220734 544170 220802 544226
rect 220858 544170 220926 544226
rect 220982 544170 251274 544226
rect 251330 544170 251398 544226
rect 251454 544170 251522 544226
rect 251578 544170 251646 544226
rect 251702 544170 281994 544226
rect 282050 544170 282118 544226
rect 282174 544170 282242 544226
rect 282298 544170 282366 544226
rect 282422 544170 312714 544226
rect 312770 544170 312838 544226
rect 312894 544170 312962 544226
rect 313018 544170 313086 544226
rect 313142 544170 343434 544226
rect 343490 544170 343558 544226
rect 343614 544170 343682 544226
rect 343738 544170 343806 544226
rect 343862 544170 374154 544226
rect 374210 544170 374278 544226
rect 374334 544170 374402 544226
rect 374458 544170 374526 544226
rect 374582 544170 404874 544226
rect 404930 544170 404998 544226
rect 405054 544170 405122 544226
rect 405178 544170 405246 544226
rect 405302 544170 435594 544226
rect 435650 544170 435718 544226
rect 435774 544170 435842 544226
rect 435898 544170 435966 544226
rect 436022 544170 466314 544226
rect 466370 544170 466438 544226
rect 466494 544170 466562 544226
rect 466618 544170 466686 544226
rect 466742 544170 497034 544226
rect 497090 544170 497158 544226
rect 497214 544170 497282 544226
rect 497338 544170 497406 544226
rect 497462 544170 527754 544226
rect 527810 544170 527878 544226
rect 527934 544170 528002 544226
rect 528058 544170 528126 544226
rect 528182 544170 558474 544226
rect 558530 544170 558598 544226
rect 558654 544170 558722 544226
rect 558778 544170 558846 544226
rect 558902 544170 589194 544226
rect 589250 544170 589318 544226
rect 589374 544170 589442 544226
rect 589498 544170 589566 544226
rect 589622 544170 596496 544226
rect 596552 544170 596620 544226
rect 596676 544170 596744 544226
rect 596800 544170 596868 544226
rect 596924 544170 597980 544226
rect -1916 544102 597980 544170
rect -1916 544046 -860 544102
rect -804 544046 -736 544102
rect -680 544046 -612 544102
rect -556 544046 -488 544102
rect -432 544046 5514 544102
rect 5570 544046 5638 544102
rect 5694 544046 5762 544102
rect 5818 544046 5886 544102
rect 5942 544046 36234 544102
rect 36290 544046 36358 544102
rect 36414 544046 36482 544102
rect 36538 544046 36606 544102
rect 36662 544046 66954 544102
rect 67010 544046 67078 544102
rect 67134 544046 67202 544102
rect 67258 544046 67326 544102
rect 67382 544046 97674 544102
rect 97730 544046 97798 544102
rect 97854 544046 97922 544102
rect 97978 544046 98046 544102
rect 98102 544046 128394 544102
rect 128450 544046 128518 544102
rect 128574 544046 128642 544102
rect 128698 544046 128766 544102
rect 128822 544046 159114 544102
rect 159170 544046 159238 544102
rect 159294 544046 159362 544102
rect 159418 544046 159486 544102
rect 159542 544046 189834 544102
rect 189890 544046 189958 544102
rect 190014 544046 190082 544102
rect 190138 544046 190206 544102
rect 190262 544046 220554 544102
rect 220610 544046 220678 544102
rect 220734 544046 220802 544102
rect 220858 544046 220926 544102
rect 220982 544046 251274 544102
rect 251330 544046 251398 544102
rect 251454 544046 251522 544102
rect 251578 544046 251646 544102
rect 251702 544046 281994 544102
rect 282050 544046 282118 544102
rect 282174 544046 282242 544102
rect 282298 544046 282366 544102
rect 282422 544046 312714 544102
rect 312770 544046 312838 544102
rect 312894 544046 312962 544102
rect 313018 544046 313086 544102
rect 313142 544046 343434 544102
rect 343490 544046 343558 544102
rect 343614 544046 343682 544102
rect 343738 544046 343806 544102
rect 343862 544046 374154 544102
rect 374210 544046 374278 544102
rect 374334 544046 374402 544102
rect 374458 544046 374526 544102
rect 374582 544046 404874 544102
rect 404930 544046 404998 544102
rect 405054 544046 405122 544102
rect 405178 544046 405246 544102
rect 405302 544046 435594 544102
rect 435650 544046 435718 544102
rect 435774 544046 435842 544102
rect 435898 544046 435966 544102
rect 436022 544046 466314 544102
rect 466370 544046 466438 544102
rect 466494 544046 466562 544102
rect 466618 544046 466686 544102
rect 466742 544046 497034 544102
rect 497090 544046 497158 544102
rect 497214 544046 497282 544102
rect 497338 544046 497406 544102
rect 497462 544046 527754 544102
rect 527810 544046 527878 544102
rect 527934 544046 528002 544102
rect 528058 544046 528126 544102
rect 528182 544046 558474 544102
rect 558530 544046 558598 544102
rect 558654 544046 558722 544102
rect 558778 544046 558846 544102
rect 558902 544046 589194 544102
rect 589250 544046 589318 544102
rect 589374 544046 589442 544102
rect 589498 544046 589566 544102
rect 589622 544046 596496 544102
rect 596552 544046 596620 544102
rect 596676 544046 596744 544102
rect 596800 544046 596868 544102
rect 596924 544046 597980 544102
rect -1916 543978 597980 544046
rect -1916 543922 -860 543978
rect -804 543922 -736 543978
rect -680 543922 -612 543978
rect -556 543922 -488 543978
rect -432 543922 5514 543978
rect 5570 543922 5638 543978
rect 5694 543922 5762 543978
rect 5818 543922 5886 543978
rect 5942 543922 36234 543978
rect 36290 543922 36358 543978
rect 36414 543922 36482 543978
rect 36538 543922 36606 543978
rect 36662 543922 66954 543978
rect 67010 543922 67078 543978
rect 67134 543922 67202 543978
rect 67258 543922 67326 543978
rect 67382 543922 97674 543978
rect 97730 543922 97798 543978
rect 97854 543922 97922 543978
rect 97978 543922 98046 543978
rect 98102 543922 128394 543978
rect 128450 543922 128518 543978
rect 128574 543922 128642 543978
rect 128698 543922 128766 543978
rect 128822 543922 159114 543978
rect 159170 543922 159238 543978
rect 159294 543922 159362 543978
rect 159418 543922 159486 543978
rect 159542 543922 189834 543978
rect 189890 543922 189958 543978
rect 190014 543922 190082 543978
rect 190138 543922 190206 543978
rect 190262 543922 220554 543978
rect 220610 543922 220678 543978
rect 220734 543922 220802 543978
rect 220858 543922 220926 543978
rect 220982 543922 251274 543978
rect 251330 543922 251398 543978
rect 251454 543922 251522 543978
rect 251578 543922 251646 543978
rect 251702 543922 281994 543978
rect 282050 543922 282118 543978
rect 282174 543922 282242 543978
rect 282298 543922 282366 543978
rect 282422 543922 312714 543978
rect 312770 543922 312838 543978
rect 312894 543922 312962 543978
rect 313018 543922 313086 543978
rect 313142 543922 343434 543978
rect 343490 543922 343558 543978
rect 343614 543922 343682 543978
rect 343738 543922 343806 543978
rect 343862 543922 374154 543978
rect 374210 543922 374278 543978
rect 374334 543922 374402 543978
rect 374458 543922 374526 543978
rect 374582 543922 404874 543978
rect 404930 543922 404998 543978
rect 405054 543922 405122 543978
rect 405178 543922 405246 543978
rect 405302 543922 435594 543978
rect 435650 543922 435718 543978
rect 435774 543922 435842 543978
rect 435898 543922 435966 543978
rect 436022 543922 466314 543978
rect 466370 543922 466438 543978
rect 466494 543922 466562 543978
rect 466618 543922 466686 543978
rect 466742 543922 497034 543978
rect 497090 543922 497158 543978
rect 497214 543922 497282 543978
rect 497338 543922 497406 543978
rect 497462 543922 527754 543978
rect 527810 543922 527878 543978
rect 527934 543922 528002 543978
rect 528058 543922 528126 543978
rect 528182 543922 558474 543978
rect 558530 543922 558598 543978
rect 558654 543922 558722 543978
rect 558778 543922 558846 543978
rect 558902 543922 589194 543978
rect 589250 543922 589318 543978
rect 589374 543922 589442 543978
rect 589498 543922 589566 543978
rect 589622 543922 596496 543978
rect 596552 543922 596620 543978
rect 596676 543922 596744 543978
rect 596800 543922 596868 543978
rect 596924 543922 597980 543978
rect -1916 543826 597980 543922
rect -1916 532350 597980 532446
rect -1916 532294 -1820 532350
rect -1764 532294 -1696 532350
rect -1640 532294 -1572 532350
rect -1516 532294 -1448 532350
rect -1392 532294 9234 532350
rect 9290 532294 9358 532350
rect 9414 532294 9482 532350
rect 9538 532294 9606 532350
rect 9662 532294 39954 532350
rect 40010 532294 40078 532350
rect 40134 532294 40202 532350
rect 40258 532294 40326 532350
rect 40382 532294 70674 532350
rect 70730 532294 70798 532350
rect 70854 532294 70922 532350
rect 70978 532294 71046 532350
rect 71102 532294 101394 532350
rect 101450 532294 101518 532350
rect 101574 532294 101642 532350
rect 101698 532294 101766 532350
rect 101822 532294 132114 532350
rect 132170 532294 132238 532350
rect 132294 532294 132362 532350
rect 132418 532294 132486 532350
rect 132542 532294 162834 532350
rect 162890 532294 162958 532350
rect 163014 532294 163082 532350
rect 163138 532294 163206 532350
rect 163262 532294 193554 532350
rect 193610 532294 193678 532350
rect 193734 532294 193802 532350
rect 193858 532294 193926 532350
rect 193982 532294 224274 532350
rect 224330 532294 224398 532350
rect 224454 532294 224522 532350
rect 224578 532294 224646 532350
rect 224702 532294 254994 532350
rect 255050 532294 255118 532350
rect 255174 532294 255242 532350
rect 255298 532294 255366 532350
rect 255422 532294 285714 532350
rect 285770 532294 285838 532350
rect 285894 532294 285962 532350
rect 286018 532294 286086 532350
rect 286142 532294 316434 532350
rect 316490 532294 316558 532350
rect 316614 532294 316682 532350
rect 316738 532294 316806 532350
rect 316862 532294 347154 532350
rect 347210 532294 347278 532350
rect 347334 532294 347402 532350
rect 347458 532294 347526 532350
rect 347582 532294 377874 532350
rect 377930 532294 377998 532350
rect 378054 532294 378122 532350
rect 378178 532294 378246 532350
rect 378302 532294 408594 532350
rect 408650 532294 408718 532350
rect 408774 532294 408842 532350
rect 408898 532294 408966 532350
rect 409022 532294 439314 532350
rect 439370 532294 439438 532350
rect 439494 532294 439562 532350
rect 439618 532294 439686 532350
rect 439742 532294 470034 532350
rect 470090 532294 470158 532350
rect 470214 532294 470282 532350
rect 470338 532294 470406 532350
rect 470462 532294 500754 532350
rect 500810 532294 500878 532350
rect 500934 532294 501002 532350
rect 501058 532294 501126 532350
rect 501182 532294 531474 532350
rect 531530 532294 531598 532350
rect 531654 532294 531722 532350
rect 531778 532294 531846 532350
rect 531902 532294 562194 532350
rect 562250 532294 562318 532350
rect 562374 532294 562442 532350
rect 562498 532294 562566 532350
rect 562622 532294 592914 532350
rect 592970 532294 593038 532350
rect 593094 532294 593162 532350
rect 593218 532294 593286 532350
rect 593342 532294 597456 532350
rect 597512 532294 597580 532350
rect 597636 532294 597704 532350
rect 597760 532294 597828 532350
rect 597884 532294 597980 532350
rect -1916 532226 597980 532294
rect -1916 532170 -1820 532226
rect -1764 532170 -1696 532226
rect -1640 532170 -1572 532226
rect -1516 532170 -1448 532226
rect -1392 532170 9234 532226
rect 9290 532170 9358 532226
rect 9414 532170 9482 532226
rect 9538 532170 9606 532226
rect 9662 532170 39954 532226
rect 40010 532170 40078 532226
rect 40134 532170 40202 532226
rect 40258 532170 40326 532226
rect 40382 532170 70674 532226
rect 70730 532170 70798 532226
rect 70854 532170 70922 532226
rect 70978 532170 71046 532226
rect 71102 532170 101394 532226
rect 101450 532170 101518 532226
rect 101574 532170 101642 532226
rect 101698 532170 101766 532226
rect 101822 532170 132114 532226
rect 132170 532170 132238 532226
rect 132294 532170 132362 532226
rect 132418 532170 132486 532226
rect 132542 532170 162834 532226
rect 162890 532170 162958 532226
rect 163014 532170 163082 532226
rect 163138 532170 163206 532226
rect 163262 532170 193554 532226
rect 193610 532170 193678 532226
rect 193734 532170 193802 532226
rect 193858 532170 193926 532226
rect 193982 532170 224274 532226
rect 224330 532170 224398 532226
rect 224454 532170 224522 532226
rect 224578 532170 224646 532226
rect 224702 532170 254994 532226
rect 255050 532170 255118 532226
rect 255174 532170 255242 532226
rect 255298 532170 255366 532226
rect 255422 532170 285714 532226
rect 285770 532170 285838 532226
rect 285894 532170 285962 532226
rect 286018 532170 286086 532226
rect 286142 532170 316434 532226
rect 316490 532170 316558 532226
rect 316614 532170 316682 532226
rect 316738 532170 316806 532226
rect 316862 532170 347154 532226
rect 347210 532170 347278 532226
rect 347334 532170 347402 532226
rect 347458 532170 347526 532226
rect 347582 532170 377874 532226
rect 377930 532170 377998 532226
rect 378054 532170 378122 532226
rect 378178 532170 378246 532226
rect 378302 532170 408594 532226
rect 408650 532170 408718 532226
rect 408774 532170 408842 532226
rect 408898 532170 408966 532226
rect 409022 532170 439314 532226
rect 439370 532170 439438 532226
rect 439494 532170 439562 532226
rect 439618 532170 439686 532226
rect 439742 532170 470034 532226
rect 470090 532170 470158 532226
rect 470214 532170 470282 532226
rect 470338 532170 470406 532226
rect 470462 532170 500754 532226
rect 500810 532170 500878 532226
rect 500934 532170 501002 532226
rect 501058 532170 501126 532226
rect 501182 532170 531474 532226
rect 531530 532170 531598 532226
rect 531654 532170 531722 532226
rect 531778 532170 531846 532226
rect 531902 532170 562194 532226
rect 562250 532170 562318 532226
rect 562374 532170 562442 532226
rect 562498 532170 562566 532226
rect 562622 532170 592914 532226
rect 592970 532170 593038 532226
rect 593094 532170 593162 532226
rect 593218 532170 593286 532226
rect 593342 532170 597456 532226
rect 597512 532170 597580 532226
rect 597636 532170 597704 532226
rect 597760 532170 597828 532226
rect 597884 532170 597980 532226
rect -1916 532102 597980 532170
rect -1916 532046 -1820 532102
rect -1764 532046 -1696 532102
rect -1640 532046 -1572 532102
rect -1516 532046 -1448 532102
rect -1392 532046 9234 532102
rect 9290 532046 9358 532102
rect 9414 532046 9482 532102
rect 9538 532046 9606 532102
rect 9662 532046 39954 532102
rect 40010 532046 40078 532102
rect 40134 532046 40202 532102
rect 40258 532046 40326 532102
rect 40382 532046 70674 532102
rect 70730 532046 70798 532102
rect 70854 532046 70922 532102
rect 70978 532046 71046 532102
rect 71102 532046 101394 532102
rect 101450 532046 101518 532102
rect 101574 532046 101642 532102
rect 101698 532046 101766 532102
rect 101822 532046 132114 532102
rect 132170 532046 132238 532102
rect 132294 532046 132362 532102
rect 132418 532046 132486 532102
rect 132542 532046 162834 532102
rect 162890 532046 162958 532102
rect 163014 532046 163082 532102
rect 163138 532046 163206 532102
rect 163262 532046 193554 532102
rect 193610 532046 193678 532102
rect 193734 532046 193802 532102
rect 193858 532046 193926 532102
rect 193982 532046 224274 532102
rect 224330 532046 224398 532102
rect 224454 532046 224522 532102
rect 224578 532046 224646 532102
rect 224702 532046 254994 532102
rect 255050 532046 255118 532102
rect 255174 532046 255242 532102
rect 255298 532046 255366 532102
rect 255422 532046 285714 532102
rect 285770 532046 285838 532102
rect 285894 532046 285962 532102
rect 286018 532046 286086 532102
rect 286142 532046 316434 532102
rect 316490 532046 316558 532102
rect 316614 532046 316682 532102
rect 316738 532046 316806 532102
rect 316862 532046 347154 532102
rect 347210 532046 347278 532102
rect 347334 532046 347402 532102
rect 347458 532046 347526 532102
rect 347582 532046 377874 532102
rect 377930 532046 377998 532102
rect 378054 532046 378122 532102
rect 378178 532046 378246 532102
rect 378302 532046 408594 532102
rect 408650 532046 408718 532102
rect 408774 532046 408842 532102
rect 408898 532046 408966 532102
rect 409022 532046 439314 532102
rect 439370 532046 439438 532102
rect 439494 532046 439562 532102
rect 439618 532046 439686 532102
rect 439742 532046 470034 532102
rect 470090 532046 470158 532102
rect 470214 532046 470282 532102
rect 470338 532046 470406 532102
rect 470462 532046 500754 532102
rect 500810 532046 500878 532102
rect 500934 532046 501002 532102
rect 501058 532046 501126 532102
rect 501182 532046 531474 532102
rect 531530 532046 531598 532102
rect 531654 532046 531722 532102
rect 531778 532046 531846 532102
rect 531902 532046 562194 532102
rect 562250 532046 562318 532102
rect 562374 532046 562442 532102
rect 562498 532046 562566 532102
rect 562622 532046 592914 532102
rect 592970 532046 593038 532102
rect 593094 532046 593162 532102
rect 593218 532046 593286 532102
rect 593342 532046 597456 532102
rect 597512 532046 597580 532102
rect 597636 532046 597704 532102
rect 597760 532046 597828 532102
rect 597884 532046 597980 532102
rect -1916 531978 597980 532046
rect -1916 531922 -1820 531978
rect -1764 531922 -1696 531978
rect -1640 531922 -1572 531978
rect -1516 531922 -1448 531978
rect -1392 531922 9234 531978
rect 9290 531922 9358 531978
rect 9414 531922 9482 531978
rect 9538 531922 9606 531978
rect 9662 531922 39954 531978
rect 40010 531922 40078 531978
rect 40134 531922 40202 531978
rect 40258 531922 40326 531978
rect 40382 531922 70674 531978
rect 70730 531922 70798 531978
rect 70854 531922 70922 531978
rect 70978 531922 71046 531978
rect 71102 531922 101394 531978
rect 101450 531922 101518 531978
rect 101574 531922 101642 531978
rect 101698 531922 101766 531978
rect 101822 531922 132114 531978
rect 132170 531922 132238 531978
rect 132294 531922 132362 531978
rect 132418 531922 132486 531978
rect 132542 531922 162834 531978
rect 162890 531922 162958 531978
rect 163014 531922 163082 531978
rect 163138 531922 163206 531978
rect 163262 531922 193554 531978
rect 193610 531922 193678 531978
rect 193734 531922 193802 531978
rect 193858 531922 193926 531978
rect 193982 531922 224274 531978
rect 224330 531922 224398 531978
rect 224454 531922 224522 531978
rect 224578 531922 224646 531978
rect 224702 531922 254994 531978
rect 255050 531922 255118 531978
rect 255174 531922 255242 531978
rect 255298 531922 255366 531978
rect 255422 531922 285714 531978
rect 285770 531922 285838 531978
rect 285894 531922 285962 531978
rect 286018 531922 286086 531978
rect 286142 531922 316434 531978
rect 316490 531922 316558 531978
rect 316614 531922 316682 531978
rect 316738 531922 316806 531978
rect 316862 531922 347154 531978
rect 347210 531922 347278 531978
rect 347334 531922 347402 531978
rect 347458 531922 347526 531978
rect 347582 531922 377874 531978
rect 377930 531922 377998 531978
rect 378054 531922 378122 531978
rect 378178 531922 378246 531978
rect 378302 531922 408594 531978
rect 408650 531922 408718 531978
rect 408774 531922 408842 531978
rect 408898 531922 408966 531978
rect 409022 531922 439314 531978
rect 439370 531922 439438 531978
rect 439494 531922 439562 531978
rect 439618 531922 439686 531978
rect 439742 531922 470034 531978
rect 470090 531922 470158 531978
rect 470214 531922 470282 531978
rect 470338 531922 470406 531978
rect 470462 531922 500754 531978
rect 500810 531922 500878 531978
rect 500934 531922 501002 531978
rect 501058 531922 501126 531978
rect 501182 531922 531474 531978
rect 531530 531922 531598 531978
rect 531654 531922 531722 531978
rect 531778 531922 531846 531978
rect 531902 531922 562194 531978
rect 562250 531922 562318 531978
rect 562374 531922 562442 531978
rect 562498 531922 562566 531978
rect 562622 531922 592914 531978
rect 592970 531922 593038 531978
rect 593094 531922 593162 531978
rect 593218 531922 593286 531978
rect 593342 531922 597456 531978
rect 597512 531922 597580 531978
rect 597636 531922 597704 531978
rect 597760 531922 597828 531978
rect 597884 531922 597980 531978
rect -1916 531826 597980 531922
rect -1916 526350 597980 526446
rect -1916 526294 -860 526350
rect -804 526294 -736 526350
rect -680 526294 -612 526350
rect -556 526294 -488 526350
rect -432 526294 5514 526350
rect 5570 526294 5638 526350
rect 5694 526294 5762 526350
rect 5818 526294 5886 526350
rect 5942 526294 36234 526350
rect 36290 526294 36358 526350
rect 36414 526294 36482 526350
rect 36538 526294 36606 526350
rect 36662 526294 66954 526350
rect 67010 526294 67078 526350
rect 67134 526294 67202 526350
rect 67258 526294 67326 526350
rect 67382 526294 97674 526350
rect 97730 526294 97798 526350
rect 97854 526294 97922 526350
rect 97978 526294 98046 526350
rect 98102 526294 128394 526350
rect 128450 526294 128518 526350
rect 128574 526294 128642 526350
rect 128698 526294 128766 526350
rect 128822 526294 159114 526350
rect 159170 526294 159238 526350
rect 159294 526294 159362 526350
rect 159418 526294 159486 526350
rect 159542 526294 189834 526350
rect 189890 526294 189958 526350
rect 190014 526294 190082 526350
rect 190138 526294 190206 526350
rect 190262 526294 220554 526350
rect 220610 526294 220678 526350
rect 220734 526294 220802 526350
rect 220858 526294 220926 526350
rect 220982 526294 251274 526350
rect 251330 526294 251398 526350
rect 251454 526294 251522 526350
rect 251578 526294 251646 526350
rect 251702 526294 281994 526350
rect 282050 526294 282118 526350
rect 282174 526294 282242 526350
rect 282298 526294 282366 526350
rect 282422 526294 312714 526350
rect 312770 526294 312838 526350
rect 312894 526294 312962 526350
rect 313018 526294 313086 526350
rect 313142 526294 343434 526350
rect 343490 526294 343558 526350
rect 343614 526294 343682 526350
rect 343738 526294 343806 526350
rect 343862 526294 374154 526350
rect 374210 526294 374278 526350
rect 374334 526294 374402 526350
rect 374458 526294 374526 526350
rect 374582 526294 404874 526350
rect 404930 526294 404998 526350
rect 405054 526294 405122 526350
rect 405178 526294 405246 526350
rect 405302 526294 435594 526350
rect 435650 526294 435718 526350
rect 435774 526294 435842 526350
rect 435898 526294 435966 526350
rect 436022 526294 466314 526350
rect 466370 526294 466438 526350
rect 466494 526294 466562 526350
rect 466618 526294 466686 526350
rect 466742 526294 497034 526350
rect 497090 526294 497158 526350
rect 497214 526294 497282 526350
rect 497338 526294 497406 526350
rect 497462 526294 527754 526350
rect 527810 526294 527878 526350
rect 527934 526294 528002 526350
rect 528058 526294 528126 526350
rect 528182 526294 558474 526350
rect 558530 526294 558598 526350
rect 558654 526294 558722 526350
rect 558778 526294 558846 526350
rect 558902 526294 589194 526350
rect 589250 526294 589318 526350
rect 589374 526294 589442 526350
rect 589498 526294 589566 526350
rect 589622 526294 596496 526350
rect 596552 526294 596620 526350
rect 596676 526294 596744 526350
rect 596800 526294 596868 526350
rect 596924 526294 597980 526350
rect -1916 526226 597980 526294
rect -1916 526170 -860 526226
rect -804 526170 -736 526226
rect -680 526170 -612 526226
rect -556 526170 -488 526226
rect -432 526170 5514 526226
rect 5570 526170 5638 526226
rect 5694 526170 5762 526226
rect 5818 526170 5886 526226
rect 5942 526170 36234 526226
rect 36290 526170 36358 526226
rect 36414 526170 36482 526226
rect 36538 526170 36606 526226
rect 36662 526170 66954 526226
rect 67010 526170 67078 526226
rect 67134 526170 67202 526226
rect 67258 526170 67326 526226
rect 67382 526170 97674 526226
rect 97730 526170 97798 526226
rect 97854 526170 97922 526226
rect 97978 526170 98046 526226
rect 98102 526170 128394 526226
rect 128450 526170 128518 526226
rect 128574 526170 128642 526226
rect 128698 526170 128766 526226
rect 128822 526170 159114 526226
rect 159170 526170 159238 526226
rect 159294 526170 159362 526226
rect 159418 526170 159486 526226
rect 159542 526170 189834 526226
rect 189890 526170 189958 526226
rect 190014 526170 190082 526226
rect 190138 526170 190206 526226
rect 190262 526170 220554 526226
rect 220610 526170 220678 526226
rect 220734 526170 220802 526226
rect 220858 526170 220926 526226
rect 220982 526170 251274 526226
rect 251330 526170 251398 526226
rect 251454 526170 251522 526226
rect 251578 526170 251646 526226
rect 251702 526170 281994 526226
rect 282050 526170 282118 526226
rect 282174 526170 282242 526226
rect 282298 526170 282366 526226
rect 282422 526170 312714 526226
rect 312770 526170 312838 526226
rect 312894 526170 312962 526226
rect 313018 526170 313086 526226
rect 313142 526170 343434 526226
rect 343490 526170 343558 526226
rect 343614 526170 343682 526226
rect 343738 526170 343806 526226
rect 343862 526170 374154 526226
rect 374210 526170 374278 526226
rect 374334 526170 374402 526226
rect 374458 526170 374526 526226
rect 374582 526170 404874 526226
rect 404930 526170 404998 526226
rect 405054 526170 405122 526226
rect 405178 526170 405246 526226
rect 405302 526170 435594 526226
rect 435650 526170 435718 526226
rect 435774 526170 435842 526226
rect 435898 526170 435966 526226
rect 436022 526170 466314 526226
rect 466370 526170 466438 526226
rect 466494 526170 466562 526226
rect 466618 526170 466686 526226
rect 466742 526170 497034 526226
rect 497090 526170 497158 526226
rect 497214 526170 497282 526226
rect 497338 526170 497406 526226
rect 497462 526170 527754 526226
rect 527810 526170 527878 526226
rect 527934 526170 528002 526226
rect 528058 526170 528126 526226
rect 528182 526170 558474 526226
rect 558530 526170 558598 526226
rect 558654 526170 558722 526226
rect 558778 526170 558846 526226
rect 558902 526170 589194 526226
rect 589250 526170 589318 526226
rect 589374 526170 589442 526226
rect 589498 526170 589566 526226
rect 589622 526170 596496 526226
rect 596552 526170 596620 526226
rect 596676 526170 596744 526226
rect 596800 526170 596868 526226
rect 596924 526170 597980 526226
rect -1916 526102 597980 526170
rect -1916 526046 -860 526102
rect -804 526046 -736 526102
rect -680 526046 -612 526102
rect -556 526046 -488 526102
rect -432 526046 5514 526102
rect 5570 526046 5638 526102
rect 5694 526046 5762 526102
rect 5818 526046 5886 526102
rect 5942 526046 36234 526102
rect 36290 526046 36358 526102
rect 36414 526046 36482 526102
rect 36538 526046 36606 526102
rect 36662 526046 66954 526102
rect 67010 526046 67078 526102
rect 67134 526046 67202 526102
rect 67258 526046 67326 526102
rect 67382 526046 97674 526102
rect 97730 526046 97798 526102
rect 97854 526046 97922 526102
rect 97978 526046 98046 526102
rect 98102 526046 128394 526102
rect 128450 526046 128518 526102
rect 128574 526046 128642 526102
rect 128698 526046 128766 526102
rect 128822 526046 159114 526102
rect 159170 526046 159238 526102
rect 159294 526046 159362 526102
rect 159418 526046 159486 526102
rect 159542 526046 189834 526102
rect 189890 526046 189958 526102
rect 190014 526046 190082 526102
rect 190138 526046 190206 526102
rect 190262 526046 220554 526102
rect 220610 526046 220678 526102
rect 220734 526046 220802 526102
rect 220858 526046 220926 526102
rect 220982 526046 251274 526102
rect 251330 526046 251398 526102
rect 251454 526046 251522 526102
rect 251578 526046 251646 526102
rect 251702 526046 281994 526102
rect 282050 526046 282118 526102
rect 282174 526046 282242 526102
rect 282298 526046 282366 526102
rect 282422 526046 312714 526102
rect 312770 526046 312838 526102
rect 312894 526046 312962 526102
rect 313018 526046 313086 526102
rect 313142 526046 343434 526102
rect 343490 526046 343558 526102
rect 343614 526046 343682 526102
rect 343738 526046 343806 526102
rect 343862 526046 374154 526102
rect 374210 526046 374278 526102
rect 374334 526046 374402 526102
rect 374458 526046 374526 526102
rect 374582 526046 404874 526102
rect 404930 526046 404998 526102
rect 405054 526046 405122 526102
rect 405178 526046 405246 526102
rect 405302 526046 435594 526102
rect 435650 526046 435718 526102
rect 435774 526046 435842 526102
rect 435898 526046 435966 526102
rect 436022 526046 466314 526102
rect 466370 526046 466438 526102
rect 466494 526046 466562 526102
rect 466618 526046 466686 526102
rect 466742 526046 497034 526102
rect 497090 526046 497158 526102
rect 497214 526046 497282 526102
rect 497338 526046 497406 526102
rect 497462 526046 527754 526102
rect 527810 526046 527878 526102
rect 527934 526046 528002 526102
rect 528058 526046 528126 526102
rect 528182 526046 558474 526102
rect 558530 526046 558598 526102
rect 558654 526046 558722 526102
rect 558778 526046 558846 526102
rect 558902 526046 589194 526102
rect 589250 526046 589318 526102
rect 589374 526046 589442 526102
rect 589498 526046 589566 526102
rect 589622 526046 596496 526102
rect 596552 526046 596620 526102
rect 596676 526046 596744 526102
rect 596800 526046 596868 526102
rect 596924 526046 597980 526102
rect -1916 525978 597980 526046
rect -1916 525922 -860 525978
rect -804 525922 -736 525978
rect -680 525922 -612 525978
rect -556 525922 -488 525978
rect -432 525922 5514 525978
rect 5570 525922 5638 525978
rect 5694 525922 5762 525978
rect 5818 525922 5886 525978
rect 5942 525922 36234 525978
rect 36290 525922 36358 525978
rect 36414 525922 36482 525978
rect 36538 525922 36606 525978
rect 36662 525922 66954 525978
rect 67010 525922 67078 525978
rect 67134 525922 67202 525978
rect 67258 525922 67326 525978
rect 67382 525922 97674 525978
rect 97730 525922 97798 525978
rect 97854 525922 97922 525978
rect 97978 525922 98046 525978
rect 98102 525922 128394 525978
rect 128450 525922 128518 525978
rect 128574 525922 128642 525978
rect 128698 525922 128766 525978
rect 128822 525922 159114 525978
rect 159170 525922 159238 525978
rect 159294 525922 159362 525978
rect 159418 525922 159486 525978
rect 159542 525922 189834 525978
rect 189890 525922 189958 525978
rect 190014 525922 190082 525978
rect 190138 525922 190206 525978
rect 190262 525922 220554 525978
rect 220610 525922 220678 525978
rect 220734 525922 220802 525978
rect 220858 525922 220926 525978
rect 220982 525922 251274 525978
rect 251330 525922 251398 525978
rect 251454 525922 251522 525978
rect 251578 525922 251646 525978
rect 251702 525922 281994 525978
rect 282050 525922 282118 525978
rect 282174 525922 282242 525978
rect 282298 525922 282366 525978
rect 282422 525922 312714 525978
rect 312770 525922 312838 525978
rect 312894 525922 312962 525978
rect 313018 525922 313086 525978
rect 313142 525922 343434 525978
rect 343490 525922 343558 525978
rect 343614 525922 343682 525978
rect 343738 525922 343806 525978
rect 343862 525922 374154 525978
rect 374210 525922 374278 525978
rect 374334 525922 374402 525978
rect 374458 525922 374526 525978
rect 374582 525922 404874 525978
rect 404930 525922 404998 525978
rect 405054 525922 405122 525978
rect 405178 525922 405246 525978
rect 405302 525922 435594 525978
rect 435650 525922 435718 525978
rect 435774 525922 435842 525978
rect 435898 525922 435966 525978
rect 436022 525922 466314 525978
rect 466370 525922 466438 525978
rect 466494 525922 466562 525978
rect 466618 525922 466686 525978
rect 466742 525922 497034 525978
rect 497090 525922 497158 525978
rect 497214 525922 497282 525978
rect 497338 525922 497406 525978
rect 497462 525922 527754 525978
rect 527810 525922 527878 525978
rect 527934 525922 528002 525978
rect 528058 525922 528126 525978
rect 528182 525922 558474 525978
rect 558530 525922 558598 525978
rect 558654 525922 558722 525978
rect 558778 525922 558846 525978
rect 558902 525922 589194 525978
rect 589250 525922 589318 525978
rect 589374 525922 589442 525978
rect 589498 525922 589566 525978
rect 589622 525922 596496 525978
rect 596552 525922 596620 525978
rect 596676 525922 596744 525978
rect 596800 525922 596868 525978
rect 596924 525922 597980 525978
rect -1916 525826 597980 525922
rect -1916 514350 597980 514446
rect -1916 514294 -1820 514350
rect -1764 514294 -1696 514350
rect -1640 514294 -1572 514350
rect -1516 514294 -1448 514350
rect -1392 514294 9234 514350
rect 9290 514294 9358 514350
rect 9414 514294 9482 514350
rect 9538 514294 9606 514350
rect 9662 514294 39954 514350
rect 40010 514294 40078 514350
rect 40134 514294 40202 514350
rect 40258 514294 40326 514350
rect 40382 514294 70674 514350
rect 70730 514294 70798 514350
rect 70854 514294 70922 514350
rect 70978 514294 71046 514350
rect 71102 514294 101394 514350
rect 101450 514294 101518 514350
rect 101574 514294 101642 514350
rect 101698 514294 101766 514350
rect 101822 514294 132114 514350
rect 132170 514294 132238 514350
rect 132294 514294 132362 514350
rect 132418 514294 132486 514350
rect 132542 514294 162834 514350
rect 162890 514294 162958 514350
rect 163014 514294 163082 514350
rect 163138 514294 163206 514350
rect 163262 514294 193554 514350
rect 193610 514294 193678 514350
rect 193734 514294 193802 514350
rect 193858 514294 193926 514350
rect 193982 514294 224274 514350
rect 224330 514294 224398 514350
rect 224454 514294 224522 514350
rect 224578 514294 224646 514350
rect 224702 514294 254994 514350
rect 255050 514294 255118 514350
rect 255174 514294 255242 514350
rect 255298 514294 255366 514350
rect 255422 514294 285714 514350
rect 285770 514294 285838 514350
rect 285894 514294 285962 514350
rect 286018 514294 286086 514350
rect 286142 514294 316434 514350
rect 316490 514294 316558 514350
rect 316614 514294 316682 514350
rect 316738 514294 316806 514350
rect 316862 514294 347154 514350
rect 347210 514294 347278 514350
rect 347334 514294 347402 514350
rect 347458 514294 347526 514350
rect 347582 514294 377874 514350
rect 377930 514294 377998 514350
rect 378054 514294 378122 514350
rect 378178 514294 378246 514350
rect 378302 514294 408594 514350
rect 408650 514294 408718 514350
rect 408774 514294 408842 514350
rect 408898 514294 408966 514350
rect 409022 514294 439314 514350
rect 439370 514294 439438 514350
rect 439494 514294 439562 514350
rect 439618 514294 439686 514350
rect 439742 514294 470034 514350
rect 470090 514294 470158 514350
rect 470214 514294 470282 514350
rect 470338 514294 470406 514350
rect 470462 514294 500754 514350
rect 500810 514294 500878 514350
rect 500934 514294 501002 514350
rect 501058 514294 501126 514350
rect 501182 514294 531474 514350
rect 531530 514294 531598 514350
rect 531654 514294 531722 514350
rect 531778 514294 531846 514350
rect 531902 514294 562194 514350
rect 562250 514294 562318 514350
rect 562374 514294 562442 514350
rect 562498 514294 562566 514350
rect 562622 514294 592914 514350
rect 592970 514294 593038 514350
rect 593094 514294 593162 514350
rect 593218 514294 593286 514350
rect 593342 514294 597456 514350
rect 597512 514294 597580 514350
rect 597636 514294 597704 514350
rect 597760 514294 597828 514350
rect 597884 514294 597980 514350
rect -1916 514226 597980 514294
rect -1916 514170 -1820 514226
rect -1764 514170 -1696 514226
rect -1640 514170 -1572 514226
rect -1516 514170 -1448 514226
rect -1392 514170 9234 514226
rect 9290 514170 9358 514226
rect 9414 514170 9482 514226
rect 9538 514170 9606 514226
rect 9662 514170 39954 514226
rect 40010 514170 40078 514226
rect 40134 514170 40202 514226
rect 40258 514170 40326 514226
rect 40382 514170 70674 514226
rect 70730 514170 70798 514226
rect 70854 514170 70922 514226
rect 70978 514170 71046 514226
rect 71102 514170 101394 514226
rect 101450 514170 101518 514226
rect 101574 514170 101642 514226
rect 101698 514170 101766 514226
rect 101822 514170 132114 514226
rect 132170 514170 132238 514226
rect 132294 514170 132362 514226
rect 132418 514170 132486 514226
rect 132542 514170 162834 514226
rect 162890 514170 162958 514226
rect 163014 514170 163082 514226
rect 163138 514170 163206 514226
rect 163262 514170 193554 514226
rect 193610 514170 193678 514226
rect 193734 514170 193802 514226
rect 193858 514170 193926 514226
rect 193982 514170 224274 514226
rect 224330 514170 224398 514226
rect 224454 514170 224522 514226
rect 224578 514170 224646 514226
rect 224702 514170 254994 514226
rect 255050 514170 255118 514226
rect 255174 514170 255242 514226
rect 255298 514170 255366 514226
rect 255422 514170 285714 514226
rect 285770 514170 285838 514226
rect 285894 514170 285962 514226
rect 286018 514170 286086 514226
rect 286142 514170 316434 514226
rect 316490 514170 316558 514226
rect 316614 514170 316682 514226
rect 316738 514170 316806 514226
rect 316862 514170 347154 514226
rect 347210 514170 347278 514226
rect 347334 514170 347402 514226
rect 347458 514170 347526 514226
rect 347582 514170 377874 514226
rect 377930 514170 377998 514226
rect 378054 514170 378122 514226
rect 378178 514170 378246 514226
rect 378302 514170 408594 514226
rect 408650 514170 408718 514226
rect 408774 514170 408842 514226
rect 408898 514170 408966 514226
rect 409022 514170 439314 514226
rect 439370 514170 439438 514226
rect 439494 514170 439562 514226
rect 439618 514170 439686 514226
rect 439742 514170 470034 514226
rect 470090 514170 470158 514226
rect 470214 514170 470282 514226
rect 470338 514170 470406 514226
rect 470462 514170 500754 514226
rect 500810 514170 500878 514226
rect 500934 514170 501002 514226
rect 501058 514170 501126 514226
rect 501182 514170 531474 514226
rect 531530 514170 531598 514226
rect 531654 514170 531722 514226
rect 531778 514170 531846 514226
rect 531902 514170 562194 514226
rect 562250 514170 562318 514226
rect 562374 514170 562442 514226
rect 562498 514170 562566 514226
rect 562622 514170 592914 514226
rect 592970 514170 593038 514226
rect 593094 514170 593162 514226
rect 593218 514170 593286 514226
rect 593342 514170 597456 514226
rect 597512 514170 597580 514226
rect 597636 514170 597704 514226
rect 597760 514170 597828 514226
rect 597884 514170 597980 514226
rect -1916 514102 597980 514170
rect -1916 514046 -1820 514102
rect -1764 514046 -1696 514102
rect -1640 514046 -1572 514102
rect -1516 514046 -1448 514102
rect -1392 514046 9234 514102
rect 9290 514046 9358 514102
rect 9414 514046 9482 514102
rect 9538 514046 9606 514102
rect 9662 514046 39954 514102
rect 40010 514046 40078 514102
rect 40134 514046 40202 514102
rect 40258 514046 40326 514102
rect 40382 514046 70674 514102
rect 70730 514046 70798 514102
rect 70854 514046 70922 514102
rect 70978 514046 71046 514102
rect 71102 514046 101394 514102
rect 101450 514046 101518 514102
rect 101574 514046 101642 514102
rect 101698 514046 101766 514102
rect 101822 514046 132114 514102
rect 132170 514046 132238 514102
rect 132294 514046 132362 514102
rect 132418 514046 132486 514102
rect 132542 514046 162834 514102
rect 162890 514046 162958 514102
rect 163014 514046 163082 514102
rect 163138 514046 163206 514102
rect 163262 514046 193554 514102
rect 193610 514046 193678 514102
rect 193734 514046 193802 514102
rect 193858 514046 193926 514102
rect 193982 514046 224274 514102
rect 224330 514046 224398 514102
rect 224454 514046 224522 514102
rect 224578 514046 224646 514102
rect 224702 514046 254994 514102
rect 255050 514046 255118 514102
rect 255174 514046 255242 514102
rect 255298 514046 255366 514102
rect 255422 514046 285714 514102
rect 285770 514046 285838 514102
rect 285894 514046 285962 514102
rect 286018 514046 286086 514102
rect 286142 514046 316434 514102
rect 316490 514046 316558 514102
rect 316614 514046 316682 514102
rect 316738 514046 316806 514102
rect 316862 514046 347154 514102
rect 347210 514046 347278 514102
rect 347334 514046 347402 514102
rect 347458 514046 347526 514102
rect 347582 514046 377874 514102
rect 377930 514046 377998 514102
rect 378054 514046 378122 514102
rect 378178 514046 378246 514102
rect 378302 514046 408594 514102
rect 408650 514046 408718 514102
rect 408774 514046 408842 514102
rect 408898 514046 408966 514102
rect 409022 514046 439314 514102
rect 439370 514046 439438 514102
rect 439494 514046 439562 514102
rect 439618 514046 439686 514102
rect 439742 514046 470034 514102
rect 470090 514046 470158 514102
rect 470214 514046 470282 514102
rect 470338 514046 470406 514102
rect 470462 514046 500754 514102
rect 500810 514046 500878 514102
rect 500934 514046 501002 514102
rect 501058 514046 501126 514102
rect 501182 514046 531474 514102
rect 531530 514046 531598 514102
rect 531654 514046 531722 514102
rect 531778 514046 531846 514102
rect 531902 514046 562194 514102
rect 562250 514046 562318 514102
rect 562374 514046 562442 514102
rect 562498 514046 562566 514102
rect 562622 514046 592914 514102
rect 592970 514046 593038 514102
rect 593094 514046 593162 514102
rect 593218 514046 593286 514102
rect 593342 514046 597456 514102
rect 597512 514046 597580 514102
rect 597636 514046 597704 514102
rect 597760 514046 597828 514102
rect 597884 514046 597980 514102
rect -1916 513978 597980 514046
rect -1916 513922 -1820 513978
rect -1764 513922 -1696 513978
rect -1640 513922 -1572 513978
rect -1516 513922 -1448 513978
rect -1392 513922 9234 513978
rect 9290 513922 9358 513978
rect 9414 513922 9482 513978
rect 9538 513922 9606 513978
rect 9662 513922 39954 513978
rect 40010 513922 40078 513978
rect 40134 513922 40202 513978
rect 40258 513922 40326 513978
rect 40382 513922 70674 513978
rect 70730 513922 70798 513978
rect 70854 513922 70922 513978
rect 70978 513922 71046 513978
rect 71102 513922 101394 513978
rect 101450 513922 101518 513978
rect 101574 513922 101642 513978
rect 101698 513922 101766 513978
rect 101822 513922 132114 513978
rect 132170 513922 132238 513978
rect 132294 513922 132362 513978
rect 132418 513922 132486 513978
rect 132542 513922 162834 513978
rect 162890 513922 162958 513978
rect 163014 513922 163082 513978
rect 163138 513922 163206 513978
rect 163262 513922 193554 513978
rect 193610 513922 193678 513978
rect 193734 513922 193802 513978
rect 193858 513922 193926 513978
rect 193982 513922 224274 513978
rect 224330 513922 224398 513978
rect 224454 513922 224522 513978
rect 224578 513922 224646 513978
rect 224702 513922 254994 513978
rect 255050 513922 255118 513978
rect 255174 513922 255242 513978
rect 255298 513922 255366 513978
rect 255422 513922 285714 513978
rect 285770 513922 285838 513978
rect 285894 513922 285962 513978
rect 286018 513922 286086 513978
rect 286142 513922 316434 513978
rect 316490 513922 316558 513978
rect 316614 513922 316682 513978
rect 316738 513922 316806 513978
rect 316862 513922 347154 513978
rect 347210 513922 347278 513978
rect 347334 513922 347402 513978
rect 347458 513922 347526 513978
rect 347582 513922 377874 513978
rect 377930 513922 377998 513978
rect 378054 513922 378122 513978
rect 378178 513922 378246 513978
rect 378302 513922 408594 513978
rect 408650 513922 408718 513978
rect 408774 513922 408842 513978
rect 408898 513922 408966 513978
rect 409022 513922 439314 513978
rect 439370 513922 439438 513978
rect 439494 513922 439562 513978
rect 439618 513922 439686 513978
rect 439742 513922 470034 513978
rect 470090 513922 470158 513978
rect 470214 513922 470282 513978
rect 470338 513922 470406 513978
rect 470462 513922 500754 513978
rect 500810 513922 500878 513978
rect 500934 513922 501002 513978
rect 501058 513922 501126 513978
rect 501182 513922 531474 513978
rect 531530 513922 531598 513978
rect 531654 513922 531722 513978
rect 531778 513922 531846 513978
rect 531902 513922 562194 513978
rect 562250 513922 562318 513978
rect 562374 513922 562442 513978
rect 562498 513922 562566 513978
rect 562622 513922 592914 513978
rect 592970 513922 593038 513978
rect 593094 513922 593162 513978
rect 593218 513922 593286 513978
rect 593342 513922 597456 513978
rect 597512 513922 597580 513978
rect 597636 513922 597704 513978
rect 597760 513922 597828 513978
rect 597884 513922 597980 513978
rect -1916 513826 597980 513922
rect -1916 508350 597980 508446
rect -1916 508294 -860 508350
rect -804 508294 -736 508350
rect -680 508294 -612 508350
rect -556 508294 -488 508350
rect -432 508294 5514 508350
rect 5570 508294 5638 508350
rect 5694 508294 5762 508350
rect 5818 508294 5886 508350
rect 5942 508294 36234 508350
rect 36290 508294 36358 508350
rect 36414 508294 36482 508350
rect 36538 508294 36606 508350
rect 36662 508294 66954 508350
rect 67010 508294 67078 508350
rect 67134 508294 67202 508350
rect 67258 508294 67326 508350
rect 67382 508294 97674 508350
rect 97730 508294 97798 508350
rect 97854 508294 97922 508350
rect 97978 508294 98046 508350
rect 98102 508294 128394 508350
rect 128450 508294 128518 508350
rect 128574 508294 128642 508350
rect 128698 508294 128766 508350
rect 128822 508294 159114 508350
rect 159170 508294 159238 508350
rect 159294 508294 159362 508350
rect 159418 508294 159486 508350
rect 159542 508294 189834 508350
rect 189890 508294 189958 508350
rect 190014 508294 190082 508350
rect 190138 508294 190206 508350
rect 190262 508294 220554 508350
rect 220610 508294 220678 508350
rect 220734 508294 220802 508350
rect 220858 508294 220926 508350
rect 220982 508294 251274 508350
rect 251330 508294 251398 508350
rect 251454 508294 251522 508350
rect 251578 508294 251646 508350
rect 251702 508294 281994 508350
rect 282050 508294 282118 508350
rect 282174 508294 282242 508350
rect 282298 508294 282366 508350
rect 282422 508294 312714 508350
rect 312770 508294 312838 508350
rect 312894 508294 312962 508350
rect 313018 508294 313086 508350
rect 313142 508294 343434 508350
rect 343490 508294 343558 508350
rect 343614 508294 343682 508350
rect 343738 508294 343806 508350
rect 343862 508294 374154 508350
rect 374210 508294 374278 508350
rect 374334 508294 374402 508350
rect 374458 508294 374526 508350
rect 374582 508294 404874 508350
rect 404930 508294 404998 508350
rect 405054 508294 405122 508350
rect 405178 508294 405246 508350
rect 405302 508294 435594 508350
rect 435650 508294 435718 508350
rect 435774 508294 435842 508350
rect 435898 508294 435966 508350
rect 436022 508294 466314 508350
rect 466370 508294 466438 508350
rect 466494 508294 466562 508350
rect 466618 508294 466686 508350
rect 466742 508294 497034 508350
rect 497090 508294 497158 508350
rect 497214 508294 497282 508350
rect 497338 508294 497406 508350
rect 497462 508294 527754 508350
rect 527810 508294 527878 508350
rect 527934 508294 528002 508350
rect 528058 508294 528126 508350
rect 528182 508294 558474 508350
rect 558530 508294 558598 508350
rect 558654 508294 558722 508350
rect 558778 508294 558846 508350
rect 558902 508294 589194 508350
rect 589250 508294 589318 508350
rect 589374 508294 589442 508350
rect 589498 508294 589566 508350
rect 589622 508294 596496 508350
rect 596552 508294 596620 508350
rect 596676 508294 596744 508350
rect 596800 508294 596868 508350
rect 596924 508294 597980 508350
rect -1916 508226 597980 508294
rect -1916 508170 -860 508226
rect -804 508170 -736 508226
rect -680 508170 -612 508226
rect -556 508170 -488 508226
rect -432 508170 5514 508226
rect 5570 508170 5638 508226
rect 5694 508170 5762 508226
rect 5818 508170 5886 508226
rect 5942 508170 36234 508226
rect 36290 508170 36358 508226
rect 36414 508170 36482 508226
rect 36538 508170 36606 508226
rect 36662 508170 66954 508226
rect 67010 508170 67078 508226
rect 67134 508170 67202 508226
rect 67258 508170 67326 508226
rect 67382 508170 97674 508226
rect 97730 508170 97798 508226
rect 97854 508170 97922 508226
rect 97978 508170 98046 508226
rect 98102 508170 128394 508226
rect 128450 508170 128518 508226
rect 128574 508170 128642 508226
rect 128698 508170 128766 508226
rect 128822 508170 159114 508226
rect 159170 508170 159238 508226
rect 159294 508170 159362 508226
rect 159418 508170 159486 508226
rect 159542 508170 189834 508226
rect 189890 508170 189958 508226
rect 190014 508170 190082 508226
rect 190138 508170 190206 508226
rect 190262 508170 220554 508226
rect 220610 508170 220678 508226
rect 220734 508170 220802 508226
rect 220858 508170 220926 508226
rect 220982 508170 251274 508226
rect 251330 508170 251398 508226
rect 251454 508170 251522 508226
rect 251578 508170 251646 508226
rect 251702 508170 281994 508226
rect 282050 508170 282118 508226
rect 282174 508170 282242 508226
rect 282298 508170 282366 508226
rect 282422 508170 312714 508226
rect 312770 508170 312838 508226
rect 312894 508170 312962 508226
rect 313018 508170 313086 508226
rect 313142 508170 343434 508226
rect 343490 508170 343558 508226
rect 343614 508170 343682 508226
rect 343738 508170 343806 508226
rect 343862 508170 374154 508226
rect 374210 508170 374278 508226
rect 374334 508170 374402 508226
rect 374458 508170 374526 508226
rect 374582 508170 404874 508226
rect 404930 508170 404998 508226
rect 405054 508170 405122 508226
rect 405178 508170 405246 508226
rect 405302 508170 435594 508226
rect 435650 508170 435718 508226
rect 435774 508170 435842 508226
rect 435898 508170 435966 508226
rect 436022 508170 466314 508226
rect 466370 508170 466438 508226
rect 466494 508170 466562 508226
rect 466618 508170 466686 508226
rect 466742 508170 497034 508226
rect 497090 508170 497158 508226
rect 497214 508170 497282 508226
rect 497338 508170 497406 508226
rect 497462 508170 527754 508226
rect 527810 508170 527878 508226
rect 527934 508170 528002 508226
rect 528058 508170 528126 508226
rect 528182 508170 558474 508226
rect 558530 508170 558598 508226
rect 558654 508170 558722 508226
rect 558778 508170 558846 508226
rect 558902 508170 589194 508226
rect 589250 508170 589318 508226
rect 589374 508170 589442 508226
rect 589498 508170 589566 508226
rect 589622 508170 596496 508226
rect 596552 508170 596620 508226
rect 596676 508170 596744 508226
rect 596800 508170 596868 508226
rect 596924 508170 597980 508226
rect -1916 508102 597980 508170
rect -1916 508046 -860 508102
rect -804 508046 -736 508102
rect -680 508046 -612 508102
rect -556 508046 -488 508102
rect -432 508046 5514 508102
rect 5570 508046 5638 508102
rect 5694 508046 5762 508102
rect 5818 508046 5886 508102
rect 5942 508046 36234 508102
rect 36290 508046 36358 508102
rect 36414 508046 36482 508102
rect 36538 508046 36606 508102
rect 36662 508046 66954 508102
rect 67010 508046 67078 508102
rect 67134 508046 67202 508102
rect 67258 508046 67326 508102
rect 67382 508046 97674 508102
rect 97730 508046 97798 508102
rect 97854 508046 97922 508102
rect 97978 508046 98046 508102
rect 98102 508046 128394 508102
rect 128450 508046 128518 508102
rect 128574 508046 128642 508102
rect 128698 508046 128766 508102
rect 128822 508046 159114 508102
rect 159170 508046 159238 508102
rect 159294 508046 159362 508102
rect 159418 508046 159486 508102
rect 159542 508046 189834 508102
rect 189890 508046 189958 508102
rect 190014 508046 190082 508102
rect 190138 508046 190206 508102
rect 190262 508046 220554 508102
rect 220610 508046 220678 508102
rect 220734 508046 220802 508102
rect 220858 508046 220926 508102
rect 220982 508046 251274 508102
rect 251330 508046 251398 508102
rect 251454 508046 251522 508102
rect 251578 508046 251646 508102
rect 251702 508046 281994 508102
rect 282050 508046 282118 508102
rect 282174 508046 282242 508102
rect 282298 508046 282366 508102
rect 282422 508046 312714 508102
rect 312770 508046 312838 508102
rect 312894 508046 312962 508102
rect 313018 508046 313086 508102
rect 313142 508046 343434 508102
rect 343490 508046 343558 508102
rect 343614 508046 343682 508102
rect 343738 508046 343806 508102
rect 343862 508046 374154 508102
rect 374210 508046 374278 508102
rect 374334 508046 374402 508102
rect 374458 508046 374526 508102
rect 374582 508046 404874 508102
rect 404930 508046 404998 508102
rect 405054 508046 405122 508102
rect 405178 508046 405246 508102
rect 405302 508046 435594 508102
rect 435650 508046 435718 508102
rect 435774 508046 435842 508102
rect 435898 508046 435966 508102
rect 436022 508046 466314 508102
rect 466370 508046 466438 508102
rect 466494 508046 466562 508102
rect 466618 508046 466686 508102
rect 466742 508046 497034 508102
rect 497090 508046 497158 508102
rect 497214 508046 497282 508102
rect 497338 508046 497406 508102
rect 497462 508046 527754 508102
rect 527810 508046 527878 508102
rect 527934 508046 528002 508102
rect 528058 508046 528126 508102
rect 528182 508046 558474 508102
rect 558530 508046 558598 508102
rect 558654 508046 558722 508102
rect 558778 508046 558846 508102
rect 558902 508046 589194 508102
rect 589250 508046 589318 508102
rect 589374 508046 589442 508102
rect 589498 508046 589566 508102
rect 589622 508046 596496 508102
rect 596552 508046 596620 508102
rect 596676 508046 596744 508102
rect 596800 508046 596868 508102
rect 596924 508046 597980 508102
rect -1916 507978 597980 508046
rect -1916 507922 -860 507978
rect -804 507922 -736 507978
rect -680 507922 -612 507978
rect -556 507922 -488 507978
rect -432 507922 5514 507978
rect 5570 507922 5638 507978
rect 5694 507922 5762 507978
rect 5818 507922 5886 507978
rect 5942 507922 36234 507978
rect 36290 507922 36358 507978
rect 36414 507922 36482 507978
rect 36538 507922 36606 507978
rect 36662 507922 66954 507978
rect 67010 507922 67078 507978
rect 67134 507922 67202 507978
rect 67258 507922 67326 507978
rect 67382 507922 97674 507978
rect 97730 507922 97798 507978
rect 97854 507922 97922 507978
rect 97978 507922 98046 507978
rect 98102 507922 128394 507978
rect 128450 507922 128518 507978
rect 128574 507922 128642 507978
rect 128698 507922 128766 507978
rect 128822 507922 159114 507978
rect 159170 507922 159238 507978
rect 159294 507922 159362 507978
rect 159418 507922 159486 507978
rect 159542 507922 189834 507978
rect 189890 507922 189958 507978
rect 190014 507922 190082 507978
rect 190138 507922 190206 507978
rect 190262 507922 220554 507978
rect 220610 507922 220678 507978
rect 220734 507922 220802 507978
rect 220858 507922 220926 507978
rect 220982 507922 251274 507978
rect 251330 507922 251398 507978
rect 251454 507922 251522 507978
rect 251578 507922 251646 507978
rect 251702 507922 281994 507978
rect 282050 507922 282118 507978
rect 282174 507922 282242 507978
rect 282298 507922 282366 507978
rect 282422 507922 312714 507978
rect 312770 507922 312838 507978
rect 312894 507922 312962 507978
rect 313018 507922 313086 507978
rect 313142 507922 343434 507978
rect 343490 507922 343558 507978
rect 343614 507922 343682 507978
rect 343738 507922 343806 507978
rect 343862 507922 374154 507978
rect 374210 507922 374278 507978
rect 374334 507922 374402 507978
rect 374458 507922 374526 507978
rect 374582 507922 404874 507978
rect 404930 507922 404998 507978
rect 405054 507922 405122 507978
rect 405178 507922 405246 507978
rect 405302 507922 435594 507978
rect 435650 507922 435718 507978
rect 435774 507922 435842 507978
rect 435898 507922 435966 507978
rect 436022 507922 466314 507978
rect 466370 507922 466438 507978
rect 466494 507922 466562 507978
rect 466618 507922 466686 507978
rect 466742 507922 497034 507978
rect 497090 507922 497158 507978
rect 497214 507922 497282 507978
rect 497338 507922 497406 507978
rect 497462 507922 527754 507978
rect 527810 507922 527878 507978
rect 527934 507922 528002 507978
rect 528058 507922 528126 507978
rect 528182 507922 558474 507978
rect 558530 507922 558598 507978
rect 558654 507922 558722 507978
rect 558778 507922 558846 507978
rect 558902 507922 589194 507978
rect 589250 507922 589318 507978
rect 589374 507922 589442 507978
rect 589498 507922 589566 507978
rect 589622 507922 596496 507978
rect 596552 507922 596620 507978
rect 596676 507922 596744 507978
rect 596800 507922 596868 507978
rect 596924 507922 597980 507978
rect -1916 507826 597980 507922
rect -1916 496350 597980 496446
rect -1916 496294 -1820 496350
rect -1764 496294 -1696 496350
rect -1640 496294 -1572 496350
rect -1516 496294 -1448 496350
rect -1392 496294 9234 496350
rect 9290 496294 9358 496350
rect 9414 496294 9482 496350
rect 9538 496294 9606 496350
rect 9662 496294 39954 496350
rect 40010 496294 40078 496350
rect 40134 496294 40202 496350
rect 40258 496294 40326 496350
rect 40382 496294 70674 496350
rect 70730 496294 70798 496350
rect 70854 496294 70922 496350
rect 70978 496294 71046 496350
rect 71102 496294 101394 496350
rect 101450 496294 101518 496350
rect 101574 496294 101642 496350
rect 101698 496294 101766 496350
rect 101822 496294 132114 496350
rect 132170 496294 132238 496350
rect 132294 496294 132362 496350
rect 132418 496294 132486 496350
rect 132542 496294 162834 496350
rect 162890 496294 162958 496350
rect 163014 496294 163082 496350
rect 163138 496294 163206 496350
rect 163262 496294 193554 496350
rect 193610 496294 193678 496350
rect 193734 496294 193802 496350
rect 193858 496294 193926 496350
rect 193982 496294 224274 496350
rect 224330 496294 224398 496350
rect 224454 496294 224522 496350
rect 224578 496294 224646 496350
rect 224702 496294 254994 496350
rect 255050 496294 255118 496350
rect 255174 496294 255242 496350
rect 255298 496294 255366 496350
rect 255422 496294 285714 496350
rect 285770 496294 285838 496350
rect 285894 496294 285962 496350
rect 286018 496294 286086 496350
rect 286142 496294 316434 496350
rect 316490 496294 316558 496350
rect 316614 496294 316682 496350
rect 316738 496294 316806 496350
rect 316862 496294 347154 496350
rect 347210 496294 347278 496350
rect 347334 496294 347402 496350
rect 347458 496294 347526 496350
rect 347582 496294 377874 496350
rect 377930 496294 377998 496350
rect 378054 496294 378122 496350
rect 378178 496294 378246 496350
rect 378302 496294 408594 496350
rect 408650 496294 408718 496350
rect 408774 496294 408842 496350
rect 408898 496294 408966 496350
rect 409022 496294 439314 496350
rect 439370 496294 439438 496350
rect 439494 496294 439562 496350
rect 439618 496294 439686 496350
rect 439742 496294 470034 496350
rect 470090 496294 470158 496350
rect 470214 496294 470282 496350
rect 470338 496294 470406 496350
rect 470462 496294 500754 496350
rect 500810 496294 500878 496350
rect 500934 496294 501002 496350
rect 501058 496294 501126 496350
rect 501182 496294 531474 496350
rect 531530 496294 531598 496350
rect 531654 496294 531722 496350
rect 531778 496294 531846 496350
rect 531902 496294 562194 496350
rect 562250 496294 562318 496350
rect 562374 496294 562442 496350
rect 562498 496294 562566 496350
rect 562622 496294 592914 496350
rect 592970 496294 593038 496350
rect 593094 496294 593162 496350
rect 593218 496294 593286 496350
rect 593342 496294 597456 496350
rect 597512 496294 597580 496350
rect 597636 496294 597704 496350
rect 597760 496294 597828 496350
rect 597884 496294 597980 496350
rect -1916 496226 597980 496294
rect -1916 496170 -1820 496226
rect -1764 496170 -1696 496226
rect -1640 496170 -1572 496226
rect -1516 496170 -1448 496226
rect -1392 496170 9234 496226
rect 9290 496170 9358 496226
rect 9414 496170 9482 496226
rect 9538 496170 9606 496226
rect 9662 496170 39954 496226
rect 40010 496170 40078 496226
rect 40134 496170 40202 496226
rect 40258 496170 40326 496226
rect 40382 496170 70674 496226
rect 70730 496170 70798 496226
rect 70854 496170 70922 496226
rect 70978 496170 71046 496226
rect 71102 496170 101394 496226
rect 101450 496170 101518 496226
rect 101574 496170 101642 496226
rect 101698 496170 101766 496226
rect 101822 496170 132114 496226
rect 132170 496170 132238 496226
rect 132294 496170 132362 496226
rect 132418 496170 132486 496226
rect 132542 496170 162834 496226
rect 162890 496170 162958 496226
rect 163014 496170 163082 496226
rect 163138 496170 163206 496226
rect 163262 496170 193554 496226
rect 193610 496170 193678 496226
rect 193734 496170 193802 496226
rect 193858 496170 193926 496226
rect 193982 496170 224274 496226
rect 224330 496170 224398 496226
rect 224454 496170 224522 496226
rect 224578 496170 224646 496226
rect 224702 496170 254994 496226
rect 255050 496170 255118 496226
rect 255174 496170 255242 496226
rect 255298 496170 255366 496226
rect 255422 496170 285714 496226
rect 285770 496170 285838 496226
rect 285894 496170 285962 496226
rect 286018 496170 286086 496226
rect 286142 496170 316434 496226
rect 316490 496170 316558 496226
rect 316614 496170 316682 496226
rect 316738 496170 316806 496226
rect 316862 496170 347154 496226
rect 347210 496170 347278 496226
rect 347334 496170 347402 496226
rect 347458 496170 347526 496226
rect 347582 496170 377874 496226
rect 377930 496170 377998 496226
rect 378054 496170 378122 496226
rect 378178 496170 378246 496226
rect 378302 496170 408594 496226
rect 408650 496170 408718 496226
rect 408774 496170 408842 496226
rect 408898 496170 408966 496226
rect 409022 496170 439314 496226
rect 439370 496170 439438 496226
rect 439494 496170 439562 496226
rect 439618 496170 439686 496226
rect 439742 496170 470034 496226
rect 470090 496170 470158 496226
rect 470214 496170 470282 496226
rect 470338 496170 470406 496226
rect 470462 496170 500754 496226
rect 500810 496170 500878 496226
rect 500934 496170 501002 496226
rect 501058 496170 501126 496226
rect 501182 496170 531474 496226
rect 531530 496170 531598 496226
rect 531654 496170 531722 496226
rect 531778 496170 531846 496226
rect 531902 496170 562194 496226
rect 562250 496170 562318 496226
rect 562374 496170 562442 496226
rect 562498 496170 562566 496226
rect 562622 496170 592914 496226
rect 592970 496170 593038 496226
rect 593094 496170 593162 496226
rect 593218 496170 593286 496226
rect 593342 496170 597456 496226
rect 597512 496170 597580 496226
rect 597636 496170 597704 496226
rect 597760 496170 597828 496226
rect 597884 496170 597980 496226
rect -1916 496102 597980 496170
rect -1916 496046 -1820 496102
rect -1764 496046 -1696 496102
rect -1640 496046 -1572 496102
rect -1516 496046 -1448 496102
rect -1392 496046 9234 496102
rect 9290 496046 9358 496102
rect 9414 496046 9482 496102
rect 9538 496046 9606 496102
rect 9662 496046 39954 496102
rect 40010 496046 40078 496102
rect 40134 496046 40202 496102
rect 40258 496046 40326 496102
rect 40382 496046 70674 496102
rect 70730 496046 70798 496102
rect 70854 496046 70922 496102
rect 70978 496046 71046 496102
rect 71102 496046 101394 496102
rect 101450 496046 101518 496102
rect 101574 496046 101642 496102
rect 101698 496046 101766 496102
rect 101822 496046 132114 496102
rect 132170 496046 132238 496102
rect 132294 496046 132362 496102
rect 132418 496046 132486 496102
rect 132542 496046 162834 496102
rect 162890 496046 162958 496102
rect 163014 496046 163082 496102
rect 163138 496046 163206 496102
rect 163262 496046 193554 496102
rect 193610 496046 193678 496102
rect 193734 496046 193802 496102
rect 193858 496046 193926 496102
rect 193982 496046 224274 496102
rect 224330 496046 224398 496102
rect 224454 496046 224522 496102
rect 224578 496046 224646 496102
rect 224702 496046 254994 496102
rect 255050 496046 255118 496102
rect 255174 496046 255242 496102
rect 255298 496046 255366 496102
rect 255422 496046 285714 496102
rect 285770 496046 285838 496102
rect 285894 496046 285962 496102
rect 286018 496046 286086 496102
rect 286142 496046 316434 496102
rect 316490 496046 316558 496102
rect 316614 496046 316682 496102
rect 316738 496046 316806 496102
rect 316862 496046 347154 496102
rect 347210 496046 347278 496102
rect 347334 496046 347402 496102
rect 347458 496046 347526 496102
rect 347582 496046 377874 496102
rect 377930 496046 377998 496102
rect 378054 496046 378122 496102
rect 378178 496046 378246 496102
rect 378302 496046 408594 496102
rect 408650 496046 408718 496102
rect 408774 496046 408842 496102
rect 408898 496046 408966 496102
rect 409022 496046 439314 496102
rect 439370 496046 439438 496102
rect 439494 496046 439562 496102
rect 439618 496046 439686 496102
rect 439742 496046 470034 496102
rect 470090 496046 470158 496102
rect 470214 496046 470282 496102
rect 470338 496046 470406 496102
rect 470462 496046 500754 496102
rect 500810 496046 500878 496102
rect 500934 496046 501002 496102
rect 501058 496046 501126 496102
rect 501182 496046 531474 496102
rect 531530 496046 531598 496102
rect 531654 496046 531722 496102
rect 531778 496046 531846 496102
rect 531902 496046 562194 496102
rect 562250 496046 562318 496102
rect 562374 496046 562442 496102
rect 562498 496046 562566 496102
rect 562622 496046 592914 496102
rect 592970 496046 593038 496102
rect 593094 496046 593162 496102
rect 593218 496046 593286 496102
rect 593342 496046 597456 496102
rect 597512 496046 597580 496102
rect 597636 496046 597704 496102
rect 597760 496046 597828 496102
rect 597884 496046 597980 496102
rect -1916 495978 597980 496046
rect -1916 495922 -1820 495978
rect -1764 495922 -1696 495978
rect -1640 495922 -1572 495978
rect -1516 495922 -1448 495978
rect -1392 495922 9234 495978
rect 9290 495922 9358 495978
rect 9414 495922 9482 495978
rect 9538 495922 9606 495978
rect 9662 495922 39954 495978
rect 40010 495922 40078 495978
rect 40134 495922 40202 495978
rect 40258 495922 40326 495978
rect 40382 495922 70674 495978
rect 70730 495922 70798 495978
rect 70854 495922 70922 495978
rect 70978 495922 71046 495978
rect 71102 495922 101394 495978
rect 101450 495922 101518 495978
rect 101574 495922 101642 495978
rect 101698 495922 101766 495978
rect 101822 495922 132114 495978
rect 132170 495922 132238 495978
rect 132294 495922 132362 495978
rect 132418 495922 132486 495978
rect 132542 495922 162834 495978
rect 162890 495922 162958 495978
rect 163014 495922 163082 495978
rect 163138 495922 163206 495978
rect 163262 495922 193554 495978
rect 193610 495922 193678 495978
rect 193734 495922 193802 495978
rect 193858 495922 193926 495978
rect 193982 495922 224274 495978
rect 224330 495922 224398 495978
rect 224454 495922 224522 495978
rect 224578 495922 224646 495978
rect 224702 495922 254994 495978
rect 255050 495922 255118 495978
rect 255174 495922 255242 495978
rect 255298 495922 255366 495978
rect 255422 495922 285714 495978
rect 285770 495922 285838 495978
rect 285894 495922 285962 495978
rect 286018 495922 286086 495978
rect 286142 495922 316434 495978
rect 316490 495922 316558 495978
rect 316614 495922 316682 495978
rect 316738 495922 316806 495978
rect 316862 495922 347154 495978
rect 347210 495922 347278 495978
rect 347334 495922 347402 495978
rect 347458 495922 347526 495978
rect 347582 495922 377874 495978
rect 377930 495922 377998 495978
rect 378054 495922 378122 495978
rect 378178 495922 378246 495978
rect 378302 495922 408594 495978
rect 408650 495922 408718 495978
rect 408774 495922 408842 495978
rect 408898 495922 408966 495978
rect 409022 495922 439314 495978
rect 439370 495922 439438 495978
rect 439494 495922 439562 495978
rect 439618 495922 439686 495978
rect 439742 495922 470034 495978
rect 470090 495922 470158 495978
rect 470214 495922 470282 495978
rect 470338 495922 470406 495978
rect 470462 495922 500754 495978
rect 500810 495922 500878 495978
rect 500934 495922 501002 495978
rect 501058 495922 501126 495978
rect 501182 495922 531474 495978
rect 531530 495922 531598 495978
rect 531654 495922 531722 495978
rect 531778 495922 531846 495978
rect 531902 495922 562194 495978
rect 562250 495922 562318 495978
rect 562374 495922 562442 495978
rect 562498 495922 562566 495978
rect 562622 495922 592914 495978
rect 592970 495922 593038 495978
rect 593094 495922 593162 495978
rect 593218 495922 593286 495978
rect 593342 495922 597456 495978
rect 597512 495922 597580 495978
rect 597636 495922 597704 495978
rect 597760 495922 597828 495978
rect 597884 495922 597980 495978
rect -1916 495826 597980 495922
rect -1916 490350 597980 490446
rect -1916 490294 -860 490350
rect -804 490294 -736 490350
rect -680 490294 -612 490350
rect -556 490294 -488 490350
rect -432 490294 5514 490350
rect 5570 490294 5638 490350
rect 5694 490294 5762 490350
rect 5818 490294 5886 490350
rect 5942 490294 36234 490350
rect 36290 490294 36358 490350
rect 36414 490294 36482 490350
rect 36538 490294 36606 490350
rect 36662 490294 66954 490350
rect 67010 490294 67078 490350
rect 67134 490294 67202 490350
rect 67258 490294 67326 490350
rect 67382 490294 97674 490350
rect 97730 490294 97798 490350
rect 97854 490294 97922 490350
rect 97978 490294 98046 490350
rect 98102 490294 128394 490350
rect 128450 490294 128518 490350
rect 128574 490294 128642 490350
rect 128698 490294 128766 490350
rect 128822 490294 159114 490350
rect 159170 490294 159238 490350
rect 159294 490294 159362 490350
rect 159418 490294 159486 490350
rect 159542 490294 189834 490350
rect 189890 490294 189958 490350
rect 190014 490294 190082 490350
rect 190138 490294 190206 490350
rect 190262 490294 220554 490350
rect 220610 490294 220678 490350
rect 220734 490294 220802 490350
rect 220858 490294 220926 490350
rect 220982 490294 251274 490350
rect 251330 490294 251398 490350
rect 251454 490294 251522 490350
rect 251578 490294 251646 490350
rect 251702 490294 281994 490350
rect 282050 490294 282118 490350
rect 282174 490294 282242 490350
rect 282298 490294 282366 490350
rect 282422 490294 312714 490350
rect 312770 490294 312838 490350
rect 312894 490294 312962 490350
rect 313018 490294 313086 490350
rect 313142 490294 343434 490350
rect 343490 490294 343558 490350
rect 343614 490294 343682 490350
rect 343738 490294 343806 490350
rect 343862 490294 374154 490350
rect 374210 490294 374278 490350
rect 374334 490294 374402 490350
rect 374458 490294 374526 490350
rect 374582 490294 404874 490350
rect 404930 490294 404998 490350
rect 405054 490294 405122 490350
rect 405178 490294 405246 490350
rect 405302 490294 435594 490350
rect 435650 490294 435718 490350
rect 435774 490294 435842 490350
rect 435898 490294 435966 490350
rect 436022 490294 466314 490350
rect 466370 490294 466438 490350
rect 466494 490294 466562 490350
rect 466618 490294 466686 490350
rect 466742 490294 497034 490350
rect 497090 490294 497158 490350
rect 497214 490294 497282 490350
rect 497338 490294 497406 490350
rect 497462 490294 527754 490350
rect 527810 490294 527878 490350
rect 527934 490294 528002 490350
rect 528058 490294 528126 490350
rect 528182 490294 558474 490350
rect 558530 490294 558598 490350
rect 558654 490294 558722 490350
rect 558778 490294 558846 490350
rect 558902 490294 589194 490350
rect 589250 490294 589318 490350
rect 589374 490294 589442 490350
rect 589498 490294 589566 490350
rect 589622 490294 596496 490350
rect 596552 490294 596620 490350
rect 596676 490294 596744 490350
rect 596800 490294 596868 490350
rect 596924 490294 597980 490350
rect -1916 490226 597980 490294
rect -1916 490170 -860 490226
rect -804 490170 -736 490226
rect -680 490170 -612 490226
rect -556 490170 -488 490226
rect -432 490170 5514 490226
rect 5570 490170 5638 490226
rect 5694 490170 5762 490226
rect 5818 490170 5886 490226
rect 5942 490170 36234 490226
rect 36290 490170 36358 490226
rect 36414 490170 36482 490226
rect 36538 490170 36606 490226
rect 36662 490170 66954 490226
rect 67010 490170 67078 490226
rect 67134 490170 67202 490226
rect 67258 490170 67326 490226
rect 67382 490170 97674 490226
rect 97730 490170 97798 490226
rect 97854 490170 97922 490226
rect 97978 490170 98046 490226
rect 98102 490170 128394 490226
rect 128450 490170 128518 490226
rect 128574 490170 128642 490226
rect 128698 490170 128766 490226
rect 128822 490170 159114 490226
rect 159170 490170 159238 490226
rect 159294 490170 159362 490226
rect 159418 490170 159486 490226
rect 159542 490170 189834 490226
rect 189890 490170 189958 490226
rect 190014 490170 190082 490226
rect 190138 490170 190206 490226
rect 190262 490170 220554 490226
rect 220610 490170 220678 490226
rect 220734 490170 220802 490226
rect 220858 490170 220926 490226
rect 220982 490170 251274 490226
rect 251330 490170 251398 490226
rect 251454 490170 251522 490226
rect 251578 490170 251646 490226
rect 251702 490170 281994 490226
rect 282050 490170 282118 490226
rect 282174 490170 282242 490226
rect 282298 490170 282366 490226
rect 282422 490170 312714 490226
rect 312770 490170 312838 490226
rect 312894 490170 312962 490226
rect 313018 490170 313086 490226
rect 313142 490170 343434 490226
rect 343490 490170 343558 490226
rect 343614 490170 343682 490226
rect 343738 490170 343806 490226
rect 343862 490170 374154 490226
rect 374210 490170 374278 490226
rect 374334 490170 374402 490226
rect 374458 490170 374526 490226
rect 374582 490170 404874 490226
rect 404930 490170 404998 490226
rect 405054 490170 405122 490226
rect 405178 490170 405246 490226
rect 405302 490170 435594 490226
rect 435650 490170 435718 490226
rect 435774 490170 435842 490226
rect 435898 490170 435966 490226
rect 436022 490170 466314 490226
rect 466370 490170 466438 490226
rect 466494 490170 466562 490226
rect 466618 490170 466686 490226
rect 466742 490170 497034 490226
rect 497090 490170 497158 490226
rect 497214 490170 497282 490226
rect 497338 490170 497406 490226
rect 497462 490170 527754 490226
rect 527810 490170 527878 490226
rect 527934 490170 528002 490226
rect 528058 490170 528126 490226
rect 528182 490170 558474 490226
rect 558530 490170 558598 490226
rect 558654 490170 558722 490226
rect 558778 490170 558846 490226
rect 558902 490170 589194 490226
rect 589250 490170 589318 490226
rect 589374 490170 589442 490226
rect 589498 490170 589566 490226
rect 589622 490170 596496 490226
rect 596552 490170 596620 490226
rect 596676 490170 596744 490226
rect 596800 490170 596868 490226
rect 596924 490170 597980 490226
rect -1916 490102 597980 490170
rect -1916 490046 -860 490102
rect -804 490046 -736 490102
rect -680 490046 -612 490102
rect -556 490046 -488 490102
rect -432 490046 5514 490102
rect 5570 490046 5638 490102
rect 5694 490046 5762 490102
rect 5818 490046 5886 490102
rect 5942 490046 36234 490102
rect 36290 490046 36358 490102
rect 36414 490046 36482 490102
rect 36538 490046 36606 490102
rect 36662 490046 66954 490102
rect 67010 490046 67078 490102
rect 67134 490046 67202 490102
rect 67258 490046 67326 490102
rect 67382 490046 97674 490102
rect 97730 490046 97798 490102
rect 97854 490046 97922 490102
rect 97978 490046 98046 490102
rect 98102 490046 128394 490102
rect 128450 490046 128518 490102
rect 128574 490046 128642 490102
rect 128698 490046 128766 490102
rect 128822 490046 159114 490102
rect 159170 490046 159238 490102
rect 159294 490046 159362 490102
rect 159418 490046 159486 490102
rect 159542 490046 189834 490102
rect 189890 490046 189958 490102
rect 190014 490046 190082 490102
rect 190138 490046 190206 490102
rect 190262 490046 220554 490102
rect 220610 490046 220678 490102
rect 220734 490046 220802 490102
rect 220858 490046 220926 490102
rect 220982 490046 251274 490102
rect 251330 490046 251398 490102
rect 251454 490046 251522 490102
rect 251578 490046 251646 490102
rect 251702 490046 281994 490102
rect 282050 490046 282118 490102
rect 282174 490046 282242 490102
rect 282298 490046 282366 490102
rect 282422 490046 312714 490102
rect 312770 490046 312838 490102
rect 312894 490046 312962 490102
rect 313018 490046 313086 490102
rect 313142 490046 343434 490102
rect 343490 490046 343558 490102
rect 343614 490046 343682 490102
rect 343738 490046 343806 490102
rect 343862 490046 374154 490102
rect 374210 490046 374278 490102
rect 374334 490046 374402 490102
rect 374458 490046 374526 490102
rect 374582 490046 404874 490102
rect 404930 490046 404998 490102
rect 405054 490046 405122 490102
rect 405178 490046 405246 490102
rect 405302 490046 435594 490102
rect 435650 490046 435718 490102
rect 435774 490046 435842 490102
rect 435898 490046 435966 490102
rect 436022 490046 466314 490102
rect 466370 490046 466438 490102
rect 466494 490046 466562 490102
rect 466618 490046 466686 490102
rect 466742 490046 497034 490102
rect 497090 490046 497158 490102
rect 497214 490046 497282 490102
rect 497338 490046 497406 490102
rect 497462 490046 527754 490102
rect 527810 490046 527878 490102
rect 527934 490046 528002 490102
rect 528058 490046 528126 490102
rect 528182 490046 558474 490102
rect 558530 490046 558598 490102
rect 558654 490046 558722 490102
rect 558778 490046 558846 490102
rect 558902 490046 589194 490102
rect 589250 490046 589318 490102
rect 589374 490046 589442 490102
rect 589498 490046 589566 490102
rect 589622 490046 596496 490102
rect 596552 490046 596620 490102
rect 596676 490046 596744 490102
rect 596800 490046 596868 490102
rect 596924 490046 597980 490102
rect -1916 489978 597980 490046
rect -1916 489922 -860 489978
rect -804 489922 -736 489978
rect -680 489922 -612 489978
rect -556 489922 -488 489978
rect -432 489922 5514 489978
rect 5570 489922 5638 489978
rect 5694 489922 5762 489978
rect 5818 489922 5886 489978
rect 5942 489922 36234 489978
rect 36290 489922 36358 489978
rect 36414 489922 36482 489978
rect 36538 489922 36606 489978
rect 36662 489922 66954 489978
rect 67010 489922 67078 489978
rect 67134 489922 67202 489978
rect 67258 489922 67326 489978
rect 67382 489922 97674 489978
rect 97730 489922 97798 489978
rect 97854 489922 97922 489978
rect 97978 489922 98046 489978
rect 98102 489922 128394 489978
rect 128450 489922 128518 489978
rect 128574 489922 128642 489978
rect 128698 489922 128766 489978
rect 128822 489922 159114 489978
rect 159170 489922 159238 489978
rect 159294 489922 159362 489978
rect 159418 489922 159486 489978
rect 159542 489922 189834 489978
rect 189890 489922 189958 489978
rect 190014 489922 190082 489978
rect 190138 489922 190206 489978
rect 190262 489922 220554 489978
rect 220610 489922 220678 489978
rect 220734 489922 220802 489978
rect 220858 489922 220926 489978
rect 220982 489922 251274 489978
rect 251330 489922 251398 489978
rect 251454 489922 251522 489978
rect 251578 489922 251646 489978
rect 251702 489922 281994 489978
rect 282050 489922 282118 489978
rect 282174 489922 282242 489978
rect 282298 489922 282366 489978
rect 282422 489922 312714 489978
rect 312770 489922 312838 489978
rect 312894 489922 312962 489978
rect 313018 489922 313086 489978
rect 313142 489922 343434 489978
rect 343490 489922 343558 489978
rect 343614 489922 343682 489978
rect 343738 489922 343806 489978
rect 343862 489922 374154 489978
rect 374210 489922 374278 489978
rect 374334 489922 374402 489978
rect 374458 489922 374526 489978
rect 374582 489922 404874 489978
rect 404930 489922 404998 489978
rect 405054 489922 405122 489978
rect 405178 489922 405246 489978
rect 405302 489922 435594 489978
rect 435650 489922 435718 489978
rect 435774 489922 435842 489978
rect 435898 489922 435966 489978
rect 436022 489922 466314 489978
rect 466370 489922 466438 489978
rect 466494 489922 466562 489978
rect 466618 489922 466686 489978
rect 466742 489922 497034 489978
rect 497090 489922 497158 489978
rect 497214 489922 497282 489978
rect 497338 489922 497406 489978
rect 497462 489922 527754 489978
rect 527810 489922 527878 489978
rect 527934 489922 528002 489978
rect 528058 489922 528126 489978
rect 528182 489922 558474 489978
rect 558530 489922 558598 489978
rect 558654 489922 558722 489978
rect 558778 489922 558846 489978
rect 558902 489922 589194 489978
rect 589250 489922 589318 489978
rect 589374 489922 589442 489978
rect 589498 489922 589566 489978
rect 589622 489922 596496 489978
rect 596552 489922 596620 489978
rect 596676 489922 596744 489978
rect 596800 489922 596868 489978
rect 596924 489922 597980 489978
rect -1916 489826 597980 489922
rect -1916 478350 597980 478446
rect -1916 478294 -1820 478350
rect -1764 478294 -1696 478350
rect -1640 478294 -1572 478350
rect -1516 478294 -1448 478350
rect -1392 478294 9234 478350
rect 9290 478294 9358 478350
rect 9414 478294 9482 478350
rect 9538 478294 9606 478350
rect 9662 478294 39954 478350
rect 40010 478294 40078 478350
rect 40134 478294 40202 478350
rect 40258 478294 40326 478350
rect 40382 478294 70674 478350
rect 70730 478294 70798 478350
rect 70854 478294 70922 478350
rect 70978 478294 71046 478350
rect 71102 478294 101394 478350
rect 101450 478294 101518 478350
rect 101574 478294 101642 478350
rect 101698 478294 101766 478350
rect 101822 478294 132114 478350
rect 132170 478294 132238 478350
rect 132294 478294 132362 478350
rect 132418 478294 132486 478350
rect 132542 478294 162834 478350
rect 162890 478294 162958 478350
rect 163014 478294 163082 478350
rect 163138 478294 163206 478350
rect 163262 478294 193554 478350
rect 193610 478294 193678 478350
rect 193734 478294 193802 478350
rect 193858 478294 193926 478350
rect 193982 478294 224274 478350
rect 224330 478294 224398 478350
rect 224454 478294 224522 478350
rect 224578 478294 224646 478350
rect 224702 478294 254994 478350
rect 255050 478294 255118 478350
rect 255174 478294 255242 478350
rect 255298 478294 255366 478350
rect 255422 478294 285714 478350
rect 285770 478294 285838 478350
rect 285894 478294 285962 478350
rect 286018 478294 286086 478350
rect 286142 478294 316434 478350
rect 316490 478294 316558 478350
rect 316614 478294 316682 478350
rect 316738 478294 316806 478350
rect 316862 478294 347154 478350
rect 347210 478294 347278 478350
rect 347334 478294 347402 478350
rect 347458 478294 347526 478350
rect 347582 478294 377874 478350
rect 377930 478294 377998 478350
rect 378054 478294 378122 478350
rect 378178 478294 378246 478350
rect 378302 478294 408594 478350
rect 408650 478294 408718 478350
rect 408774 478294 408842 478350
rect 408898 478294 408966 478350
rect 409022 478294 439314 478350
rect 439370 478294 439438 478350
rect 439494 478294 439562 478350
rect 439618 478294 439686 478350
rect 439742 478294 470034 478350
rect 470090 478294 470158 478350
rect 470214 478294 470282 478350
rect 470338 478294 470406 478350
rect 470462 478294 500754 478350
rect 500810 478294 500878 478350
rect 500934 478294 501002 478350
rect 501058 478294 501126 478350
rect 501182 478294 531474 478350
rect 531530 478294 531598 478350
rect 531654 478294 531722 478350
rect 531778 478294 531846 478350
rect 531902 478294 562194 478350
rect 562250 478294 562318 478350
rect 562374 478294 562442 478350
rect 562498 478294 562566 478350
rect 562622 478294 592914 478350
rect 592970 478294 593038 478350
rect 593094 478294 593162 478350
rect 593218 478294 593286 478350
rect 593342 478294 597456 478350
rect 597512 478294 597580 478350
rect 597636 478294 597704 478350
rect 597760 478294 597828 478350
rect 597884 478294 597980 478350
rect -1916 478226 597980 478294
rect -1916 478170 -1820 478226
rect -1764 478170 -1696 478226
rect -1640 478170 -1572 478226
rect -1516 478170 -1448 478226
rect -1392 478170 9234 478226
rect 9290 478170 9358 478226
rect 9414 478170 9482 478226
rect 9538 478170 9606 478226
rect 9662 478170 39954 478226
rect 40010 478170 40078 478226
rect 40134 478170 40202 478226
rect 40258 478170 40326 478226
rect 40382 478170 70674 478226
rect 70730 478170 70798 478226
rect 70854 478170 70922 478226
rect 70978 478170 71046 478226
rect 71102 478170 101394 478226
rect 101450 478170 101518 478226
rect 101574 478170 101642 478226
rect 101698 478170 101766 478226
rect 101822 478170 132114 478226
rect 132170 478170 132238 478226
rect 132294 478170 132362 478226
rect 132418 478170 132486 478226
rect 132542 478170 162834 478226
rect 162890 478170 162958 478226
rect 163014 478170 163082 478226
rect 163138 478170 163206 478226
rect 163262 478170 193554 478226
rect 193610 478170 193678 478226
rect 193734 478170 193802 478226
rect 193858 478170 193926 478226
rect 193982 478170 224274 478226
rect 224330 478170 224398 478226
rect 224454 478170 224522 478226
rect 224578 478170 224646 478226
rect 224702 478170 254994 478226
rect 255050 478170 255118 478226
rect 255174 478170 255242 478226
rect 255298 478170 255366 478226
rect 255422 478170 285714 478226
rect 285770 478170 285838 478226
rect 285894 478170 285962 478226
rect 286018 478170 286086 478226
rect 286142 478170 316434 478226
rect 316490 478170 316558 478226
rect 316614 478170 316682 478226
rect 316738 478170 316806 478226
rect 316862 478170 347154 478226
rect 347210 478170 347278 478226
rect 347334 478170 347402 478226
rect 347458 478170 347526 478226
rect 347582 478170 377874 478226
rect 377930 478170 377998 478226
rect 378054 478170 378122 478226
rect 378178 478170 378246 478226
rect 378302 478170 408594 478226
rect 408650 478170 408718 478226
rect 408774 478170 408842 478226
rect 408898 478170 408966 478226
rect 409022 478170 439314 478226
rect 439370 478170 439438 478226
rect 439494 478170 439562 478226
rect 439618 478170 439686 478226
rect 439742 478170 470034 478226
rect 470090 478170 470158 478226
rect 470214 478170 470282 478226
rect 470338 478170 470406 478226
rect 470462 478170 500754 478226
rect 500810 478170 500878 478226
rect 500934 478170 501002 478226
rect 501058 478170 501126 478226
rect 501182 478170 531474 478226
rect 531530 478170 531598 478226
rect 531654 478170 531722 478226
rect 531778 478170 531846 478226
rect 531902 478170 562194 478226
rect 562250 478170 562318 478226
rect 562374 478170 562442 478226
rect 562498 478170 562566 478226
rect 562622 478170 592914 478226
rect 592970 478170 593038 478226
rect 593094 478170 593162 478226
rect 593218 478170 593286 478226
rect 593342 478170 597456 478226
rect 597512 478170 597580 478226
rect 597636 478170 597704 478226
rect 597760 478170 597828 478226
rect 597884 478170 597980 478226
rect -1916 478102 597980 478170
rect -1916 478046 -1820 478102
rect -1764 478046 -1696 478102
rect -1640 478046 -1572 478102
rect -1516 478046 -1448 478102
rect -1392 478046 9234 478102
rect 9290 478046 9358 478102
rect 9414 478046 9482 478102
rect 9538 478046 9606 478102
rect 9662 478046 39954 478102
rect 40010 478046 40078 478102
rect 40134 478046 40202 478102
rect 40258 478046 40326 478102
rect 40382 478046 70674 478102
rect 70730 478046 70798 478102
rect 70854 478046 70922 478102
rect 70978 478046 71046 478102
rect 71102 478046 101394 478102
rect 101450 478046 101518 478102
rect 101574 478046 101642 478102
rect 101698 478046 101766 478102
rect 101822 478046 132114 478102
rect 132170 478046 132238 478102
rect 132294 478046 132362 478102
rect 132418 478046 132486 478102
rect 132542 478046 162834 478102
rect 162890 478046 162958 478102
rect 163014 478046 163082 478102
rect 163138 478046 163206 478102
rect 163262 478046 193554 478102
rect 193610 478046 193678 478102
rect 193734 478046 193802 478102
rect 193858 478046 193926 478102
rect 193982 478046 224274 478102
rect 224330 478046 224398 478102
rect 224454 478046 224522 478102
rect 224578 478046 224646 478102
rect 224702 478046 254994 478102
rect 255050 478046 255118 478102
rect 255174 478046 255242 478102
rect 255298 478046 255366 478102
rect 255422 478046 285714 478102
rect 285770 478046 285838 478102
rect 285894 478046 285962 478102
rect 286018 478046 286086 478102
rect 286142 478046 316434 478102
rect 316490 478046 316558 478102
rect 316614 478046 316682 478102
rect 316738 478046 316806 478102
rect 316862 478046 347154 478102
rect 347210 478046 347278 478102
rect 347334 478046 347402 478102
rect 347458 478046 347526 478102
rect 347582 478046 377874 478102
rect 377930 478046 377998 478102
rect 378054 478046 378122 478102
rect 378178 478046 378246 478102
rect 378302 478046 408594 478102
rect 408650 478046 408718 478102
rect 408774 478046 408842 478102
rect 408898 478046 408966 478102
rect 409022 478046 439314 478102
rect 439370 478046 439438 478102
rect 439494 478046 439562 478102
rect 439618 478046 439686 478102
rect 439742 478046 470034 478102
rect 470090 478046 470158 478102
rect 470214 478046 470282 478102
rect 470338 478046 470406 478102
rect 470462 478046 500754 478102
rect 500810 478046 500878 478102
rect 500934 478046 501002 478102
rect 501058 478046 501126 478102
rect 501182 478046 531474 478102
rect 531530 478046 531598 478102
rect 531654 478046 531722 478102
rect 531778 478046 531846 478102
rect 531902 478046 562194 478102
rect 562250 478046 562318 478102
rect 562374 478046 562442 478102
rect 562498 478046 562566 478102
rect 562622 478046 592914 478102
rect 592970 478046 593038 478102
rect 593094 478046 593162 478102
rect 593218 478046 593286 478102
rect 593342 478046 597456 478102
rect 597512 478046 597580 478102
rect 597636 478046 597704 478102
rect 597760 478046 597828 478102
rect 597884 478046 597980 478102
rect -1916 477978 597980 478046
rect -1916 477922 -1820 477978
rect -1764 477922 -1696 477978
rect -1640 477922 -1572 477978
rect -1516 477922 -1448 477978
rect -1392 477922 9234 477978
rect 9290 477922 9358 477978
rect 9414 477922 9482 477978
rect 9538 477922 9606 477978
rect 9662 477922 39954 477978
rect 40010 477922 40078 477978
rect 40134 477922 40202 477978
rect 40258 477922 40326 477978
rect 40382 477922 70674 477978
rect 70730 477922 70798 477978
rect 70854 477922 70922 477978
rect 70978 477922 71046 477978
rect 71102 477922 101394 477978
rect 101450 477922 101518 477978
rect 101574 477922 101642 477978
rect 101698 477922 101766 477978
rect 101822 477922 132114 477978
rect 132170 477922 132238 477978
rect 132294 477922 132362 477978
rect 132418 477922 132486 477978
rect 132542 477922 162834 477978
rect 162890 477922 162958 477978
rect 163014 477922 163082 477978
rect 163138 477922 163206 477978
rect 163262 477922 193554 477978
rect 193610 477922 193678 477978
rect 193734 477922 193802 477978
rect 193858 477922 193926 477978
rect 193982 477922 224274 477978
rect 224330 477922 224398 477978
rect 224454 477922 224522 477978
rect 224578 477922 224646 477978
rect 224702 477922 254994 477978
rect 255050 477922 255118 477978
rect 255174 477922 255242 477978
rect 255298 477922 255366 477978
rect 255422 477922 285714 477978
rect 285770 477922 285838 477978
rect 285894 477922 285962 477978
rect 286018 477922 286086 477978
rect 286142 477922 316434 477978
rect 316490 477922 316558 477978
rect 316614 477922 316682 477978
rect 316738 477922 316806 477978
rect 316862 477922 347154 477978
rect 347210 477922 347278 477978
rect 347334 477922 347402 477978
rect 347458 477922 347526 477978
rect 347582 477922 377874 477978
rect 377930 477922 377998 477978
rect 378054 477922 378122 477978
rect 378178 477922 378246 477978
rect 378302 477922 408594 477978
rect 408650 477922 408718 477978
rect 408774 477922 408842 477978
rect 408898 477922 408966 477978
rect 409022 477922 439314 477978
rect 439370 477922 439438 477978
rect 439494 477922 439562 477978
rect 439618 477922 439686 477978
rect 439742 477922 470034 477978
rect 470090 477922 470158 477978
rect 470214 477922 470282 477978
rect 470338 477922 470406 477978
rect 470462 477922 500754 477978
rect 500810 477922 500878 477978
rect 500934 477922 501002 477978
rect 501058 477922 501126 477978
rect 501182 477922 531474 477978
rect 531530 477922 531598 477978
rect 531654 477922 531722 477978
rect 531778 477922 531846 477978
rect 531902 477922 562194 477978
rect 562250 477922 562318 477978
rect 562374 477922 562442 477978
rect 562498 477922 562566 477978
rect 562622 477922 592914 477978
rect 592970 477922 593038 477978
rect 593094 477922 593162 477978
rect 593218 477922 593286 477978
rect 593342 477922 597456 477978
rect 597512 477922 597580 477978
rect 597636 477922 597704 477978
rect 597760 477922 597828 477978
rect 597884 477922 597980 477978
rect -1916 477826 597980 477922
rect -1916 472350 597980 472446
rect -1916 472294 -860 472350
rect -804 472294 -736 472350
rect -680 472294 -612 472350
rect -556 472294 -488 472350
rect -432 472294 5514 472350
rect 5570 472294 5638 472350
rect 5694 472294 5762 472350
rect 5818 472294 5886 472350
rect 5942 472294 36234 472350
rect 36290 472294 36358 472350
rect 36414 472294 36482 472350
rect 36538 472294 36606 472350
rect 36662 472294 66954 472350
rect 67010 472294 67078 472350
rect 67134 472294 67202 472350
rect 67258 472294 67326 472350
rect 67382 472294 97674 472350
rect 97730 472294 97798 472350
rect 97854 472294 97922 472350
rect 97978 472294 98046 472350
rect 98102 472294 128394 472350
rect 128450 472294 128518 472350
rect 128574 472294 128642 472350
rect 128698 472294 128766 472350
rect 128822 472294 159114 472350
rect 159170 472294 159238 472350
rect 159294 472294 159362 472350
rect 159418 472294 159486 472350
rect 159542 472294 189834 472350
rect 189890 472294 189958 472350
rect 190014 472294 190082 472350
rect 190138 472294 190206 472350
rect 190262 472294 220554 472350
rect 220610 472294 220678 472350
rect 220734 472294 220802 472350
rect 220858 472294 220926 472350
rect 220982 472294 251274 472350
rect 251330 472294 251398 472350
rect 251454 472294 251522 472350
rect 251578 472294 251646 472350
rect 251702 472294 281994 472350
rect 282050 472294 282118 472350
rect 282174 472294 282242 472350
rect 282298 472294 282366 472350
rect 282422 472294 312714 472350
rect 312770 472294 312838 472350
rect 312894 472294 312962 472350
rect 313018 472294 313086 472350
rect 313142 472294 343434 472350
rect 343490 472294 343558 472350
rect 343614 472294 343682 472350
rect 343738 472294 343806 472350
rect 343862 472294 374154 472350
rect 374210 472294 374278 472350
rect 374334 472294 374402 472350
rect 374458 472294 374526 472350
rect 374582 472294 404874 472350
rect 404930 472294 404998 472350
rect 405054 472294 405122 472350
rect 405178 472294 405246 472350
rect 405302 472294 435594 472350
rect 435650 472294 435718 472350
rect 435774 472294 435842 472350
rect 435898 472294 435966 472350
rect 436022 472294 466314 472350
rect 466370 472294 466438 472350
rect 466494 472294 466562 472350
rect 466618 472294 466686 472350
rect 466742 472294 497034 472350
rect 497090 472294 497158 472350
rect 497214 472294 497282 472350
rect 497338 472294 497406 472350
rect 497462 472294 527754 472350
rect 527810 472294 527878 472350
rect 527934 472294 528002 472350
rect 528058 472294 528126 472350
rect 528182 472294 558474 472350
rect 558530 472294 558598 472350
rect 558654 472294 558722 472350
rect 558778 472294 558846 472350
rect 558902 472294 589194 472350
rect 589250 472294 589318 472350
rect 589374 472294 589442 472350
rect 589498 472294 589566 472350
rect 589622 472294 596496 472350
rect 596552 472294 596620 472350
rect 596676 472294 596744 472350
rect 596800 472294 596868 472350
rect 596924 472294 597980 472350
rect -1916 472226 597980 472294
rect -1916 472170 -860 472226
rect -804 472170 -736 472226
rect -680 472170 -612 472226
rect -556 472170 -488 472226
rect -432 472170 5514 472226
rect 5570 472170 5638 472226
rect 5694 472170 5762 472226
rect 5818 472170 5886 472226
rect 5942 472170 36234 472226
rect 36290 472170 36358 472226
rect 36414 472170 36482 472226
rect 36538 472170 36606 472226
rect 36662 472170 66954 472226
rect 67010 472170 67078 472226
rect 67134 472170 67202 472226
rect 67258 472170 67326 472226
rect 67382 472170 97674 472226
rect 97730 472170 97798 472226
rect 97854 472170 97922 472226
rect 97978 472170 98046 472226
rect 98102 472170 128394 472226
rect 128450 472170 128518 472226
rect 128574 472170 128642 472226
rect 128698 472170 128766 472226
rect 128822 472170 159114 472226
rect 159170 472170 159238 472226
rect 159294 472170 159362 472226
rect 159418 472170 159486 472226
rect 159542 472170 189834 472226
rect 189890 472170 189958 472226
rect 190014 472170 190082 472226
rect 190138 472170 190206 472226
rect 190262 472170 220554 472226
rect 220610 472170 220678 472226
rect 220734 472170 220802 472226
rect 220858 472170 220926 472226
rect 220982 472170 251274 472226
rect 251330 472170 251398 472226
rect 251454 472170 251522 472226
rect 251578 472170 251646 472226
rect 251702 472170 281994 472226
rect 282050 472170 282118 472226
rect 282174 472170 282242 472226
rect 282298 472170 282366 472226
rect 282422 472170 312714 472226
rect 312770 472170 312838 472226
rect 312894 472170 312962 472226
rect 313018 472170 313086 472226
rect 313142 472170 343434 472226
rect 343490 472170 343558 472226
rect 343614 472170 343682 472226
rect 343738 472170 343806 472226
rect 343862 472170 374154 472226
rect 374210 472170 374278 472226
rect 374334 472170 374402 472226
rect 374458 472170 374526 472226
rect 374582 472170 404874 472226
rect 404930 472170 404998 472226
rect 405054 472170 405122 472226
rect 405178 472170 405246 472226
rect 405302 472170 435594 472226
rect 435650 472170 435718 472226
rect 435774 472170 435842 472226
rect 435898 472170 435966 472226
rect 436022 472170 466314 472226
rect 466370 472170 466438 472226
rect 466494 472170 466562 472226
rect 466618 472170 466686 472226
rect 466742 472170 497034 472226
rect 497090 472170 497158 472226
rect 497214 472170 497282 472226
rect 497338 472170 497406 472226
rect 497462 472170 527754 472226
rect 527810 472170 527878 472226
rect 527934 472170 528002 472226
rect 528058 472170 528126 472226
rect 528182 472170 558474 472226
rect 558530 472170 558598 472226
rect 558654 472170 558722 472226
rect 558778 472170 558846 472226
rect 558902 472170 589194 472226
rect 589250 472170 589318 472226
rect 589374 472170 589442 472226
rect 589498 472170 589566 472226
rect 589622 472170 596496 472226
rect 596552 472170 596620 472226
rect 596676 472170 596744 472226
rect 596800 472170 596868 472226
rect 596924 472170 597980 472226
rect -1916 472102 597980 472170
rect -1916 472046 -860 472102
rect -804 472046 -736 472102
rect -680 472046 -612 472102
rect -556 472046 -488 472102
rect -432 472046 5514 472102
rect 5570 472046 5638 472102
rect 5694 472046 5762 472102
rect 5818 472046 5886 472102
rect 5942 472046 36234 472102
rect 36290 472046 36358 472102
rect 36414 472046 36482 472102
rect 36538 472046 36606 472102
rect 36662 472046 66954 472102
rect 67010 472046 67078 472102
rect 67134 472046 67202 472102
rect 67258 472046 67326 472102
rect 67382 472046 97674 472102
rect 97730 472046 97798 472102
rect 97854 472046 97922 472102
rect 97978 472046 98046 472102
rect 98102 472046 128394 472102
rect 128450 472046 128518 472102
rect 128574 472046 128642 472102
rect 128698 472046 128766 472102
rect 128822 472046 159114 472102
rect 159170 472046 159238 472102
rect 159294 472046 159362 472102
rect 159418 472046 159486 472102
rect 159542 472046 189834 472102
rect 189890 472046 189958 472102
rect 190014 472046 190082 472102
rect 190138 472046 190206 472102
rect 190262 472046 220554 472102
rect 220610 472046 220678 472102
rect 220734 472046 220802 472102
rect 220858 472046 220926 472102
rect 220982 472046 251274 472102
rect 251330 472046 251398 472102
rect 251454 472046 251522 472102
rect 251578 472046 251646 472102
rect 251702 472046 281994 472102
rect 282050 472046 282118 472102
rect 282174 472046 282242 472102
rect 282298 472046 282366 472102
rect 282422 472046 312714 472102
rect 312770 472046 312838 472102
rect 312894 472046 312962 472102
rect 313018 472046 313086 472102
rect 313142 472046 343434 472102
rect 343490 472046 343558 472102
rect 343614 472046 343682 472102
rect 343738 472046 343806 472102
rect 343862 472046 374154 472102
rect 374210 472046 374278 472102
rect 374334 472046 374402 472102
rect 374458 472046 374526 472102
rect 374582 472046 404874 472102
rect 404930 472046 404998 472102
rect 405054 472046 405122 472102
rect 405178 472046 405246 472102
rect 405302 472046 435594 472102
rect 435650 472046 435718 472102
rect 435774 472046 435842 472102
rect 435898 472046 435966 472102
rect 436022 472046 466314 472102
rect 466370 472046 466438 472102
rect 466494 472046 466562 472102
rect 466618 472046 466686 472102
rect 466742 472046 497034 472102
rect 497090 472046 497158 472102
rect 497214 472046 497282 472102
rect 497338 472046 497406 472102
rect 497462 472046 527754 472102
rect 527810 472046 527878 472102
rect 527934 472046 528002 472102
rect 528058 472046 528126 472102
rect 528182 472046 558474 472102
rect 558530 472046 558598 472102
rect 558654 472046 558722 472102
rect 558778 472046 558846 472102
rect 558902 472046 589194 472102
rect 589250 472046 589318 472102
rect 589374 472046 589442 472102
rect 589498 472046 589566 472102
rect 589622 472046 596496 472102
rect 596552 472046 596620 472102
rect 596676 472046 596744 472102
rect 596800 472046 596868 472102
rect 596924 472046 597980 472102
rect -1916 471978 597980 472046
rect -1916 471922 -860 471978
rect -804 471922 -736 471978
rect -680 471922 -612 471978
rect -556 471922 -488 471978
rect -432 471922 5514 471978
rect 5570 471922 5638 471978
rect 5694 471922 5762 471978
rect 5818 471922 5886 471978
rect 5942 471922 36234 471978
rect 36290 471922 36358 471978
rect 36414 471922 36482 471978
rect 36538 471922 36606 471978
rect 36662 471922 66954 471978
rect 67010 471922 67078 471978
rect 67134 471922 67202 471978
rect 67258 471922 67326 471978
rect 67382 471922 97674 471978
rect 97730 471922 97798 471978
rect 97854 471922 97922 471978
rect 97978 471922 98046 471978
rect 98102 471922 128394 471978
rect 128450 471922 128518 471978
rect 128574 471922 128642 471978
rect 128698 471922 128766 471978
rect 128822 471922 159114 471978
rect 159170 471922 159238 471978
rect 159294 471922 159362 471978
rect 159418 471922 159486 471978
rect 159542 471922 189834 471978
rect 189890 471922 189958 471978
rect 190014 471922 190082 471978
rect 190138 471922 190206 471978
rect 190262 471922 220554 471978
rect 220610 471922 220678 471978
rect 220734 471922 220802 471978
rect 220858 471922 220926 471978
rect 220982 471922 251274 471978
rect 251330 471922 251398 471978
rect 251454 471922 251522 471978
rect 251578 471922 251646 471978
rect 251702 471922 281994 471978
rect 282050 471922 282118 471978
rect 282174 471922 282242 471978
rect 282298 471922 282366 471978
rect 282422 471922 312714 471978
rect 312770 471922 312838 471978
rect 312894 471922 312962 471978
rect 313018 471922 313086 471978
rect 313142 471922 343434 471978
rect 343490 471922 343558 471978
rect 343614 471922 343682 471978
rect 343738 471922 343806 471978
rect 343862 471922 374154 471978
rect 374210 471922 374278 471978
rect 374334 471922 374402 471978
rect 374458 471922 374526 471978
rect 374582 471922 404874 471978
rect 404930 471922 404998 471978
rect 405054 471922 405122 471978
rect 405178 471922 405246 471978
rect 405302 471922 435594 471978
rect 435650 471922 435718 471978
rect 435774 471922 435842 471978
rect 435898 471922 435966 471978
rect 436022 471922 466314 471978
rect 466370 471922 466438 471978
rect 466494 471922 466562 471978
rect 466618 471922 466686 471978
rect 466742 471922 497034 471978
rect 497090 471922 497158 471978
rect 497214 471922 497282 471978
rect 497338 471922 497406 471978
rect 497462 471922 527754 471978
rect 527810 471922 527878 471978
rect 527934 471922 528002 471978
rect 528058 471922 528126 471978
rect 528182 471922 558474 471978
rect 558530 471922 558598 471978
rect 558654 471922 558722 471978
rect 558778 471922 558846 471978
rect 558902 471922 589194 471978
rect 589250 471922 589318 471978
rect 589374 471922 589442 471978
rect 589498 471922 589566 471978
rect 589622 471922 596496 471978
rect 596552 471922 596620 471978
rect 596676 471922 596744 471978
rect 596800 471922 596868 471978
rect 596924 471922 597980 471978
rect -1916 471826 597980 471922
rect -1916 460350 597980 460446
rect -1916 460294 -1820 460350
rect -1764 460294 -1696 460350
rect -1640 460294 -1572 460350
rect -1516 460294 -1448 460350
rect -1392 460294 9234 460350
rect 9290 460294 9358 460350
rect 9414 460294 9482 460350
rect 9538 460294 9606 460350
rect 9662 460294 39954 460350
rect 40010 460294 40078 460350
rect 40134 460294 40202 460350
rect 40258 460294 40326 460350
rect 40382 460294 70674 460350
rect 70730 460294 70798 460350
rect 70854 460294 70922 460350
rect 70978 460294 71046 460350
rect 71102 460294 101394 460350
rect 101450 460294 101518 460350
rect 101574 460294 101642 460350
rect 101698 460294 101766 460350
rect 101822 460294 132114 460350
rect 132170 460294 132238 460350
rect 132294 460294 132362 460350
rect 132418 460294 132486 460350
rect 132542 460294 162834 460350
rect 162890 460294 162958 460350
rect 163014 460294 163082 460350
rect 163138 460294 163206 460350
rect 163262 460294 193554 460350
rect 193610 460294 193678 460350
rect 193734 460294 193802 460350
rect 193858 460294 193926 460350
rect 193982 460294 224274 460350
rect 224330 460294 224398 460350
rect 224454 460294 224522 460350
rect 224578 460294 224646 460350
rect 224702 460294 254994 460350
rect 255050 460294 255118 460350
rect 255174 460294 255242 460350
rect 255298 460294 255366 460350
rect 255422 460294 285714 460350
rect 285770 460294 285838 460350
rect 285894 460294 285962 460350
rect 286018 460294 286086 460350
rect 286142 460294 316434 460350
rect 316490 460294 316558 460350
rect 316614 460294 316682 460350
rect 316738 460294 316806 460350
rect 316862 460294 347154 460350
rect 347210 460294 347278 460350
rect 347334 460294 347402 460350
rect 347458 460294 347526 460350
rect 347582 460294 377874 460350
rect 377930 460294 377998 460350
rect 378054 460294 378122 460350
rect 378178 460294 378246 460350
rect 378302 460294 408594 460350
rect 408650 460294 408718 460350
rect 408774 460294 408842 460350
rect 408898 460294 408966 460350
rect 409022 460294 439314 460350
rect 439370 460294 439438 460350
rect 439494 460294 439562 460350
rect 439618 460294 439686 460350
rect 439742 460294 470034 460350
rect 470090 460294 470158 460350
rect 470214 460294 470282 460350
rect 470338 460294 470406 460350
rect 470462 460294 500754 460350
rect 500810 460294 500878 460350
rect 500934 460294 501002 460350
rect 501058 460294 501126 460350
rect 501182 460294 531474 460350
rect 531530 460294 531598 460350
rect 531654 460294 531722 460350
rect 531778 460294 531846 460350
rect 531902 460294 562194 460350
rect 562250 460294 562318 460350
rect 562374 460294 562442 460350
rect 562498 460294 562566 460350
rect 562622 460294 592914 460350
rect 592970 460294 593038 460350
rect 593094 460294 593162 460350
rect 593218 460294 593286 460350
rect 593342 460294 597456 460350
rect 597512 460294 597580 460350
rect 597636 460294 597704 460350
rect 597760 460294 597828 460350
rect 597884 460294 597980 460350
rect -1916 460226 597980 460294
rect -1916 460170 -1820 460226
rect -1764 460170 -1696 460226
rect -1640 460170 -1572 460226
rect -1516 460170 -1448 460226
rect -1392 460170 9234 460226
rect 9290 460170 9358 460226
rect 9414 460170 9482 460226
rect 9538 460170 9606 460226
rect 9662 460170 39954 460226
rect 40010 460170 40078 460226
rect 40134 460170 40202 460226
rect 40258 460170 40326 460226
rect 40382 460170 70674 460226
rect 70730 460170 70798 460226
rect 70854 460170 70922 460226
rect 70978 460170 71046 460226
rect 71102 460170 101394 460226
rect 101450 460170 101518 460226
rect 101574 460170 101642 460226
rect 101698 460170 101766 460226
rect 101822 460170 132114 460226
rect 132170 460170 132238 460226
rect 132294 460170 132362 460226
rect 132418 460170 132486 460226
rect 132542 460170 162834 460226
rect 162890 460170 162958 460226
rect 163014 460170 163082 460226
rect 163138 460170 163206 460226
rect 163262 460170 193554 460226
rect 193610 460170 193678 460226
rect 193734 460170 193802 460226
rect 193858 460170 193926 460226
rect 193982 460170 224274 460226
rect 224330 460170 224398 460226
rect 224454 460170 224522 460226
rect 224578 460170 224646 460226
rect 224702 460170 254994 460226
rect 255050 460170 255118 460226
rect 255174 460170 255242 460226
rect 255298 460170 255366 460226
rect 255422 460170 285714 460226
rect 285770 460170 285838 460226
rect 285894 460170 285962 460226
rect 286018 460170 286086 460226
rect 286142 460170 316434 460226
rect 316490 460170 316558 460226
rect 316614 460170 316682 460226
rect 316738 460170 316806 460226
rect 316862 460170 347154 460226
rect 347210 460170 347278 460226
rect 347334 460170 347402 460226
rect 347458 460170 347526 460226
rect 347582 460170 377874 460226
rect 377930 460170 377998 460226
rect 378054 460170 378122 460226
rect 378178 460170 378246 460226
rect 378302 460170 408594 460226
rect 408650 460170 408718 460226
rect 408774 460170 408842 460226
rect 408898 460170 408966 460226
rect 409022 460170 439314 460226
rect 439370 460170 439438 460226
rect 439494 460170 439562 460226
rect 439618 460170 439686 460226
rect 439742 460170 470034 460226
rect 470090 460170 470158 460226
rect 470214 460170 470282 460226
rect 470338 460170 470406 460226
rect 470462 460170 500754 460226
rect 500810 460170 500878 460226
rect 500934 460170 501002 460226
rect 501058 460170 501126 460226
rect 501182 460170 531474 460226
rect 531530 460170 531598 460226
rect 531654 460170 531722 460226
rect 531778 460170 531846 460226
rect 531902 460170 562194 460226
rect 562250 460170 562318 460226
rect 562374 460170 562442 460226
rect 562498 460170 562566 460226
rect 562622 460170 592914 460226
rect 592970 460170 593038 460226
rect 593094 460170 593162 460226
rect 593218 460170 593286 460226
rect 593342 460170 597456 460226
rect 597512 460170 597580 460226
rect 597636 460170 597704 460226
rect 597760 460170 597828 460226
rect 597884 460170 597980 460226
rect -1916 460102 597980 460170
rect -1916 460046 -1820 460102
rect -1764 460046 -1696 460102
rect -1640 460046 -1572 460102
rect -1516 460046 -1448 460102
rect -1392 460046 9234 460102
rect 9290 460046 9358 460102
rect 9414 460046 9482 460102
rect 9538 460046 9606 460102
rect 9662 460046 39954 460102
rect 40010 460046 40078 460102
rect 40134 460046 40202 460102
rect 40258 460046 40326 460102
rect 40382 460046 70674 460102
rect 70730 460046 70798 460102
rect 70854 460046 70922 460102
rect 70978 460046 71046 460102
rect 71102 460046 101394 460102
rect 101450 460046 101518 460102
rect 101574 460046 101642 460102
rect 101698 460046 101766 460102
rect 101822 460046 132114 460102
rect 132170 460046 132238 460102
rect 132294 460046 132362 460102
rect 132418 460046 132486 460102
rect 132542 460046 162834 460102
rect 162890 460046 162958 460102
rect 163014 460046 163082 460102
rect 163138 460046 163206 460102
rect 163262 460046 193554 460102
rect 193610 460046 193678 460102
rect 193734 460046 193802 460102
rect 193858 460046 193926 460102
rect 193982 460046 224274 460102
rect 224330 460046 224398 460102
rect 224454 460046 224522 460102
rect 224578 460046 224646 460102
rect 224702 460046 254994 460102
rect 255050 460046 255118 460102
rect 255174 460046 255242 460102
rect 255298 460046 255366 460102
rect 255422 460046 285714 460102
rect 285770 460046 285838 460102
rect 285894 460046 285962 460102
rect 286018 460046 286086 460102
rect 286142 460046 316434 460102
rect 316490 460046 316558 460102
rect 316614 460046 316682 460102
rect 316738 460046 316806 460102
rect 316862 460046 347154 460102
rect 347210 460046 347278 460102
rect 347334 460046 347402 460102
rect 347458 460046 347526 460102
rect 347582 460046 377874 460102
rect 377930 460046 377998 460102
rect 378054 460046 378122 460102
rect 378178 460046 378246 460102
rect 378302 460046 408594 460102
rect 408650 460046 408718 460102
rect 408774 460046 408842 460102
rect 408898 460046 408966 460102
rect 409022 460046 439314 460102
rect 439370 460046 439438 460102
rect 439494 460046 439562 460102
rect 439618 460046 439686 460102
rect 439742 460046 470034 460102
rect 470090 460046 470158 460102
rect 470214 460046 470282 460102
rect 470338 460046 470406 460102
rect 470462 460046 500754 460102
rect 500810 460046 500878 460102
rect 500934 460046 501002 460102
rect 501058 460046 501126 460102
rect 501182 460046 531474 460102
rect 531530 460046 531598 460102
rect 531654 460046 531722 460102
rect 531778 460046 531846 460102
rect 531902 460046 562194 460102
rect 562250 460046 562318 460102
rect 562374 460046 562442 460102
rect 562498 460046 562566 460102
rect 562622 460046 592914 460102
rect 592970 460046 593038 460102
rect 593094 460046 593162 460102
rect 593218 460046 593286 460102
rect 593342 460046 597456 460102
rect 597512 460046 597580 460102
rect 597636 460046 597704 460102
rect 597760 460046 597828 460102
rect 597884 460046 597980 460102
rect -1916 459978 597980 460046
rect -1916 459922 -1820 459978
rect -1764 459922 -1696 459978
rect -1640 459922 -1572 459978
rect -1516 459922 -1448 459978
rect -1392 459922 9234 459978
rect 9290 459922 9358 459978
rect 9414 459922 9482 459978
rect 9538 459922 9606 459978
rect 9662 459922 39954 459978
rect 40010 459922 40078 459978
rect 40134 459922 40202 459978
rect 40258 459922 40326 459978
rect 40382 459922 70674 459978
rect 70730 459922 70798 459978
rect 70854 459922 70922 459978
rect 70978 459922 71046 459978
rect 71102 459922 101394 459978
rect 101450 459922 101518 459978
rect 101574 459922 101642 459978
rect 101698 459922 101766 459978
rect 101822 459922 132114 459978
rect 132170 459922 132238 459978
rect 132294 459922 132362 459978
rect 132418 459922 132486 459978
rect 132542 459922 162834 459978
rect 162890 459922 162958 459978
rect 163014 459922 163082 459978
rect 163138 459922 163206 459978
rect 163262 459922 193554 459978
rect 193610 459922 193678 459978
rect 193734 459922 193802 459978
rect 193858 459922 193926 459978
rect 193982 459922 224274 459978
rect 224330 459922 224398 459978
rect 224454 459922 224522 459978
rect 224578 459922 224646 459978
rect 224702 459922 254994 459978
rect 255050 459922 255118 459978
rect 255174 459922 255242 459978
rect 255298 459922 255366 459978
rect 255422 459922 285714 459978
rect 285770 459922 285838 459978
rect 285894 459922 285962 459978
rect 286018 459922 286086 459978
rect 286142 459922 316434 459978
rect 316490 459922 316558 459978
rect 316614 459922 316682 459978
rect 316738 459922 316806 459978
rect 316862 459922 347154 459978
rect 347210 459922 347278 459978
rect 347334 459922 347402 459978
rect 347458 459922 347526 459978
rect 347582 459922 377874 459978
rect 377930 459922 377998 459978
rect 378054 459922 378122 459978
rect 378178 459922 378246 459978
rect 378302 459922 408594 459978
rect 408650 459922 408718 459978
rect 408774 459922 408842 459978
rect 408898 459922 408966 459978
rect 409022 459922 439314 459978
rect 439370 459922 439438 459978
rect 439494 459922 439562 459978
rect 439618 459922 439686 459978
rect 439742 459922 470034 459978
rect 470090 459922 470158 459978
rect 470214 459922 470282 459978
rect 470338 459922 470406 459978
rect 470462 459922 500754 459978
rect 500810 459922 500878 459978
rect 500934 459922 501002 459978
rect 501058 459922 501126 459978
rect 501182 459922 531474 459978
rect 531530 459922 531598 459978
rect 531654 459922 531722 459978
rect 531778 459922 531846 459978
rect 531902 459922 562194 459978
rect 562250 459922 562318 459978
rect 562374 459922 562442 459978
rect 562498 459922 562566 459978
rect 562622 459922 592914 459978
rect 592970 459922 593038 459978
rect 593094 459922 593162 459978
rect 593218 459922 593286 459978
rect 593342 459922 597456 459978
rect 597512 459922 597580 459978
rect 597636 459922 597704 459978
rect 597760 459922 597828 459978
rect 597884 459922 597980 459978
rect -1916 459826 597980 459922
rect -1916 454350 597980 454446
rect -1916 454294 -860 454350
rect -804 454294 -736 454350
rect -680 454294 -612 454350
rect -556 454294 -488 454350
rect -432 454294 5514 454350
rect 5570 454294 5638 454350
rect 5694 454294 5762 454350
rect 5818 454294 5886 454350
rect 5942 454294 36234 454350
rect 36290 454294 36358 454350
rect 36414 454294 36482 454350
rect 36538 454294 36606 454350
rect 36662 454294 66954 454350
rect 67010 454294 67078 454350
rect 67134 454294 67202 454350
rect 67258 454294 67326 454350
rect 67382 454294 97674 454350
rect 97730 454294 97798 454350
rect 97854 454294 97922 454350
rect 97978 454294 98046 454350
rect 98102 454294 128394 454350
rect 128450 454294 128518 454350
rect 128574 454294 128642 454350
rect 128698 454294 128766 454350
rect 128822 454294 159114 454350
rect 159170 454294 159238 454350
rect 159294 454294 159362 454350
rect 159418 454294 159486 454350
rect 159542 454294 189834 454350
rect 189890 454294 189958 454350
rect 190014 454294 190082 454350
rect 190138 454294 190206 454350
rect 190262 454294 220554 454350
rect 220610 454294 220678 454350
rect 220734 454294 220802 454350
rect 220858 454294 220926 454350
rect 220982 454294 251274 454350
rect 251330 454294 251398 454350
rect 251454 454294 251522 454350
rect 251578 454294 251646 454350
rect 251702 454294 281994 454350
rect 282050 454294 282118 454350
rect 282174 454294 282242 454350
rect 282298 454294 282366 454350
rect 282422 454294 312714 454350
rect 312770 454294 312838 454350
rect 312894 454294 312962 454350
rect 313018 454294 313086 454350
rect 313142 454294 343434 454350
rect 343490 454294 343558 454350
rect 343614 454294 343682 454350
rect 343738 454294 343806 454350
rect 343862 454294 374154 454350
rect 374210 454294 374278 454350
rect 374334 454294 374402 454350
rect 374458 454294 374526 454350
rect 374582 454294 404874 454350
rect 404930 454294 404998 454350
rect 405054 454294 405122 454350
rect 405178 454294 405246 454350
rect 405302 454294 435594 454350
rect 435650 454294 435718 454350
rect 435774 454294 435842 454350
rect 435898 454294 435966 454350
rect 436022 454294 466314 454350
rect 466370 454294 466438 454350
rect 466494 454294 466562 454350
rect 466618 454294 466686 454350
rect 466742 454294 497034 454350
rect 497090 454294 497158 454350
rect 497214 454294 497282 454350
rect 497338 454294 497406 454350
rect 497462 454294 527754 454350
rect 527810 454294 527878 454350
rect 527934 454294 528002 454350
rect 528058 454294 528126 454350
rect 528182 454294 558474 454350
rect 558530 454294 558598 454350
rect 558654 454294 558722 454350
rect 558778 454294 558846 454350
rect 558902 454294 589194 454350
rect 589250 454294 589318 454350
rect 589374 454294 589442 454350
rect 589498 454294 589566 454350
rect 589622 454294 596496 454350
rect 596552 454294 596620 454350
rect 596676 454294 596744 454350
rect 596800 454294 596868 454350
rect 596924 454294 597980 454350
rect -1916 454226 597980 454294
rect -1916 454170 -860 454226
rect -804 454170 -736 454226
rect -680 454170 -612 454226
rect -556 454170 -488 454226
rect -432 454170 5514 454226
rect 5570 454170 5638 454226
rect 5694 454170 5762 454226
rect 5818 454170 5886 454226
rect 5942 454170 36234 454226
rect 36290 454170 36358 454226
rect 36414 454170 36482 454226
rect 36538 454170 36606 454226
rect 36662 454170 66954 454226
rect 67010 454170 67078 454226
rect 67134 454170 67202 454226
rect 67258 454170 67326 454226
rect 67382 454170 97674 454226
rect 97730 454170 97798 454226
rect 97854 454170 97922 454226
rect 97978 454170 98046 454226
rect 98102 454170 128394 454226
rect 128450 454170 128518 454226
rect 128574 454170 128642 454226
rect 128698 454170 128766 454226
rect 128822 454170 159114 454226
rect 159170 454170 159238 454226
rect 159294 454170 159362 454226
rect 159418 454170 159486 454226
rect 159542 454170 189834 454226
rect 189890 454170 189958 454226
rect 190014 454170 190082 454226
rect 190138 454170 190206 454226
rect 190262 454170 220554 454226
rect 220610 454170 220678 454226
rect 220734 454170 220802 454226
rect 220858 454170 220926 454226
rect 220982 454170 251274 454226
rect 251330 454170 251398 454226
rect 251454 454170 251522 454226
rect 251578 454170 251646 454226
rect 251702 454170 281994 454226
rect 282050 454170 282118 454226
rect 282174 454170 282242 454226
rect 282298 454170 282366 454226
rect 282422 454170 312714 454226
rect 312770 454170 312838 454226
rect 312894 454170 312962 454226
rect 313018 454170 313086 454226
rect 313142 454170 343434 454226
rect 343490 454170 343558 454226
rect 343614 454170 343682 454226
rect 343738 454170 343806 454226
rect 343862 454170 374154 454226
rect 374210 454170 374278 454226
rect 374334 454170 374402 454226
rect 374458 454170 374526 454226
rect 374582 454170 404874 454226
rect 404930 454170 404998 454226
rect 405054 454170 405122 454226
rect 405178 454170 405246 454226
rect 405302 454170 435594 454226
rect 435650 454170 435718 454226
rect 435774 454170 435842 454226
rect 435898 454170 435966 454226
rect 436022 454170 466314 454226
rect 466370 454170 466438 454226
rect 466494 454170 466562 454226
rect 466618 454170 466686 454226
rect 466742 454170 497034 454226
rect 497090 454170 497158 454226
rect 497214 454170 497282 454226
rect 497338 454170 497406 454226
rect 497462 454170 527754 454226
rect 527810 454170 527878 454226
rect 527934 454170 528002 454226
rect 528058 454170 528126 454226
rect 528182 454170 558474 454226
rect 558530 454170 558598 454226
rect 558654 454170 558722 454226
rect 558778 454170 558846 454226
rect 558902 454170 589194 454226
rect 589250 454170 589318 454226
rect 589374 454170 589442 454226
rect 589498 454170 589566 454226
rect 589622 454170 596496 454226
rect 596552 454170 596620 454226
rect 596676 454170 596744 454226
rect 596800 454170 596868 454226
rect 596924 454170 597980 454226
rect -1916 454102 597980 454170
rect -1916 454046 -860 454102
rect -804 454046 -736 454102
rect -680 454046 -612 454102
rect -556 454046 -488 454102
rect -432 454046 5514 454102
rect 5570 454046 5638 454102
rect 5694 454046 5762 454102
rect 5818 454046 5886 454102
rect 5942 454046 36234 454102
rect 36290 454046 36358 454102
rect 36414 454046 36482 454102
rect 36538 454046 36606 454102
rect 36662 454046 66954 454102
rect 67010 454046 67078 454102
rect 67134 454046 67202 454102
rect 67258 454046 67326 454102
rect 67382 454046 97674 454102
rect 97730 454046 97798 454102
rect 97854 454046 97922 454102
rect 97978 454046 98046 454102
rect 98102 454046 128394 454102
rect 128450 454046 128518 454102
rect 128574 454046 128642 454102
rect 128698 454046 128766 454102
rect 128822 454046 159114 454102
rect 159170 454046 159238 454102
rect 159294 454046 159362 454102
rect 159418 454046 159486 454102
rect 159542 454046 189834 454102
rect 189890 454046 189958 454102
rect 190014 454046 190082 454102
rect 190138 454046 190206 454102
rect 190262 454046 220554 454102
rect 220610 454046 220678 454102
rect 220734 454046 220802 454102
rect 220858 454046 220926 454102
rect 220982 454046 251274 454102
rect 251330 454046 251398 454102
rect 251454 454046 251522 454102
rect 251578 454046 251646 454102
rect 251702 454046 281994 454102
rect 282050 454046 282118 454102
rect 282174 454046 282242 454102
rect 282298 454046 282366 454102
rect 282422 454046 312714 454102
rect 312770 454046 312838 454102
rect 312894 454046 312962 454102
rect 313018 454046 313086 454102
rect 313142 454046 343434 454102
rect 343490 454046 343558 454102
rect 343614 454046 343682 454102
rect 343738 454046 343806 454102
rect 343862 454046 374154 454102
rect 374210 454046 374278 454102
rect 374334 454046 374402 454102
rect 374458 454046 374526 454102
rect 374582 454046 404874 454102
rect 404930 454046 404998 454102
rect 405054 454046 405122 454102
rect 405178 454046 405246 454102
rect 405302 454046 435594 454102
rect 435650 454046 435718 454102
rect 435774 454046 435842 454102
rect 435898 454046 435966 454102
rect 436022 454046 466314 454102
rect 466370 454046 466438 454102
rect 466494 454046 466562 454102
rect 466618 454046 466686 454102
rect 466742 454046 497034 454102
rect 497090 454046 497158 454102
rect 497214 454046 497282 454102
rect 497338 454046 497406 454102
rect 497462 454046 527754 454102
rect 527810 454046 527878 454102
rect 527934 454046 528002 454102
rect 528058 454046 528126 454102
rect 528182 454046 558474 454102
rect 558530 454046 558598 454102
rect 558654 454046 558722 454102
rect 558778 454046 558846 454102
rect 558902 454046 589194 454102
rect 589250 454046 589318 454102
rect 589374 454046 589442 454102
rect 589498 454046 589566 454102
rect 589622 454046 596496 454102
rect 596552 454046 596620 454102
rect 596676 454046 596744 454102
rect 596800 454046 596868 454102
rect 596924 454046 597980 454102
rect -1916 453978 597980 454046
rect -1916 453922 -860 453978
rect -804 453922 -736 453978
rect -680 453922 -612 453978
rect -556 453922 -488 453978
rect -432 453922 5514 453978
rect 5570 453922 5638 453978
rect 5694 453922 5762 453978
rect 5818 453922 5886 453978
rect 5942 453922 36234 453978
rect 36290 453922 36358 453978
rect 36414 453922 36482 453978
rect 36538 453922 36606 453978
rect 36662 453922 66954 453978
rect 67010 453922 67078 453978
rect 67134 453922 67202 453978
rect 67258 453922 67326 453978
rect 67382 453922 97674 453978
rect 97730 453922 97798 453978
rect 97854 453922 97922 453978
rect 97978 453922 98046 453978
rect 98102 453922 128394 453978
rect 128450 453922 128518 453978
rect 128574 453922 128642 453978
rect 128698 453922 128766 453978
rect 128822 453922 159114 453978
rect 159170 453922 159238 453978
rect 159294 453922 159362 453978
rect 159418 453922 159486 453978
rect 159542 453922 189834 453978
rect 189890 453922 189958 453978
rect 190014 453922 190082 453978
rect 190138 453922 190206 453978
rect 190262 453922 220554 453978
rect 220610 453922 220678 453978
rect 220734 453922 220802 453978
rect 220858 453922 220926 453978
rect 220982 453922 251274 453978
rect 251330 453922 251398 453978
rect 251454 453922 251522 453978
rect 251578 453922 251646 453978
rect 251702 453922 281994 453978
rect 282050 453922 282118 453978
rect 282174 453922 282242 453978
rect 282298 453922 282366 453978
rect 282422 453922 312714 453978
rect 312770 453922 312838 453978
rect 312894 453922 312962 453978
rect 313018 453922 313086 453978
rect 313142 453922 343434 453978
rect 343490 453922 343558 453978
rect 343614 453922 343682 453978
rect 343738 453922 343806 453978
rect 343862 453922 374154 453978
rect 374210 453922 374278 453978
rect 374334 453922 374402 453978
rect 374458 453922 374526 453978
rect 374582 453922 404874 453978
rect 404930 453922 404998 453978
rect 405054 453922 405122 453978
rect 405178 453922 405246 453978
rect 405302 453922 435594 453978
rect 435650 453922 435718 453978
rect 435774 453922 435842 453978
rect 435898 453922 435966 453978
rect 436022 453922 466314 453978
rect 466370 453922 466438 453978
rect 466494 453922 466562 453978
rect 466618 453922 466686 453978
rect 466742 453922 497034 453978
rect 497090 453922 497158 453978
rect 497214 453922 497282 453978
rect 497338 453922 497406 453978
rect 497462 453922 527754 453978
rect 527810 453922 527878 453978
rect 527934 453922 528002 453978
rect 528058 453922 528126 453978
rect 528182 453922 558474 453978
rect 558530 453922 558598 453978
rect 558654 453922 558722 453978
rect 558778 453922 558846 453978
rect 558902 453922 589194 453978
rect 589250 453922 589318 453978
rect 589374 453922 589442 453978
rect 589498 453922 589566 453978
rect 589622 453922 596496 453978
rect 596552 453922 596620 453978
rect 596676 453922 596744 453978
rect 596800 453922 596868 453978
rect 596924 453922 597980 453978
rect -1916 453826 597980 453922
rect -1916 442350 597980 442446
rect -1916 442294 -1820 442350
rect -1764 442294 -1696 442350
rect -1640 442294 -1572 442350
rect -1516 442294 -1448 442350
rect -1392 442294 9234 442350
rect 9290 442294 9358 442350
rect 9414 442294 9482 442350
rect 9538 442294 9606 442350
rect 9662 442294 39954 442350
rect 40010 442294 40078 442350
rect 40134 442294 40202 442350
rect 40258 442294 40326 442350
rect 40382 442294 70674 442350
rect 70730 442294 70798 442350
rect 70854 442294 70922 442350
rect 70978 442294 71046 442350
rect 71102 442294 101394 442350
rect 101450 442294 101518 442350
rect 101574 442294 101642 442350
rect 101698 442294 101766 442350
rect 101822 442294 132114 442350
rect 132170 442294 132238 442350
rect 132294 442294 132362 442350
rect 132418 442294 132486 442350
rect 132542 442294 162834 442350
rect 162890 442294 162958 442350
rect 163014 442294 163082 442350
rect 163138 442294 163206 442350
rect 163262 442294 193554 442350
rect 193610 442294 193678 442350
rect 193734 442294 193802 442350
rect 193858 442294 193926 442350
rect 193982 442294 224274 442350
rect 224330 442294 224398 442350
rect 224454 442294 224522 442350
rect 224578 442294 224646 442350
rect 224702 442294 254994 442350
rect 255050 442294 255118 442350
rect 255174 442294 255242 442350
rect 255298 442294 255366 442350
rect 255422 442294 285714 442350
rect 285770 442294 285838 442350
rect 285894 442294 285962 442350
rect 286018 442294 286086 442350
rect 286142 442294 316434 442350
rect 316490 442294 316558 442350
rect 316614 442294 316682 442350
rect 316738 442294 316806 442350
rect 316862 442294 347154 442350
rect 347210 442294 347278 442350
rect 347334 442294 347402 442350
rect 347458 442294 347526 442350
rect 347582 442294 377874 442350
rect 377930 442294 377998 442350
rect 378054 442294 378122 442350
rect 378178 442294 378246 442350
rect 378302 442294 408594 442350
rect 408650 442294 408718 442350
rect 408774 442294 408842 442350
rect 408898 442294 408966 442350
rect 409022 442294 439314 442350
rect 439370 442294 439438 442350
rect 439494 442294 439562 442350
rect 439618 442294 439686 442350
rect 439742 442294 470034 442350
rect 470090 442294 470158 442350
rect 470214 442294 470282 442350
rect 470338 442294 470406 442350
rect 470462 442294 500754 442350
rect 500810 442294 500878 442350
rect 500934 442294 501002 442350
rect 501058 442294 501126 442350
rect 501182 442294 531474 442350
rect 531530 442294 531598 442350
rect 531654 442294 531722 442350
rect 531778 442294 531846 442350
rect 531902 442294 562194 442350
rect 562250 442294 562318 442350
rect 562374 442294 562442 442350
rect 562498 442294 562566 442350
rect 562622 442294 592914 442350
rect 592970 442294 593038 442350
rect 593094 442294 593162 442350
rect 593218 442294 593286 442350
rect 593342 442294 597456 442350
rect 597512 442294 597580 442350
rect 597636 442294 597704 442350
rect 597760 442294 597828 442350
rect 597884 442294 597980 442350
rect -1916 442226 597980 442294
rect -1916 442170 -1820 442226
rect -1764 442170 -1696 442226
rect -1640 442170 -1572 442226
rect -1516 442170 -1448 442226
rect -1392 442170 9234 442226
rect 9290 442170 9358 442226
rect 9414 442170 9482 442226
rect 9538 442170 9606 442226
rect 9662 442170 39954 442226
rect 40010 442170 40078 442226
rect 40134 442170 40202 442226
rect 40258 442170 40326 442226
rect 40382 442170 70674 442226
rect 70730 442170 70798 442226
rect 70854 442170 70922 442226
rect 70978 442170 71046 442226
rect 71102 442170 101394 442226
rect 101450 442170 101518 442226
rect 101574 442170 101642 442226
rect 101698 442170 101766 442226
rect 101822 442170 132114 442226
rect 132170 442170 132238 442226
rect 132294 442170 132362 442226
rect 132418 442170 132486 442226
rect 132542 442170 162834 442226
rect 162890 442170 162958 442226
rect 163014 442170 163082 442226
rect 163138 442170 163206 442226
rect 163262 442170 193554 442226
rect 193610 442170 193678 442226
rect 193734 442170 193802 442226
rect 193858 442170 193926 442226
rect 193982 442170 224274 442226
rect 224330 442170 224398 442226
rect 224454 442170 224522 442226
rect 224578 442170 224646 442226
rect 224702 442170 254994 442226
rect 255050 442170 255118 442226
rect 255174 442170 255242 442226
rect 255298 442170 255366 442226
rect 255422 442170 285714 442226
rect 285770 442170 285838 442226
rect 285894 442170 285962 442226
rect 286018 442170 286086 442226
rect 286142 442170 316434 442226
rect 316490 442170 316558 442226
rect 316614 442170 316682 442226
rect 316738 442170 316806 442226
rect 316862 442170 347154 442226
rect 347210 442170 347278 442226
rect 347334 442170 347402 442226
rect 347458 442170 347526 442226
rect 347582 442170 377874 442226
rect 377930 442170 377998 442226
rect 378054 442170 378122 442226
rect 378178 442170 378246 442226
rect 378302 442170 408594 442226
rect 408650 442170 408718 442226
rect 408774 442170 408842 442226
rect 408898 442170 408966 442226
rect 409022 442170 439314 442226
rect 439370 442170 439438 442226
rect 439494 442170 439562 442226
rect 439618 442170 439686 442226
rect 439742 442170 470034 442226
rect 470090 442170 470158 442226
rect 470214 442170 470282 442226
rect 470338 442170 470406 442226
rect 470462 442170 500754 442226
rect 500810 442170 500878 442226
rect 500934 442170 501002 442226
rect 501058 442170 501126 442226
rect 501182 442170 531474 442226
rect 531530 442170 531598 442226
rect 531654 442170 531722 442226
rect 531778 442170 531846 442226
rect 531902 442170 562194 442226
rect 562250 442170 562318 442226
rect 562374 442170 562442 442226
rect 562498 442170 562566 442226
rect 562622 442170 592914 442226
rect 592970 442170 593038 442226
rect 593094 442170 593162 442226
rect 593218 442170 593286 442226
rect 593342 442170 597456 442226
rect 597512 442170 597580 442226
rect 597636 442170 597704 442226
rect 597760 442170 597828 442226
rect 597884 442170 597980 442226
rect -1916 442102 597980 442170
rect -1916 442046 -1820 442102
rect -1764 442046 -1696 442102
rect -1640 442046 -1572 442102
rect -1516 442046 -1448 442102
rect -1392 442046 9234 442102
rect 9290 442046 9358 442102
rect 9414 442046 9482 442102
rect 9538 442046 9606 442102
rect 9662 442046 39954 442102
rect 40010 442046 40078 442102
rect 40134 442046 40202 442102
rect 40258 442046 40326 442102
rect 40382 442046 70674 442102
rect 70730 442046 70798 442102
rect 70854 442046 70922 442102
rect 70978 442046 71046 442102
rect 71102 442046 101394 442102
rect 101450 442046 101518 442102
rect 101574 442046 101642 442102
rect 101698 442046 101766 442102
rect 101822 442046 132114 442102
rect 132170 442046 132238 442102
rect 132294 442046 132362 442102
rect 132418 442046 132486 442102
rect 132542 442046 162834 442102
rect 162890 442046 162958 442102
rect 163014 442046 163082 442102
rect 163138 442046 163206 442102
rect 163262 442046 193554 442102
rect 193610 442046 193678 442102
rect 193734 442046 193802 442102
rect 193858 442046 193926 442102
rect 193982 442046 224274 442102
rect 224330 442046 224398 442102
rect 224454 442046 224522 442102
rect 224578 442046 224646 442102
rect 224702 442046 254994 442102
rect 255050 442046 255118 442102
rect 255174 442046 255242 442102
rect 255298 442046 255366 442102
rect 255422 442046 285714 442102
rect 285770 442046 285838 442102
rect 285894 442046 285962 442102
rect 286018 442046 286086 442102
rect 286142 442046 316434 442102
rect 316490 442046 316558 442102
rect 316614 442046 316682 442102
rect 316738 442046 316806 442102
rect 316862 442046 347154 442102
rect 347210 442046 347278 442102
rect 347334 442046 347402 442102
rect 347458 442046 347526 442102
rect 347582 442046 377874 442102
rect 377930 442046 377998 442102
rect 378054 442046 378122 442102
rect 378178 442046 378246 442102
rect 378302 442046 408594 442102
rect 408650 442046 408718 442102
rect 408774 442046 408842 442102
rect 408898 442046 408966 442102
rect 409022 442046 439314 442102
rect 439370 442046 439438 442102
rect 439494 442046 439562 442102
rect 439618 442046 439686 442102
rect 439742 442046 470034 442102
rect 470090 442046 470158 442102
rect 470214 442046 470282 442102
rect 470338 442046 470406 442102
rect 470462 442046 500754 442102
rect 500810 442046 500878 442102
rect 500934 442046 501002 442102
rect 501058 442046 501126 442102
rect 501182 442046 531474 442102
rect 531530 442046 531598 442102
rect 531654 442046 531722 442102
rect 531778 442046 531846 442102
rect 531902 442046 562194 442102
rect 562250 442046 562318 442102
rect 562374 442046 562442 442102
rect 562498 442046 562566 442102
rect 562622 442046 592914 442102
rect 592970 442046 593038 442102
rect 593094 442046 593162 442102
rect 593218 442046 593286 442102
rect 593342 442046 597456 442102
rect 597512 442046 597580 442102
rect 597636 442046 597704 442102
rect 597760 442046 597828 442102
rect 597884 442046 597980 442102
rect -1916 441978 597980 442046
rect -1916 441922 -1820 441978
rect -1764 441922 -1696 441978
rect -1640 441922 -1572 441978
rect -1516 441922 -1448 441978
rect -1392 441922 9234 441978
rect 9290 441922 9358 441978
rect 9414 441922 9482 441978
rect 9538 441922 9606 441978
rect 9662 441922 39954 441978
rect 40010 441922 40078 441978
rect 40134 441922 40202 441978
rect 40258 441922 40326 441978
rect 40382 441922 70674 441978
rect 70730 441922 70798 441978
rect 70854 441922 70922 441978
rect 70978 441922 71046 441978
rect 71102 441922 101394 441978
rect 101450 441922 101518 441978
rect 101574 441922 101642 441978
rect 101698 441922 101766 441978
rect 101822 441922 132114 441978
rect 132170 441922 132238 441978
rect 132294 441922 132362 441978
rect 132418 441922 132486 441978
rect 132542 441922 162834 441978
rect 162890 441922 162958 441978
rect 163014 441922 163082 441978
rect 163138 441922 163206 441978
rect 163262 441922 193554 441978
rect 193610 441922 193678 441978
rect 193734 441922 193802 441978
rect 193858 441922 193926 441978
rect 193982 441922 224274 441978
rect 224330 441922 224398 441978
rect 224454 441922 224522 441978
rect 224578 441922 224646 441978
rect 224702 441922 254994 441978
rect 255050 441922 255118 441978
rect 255174 441922 255242 441978
rect 255298 441922 255366 441978
rect 255422 441922 285714 441978
rect 285770 441922 285838 441978
rect 285894 441922 285962 441978
rect 286018 441922 286086 441978
rect 286142 441922 316434 441978
rect 316490 441922 316558 441978
rect 316614 441922 316682 441978
rect 316738 441922 316806 441978
rect 316862 441922 347154 441978
rect 347210 441922 347278 441978
rect 347334 441922 347402 441978
rect 347458 441922 347526 441978
rect 347582 441922 377874 441978
rect 377930 441922 377998 441978
rect 378054 441922 378122 441978
rect 378178 441922 378246 441978
rect 378302 441922 408594 441978
rect 408650 441922 408718 441978
rect 408774 441922 408842 441978
rect 408898 441922 408966 441978
rect 409022 441922 439314 441978
rect 439370 441922 439438 441978
rect 439494 441922 439562 441978
rect 439618 441922 439686 441978
rect 439742 441922 470034 441978
rect 470090 441922 470158 441978
rect 470214 441922 470282 441978
rect 470338 441922 470406 441978
rect 470462 441922 500754 441978
rect 500810 441922 500878 441978
rect 500934 441922 501002 441978
rect 501058 441922 501126 441978
rect 501182 441922 531474 441978
rect 531530 441922 531598 441978
rect 531654 441922 531722 441978
rect 531778 441922 531846 441978
rect 531902 441922 562194 441978
rect 562250 441922 562318 441978
rect 562374 441922 562442 441978
rect 562498 441922 562566 441978
rect 562622 441922 592914 441978
rect 592970 441922 593038 441978
rect 593094 441922 593162 441978
rect 593218 441922 593286 441978
rect 593342 441922 597456 441978
rect 597512 441922 597580 441978
rect 597636 441922 597704 441978
rect 597760 441922 597828 441978
rect 597884 441922 597980 441978
rect -1916 441826 597980 441922
rect -1916 436350 597980 436446
rect -1916 436294 -860 436350
rect -804 436294 -736 436350
rect -680 436294 -612 436350
rect -556 436294 -488 436350
rect -432 436294 5514 436350
rect 5570 436294 5638 436350
rect 5694 436294 5762 436350
rect 5818 436294 5886 436350
rect 5942 436294 36234 436350
rect 36290 436294 36358 436350
rect 36414 436294 36482 436350
rect 36538 436294 36606 436350
rect 36662 436294 66954 436350
rect 67010 436294 67078 436350
rect 67134 436294 67202 436350
rect 67258 436294 67326 436350
rect 67382 436294 97674 436350
rect 97730 436294 97798 436350
rect 97854 436294 97922 436350
rect 97978 436294 98046 436350
rect 98102 436294 128394 436350
rect 128450 436294 128518 436350
rect 128574 436294 128642 436350
rect 128698 436294 128766 436350
rect 128822 436294 159114 436350
rect 159170 436294 159238 436350
rect 159294 436294 159362 436350
rect 159418 436294 159486 436350
rect 159542 436294 189834 436350
rect 189890 436294 189958 436350
rect 190014 436294 190082 436350
rect 190138 436294 190206 436350
rect 190262 436294 220554 436350
rect 220610 436294 220678 436350
rect 220734 436294 220802 436350
rect 220858 436294 220926 436350
rect 220982 436294 251274 436350
rect 251330 436294 251398 436350
rect 251454 436294 251522 436350
rect 251578 436294 251646 436350
rect 251702 436294 281994 436350
rect 282050 436294 282118 436350
rect 282174 436294 282242 436350
rect 282298 436294 282366 436350
rect 282422 436294 312714 436350
rect 312770 436294 312838 436350
rect 312894 436294 312962 436350
rect 313018 436294 313086 436350
rect 313142 436294 343434 436350
rect 343490 436294 343558 436350
rect 343614 436294 343682 436350
rect 343738 436294 343806 436350
rect 343862 436294 374154 436350
rect 374210 436294 374278 436350
rect 374334 436294 374402 436350
rect 374458 436294 374526 436350
rect 374582 436294 404874 436350
rect 404930 436294 404998 436350
rect 405054 436294 405122 436350
rect 405178 436294 405246 436350
rect 405302 436294 435594 436350
rect 435650 436294 435718 436350
rect 435774 436294 435842 436350
rect 435898 436294 435966 436350
rect 436022 436294 466314 436350
rect 466370 436294 466438 436350
rect 466494 436294 466562 436350
rect 466618 436294 466686 436350
rect 466742 436294 497034 436350
rect 497090 436294 497158 436350
rect 497214 436294 497282 436350
rect 497338 436294 497406 436350
rect 497462 436294 527754 436350
rect 527810 436294 527878 436350
rect 527934 436294 528002 436350
rect 528058 436294 528126 436350
rect 528182 436294 558474 436350
rect 558530 436294 558598 436350
rect 558654 436294 558722 436350
rect 558778 436294 558846 436350
rect 558902 436294 589194 436350
rect 589250 436294 589318 436350
rect 589374 436294 589442 436350
rect 589498 436294 589566 436350
rect 589622 436294 596496 436350
rect 596552 436294 596620 436350
rect 596676 436294 596744 436350
rect 596800 436294 596868 436350
rect 596924 436294 597980 436350
rect -1916 436226 597980 436294
rect -1916 436170 -860 436226
rect -804 436170 -736 436226
rect -680 436170 -612 436226
rect -556 436170 -488 436226
rect -432 436170 5514 436226
rect 5570 436170 5638 436226
rect 5694 436170 5762 436226
rect 5818 436170 5886 436226
rect 5942 436170 36234 436226
rect 36290 436170 36358 436226
rect 36414 436170 36482 436226
rect 36538 436170 36606 436226
rect 36662 436170 66954 436226
rect 67010 436170 67078 436226
rect 67134 436170 67202 436226
rect 67258 436170 67326 436226
rect 67382 436170 97674 436226
rect 97730 436170 97798 436226
rect 97854 436170 97922 436226
rect 97978 436170 98046 436226
rect 98102 436170 128394 436226
rect 128450 436170 128518 436226
rect 128574 436170 128642 436226
rect 128698 436170 128766 436226
rect 128822 436170 159114 436226
rect 159170 436170 159238 436226
rect 159294 436170 159362 436226
rect 159418 436170 159486 436226
rect 159542 436170 189834 436226
rect 189890 436170 189958 436226
rect 190014 436170 190082 436226
rect 190138 436170 190206 436226
rect 190262 436170 220554 436226
rect 220610 436170 220678 436226
rect 220734 436170 220802 436226
rect 220858 436170 220926 436226
rect 220982 436170 251274 436226
rect 251330 436170 251398 436226
rect 251454 436170 251522 436226
rect 251578 436170 251646 436226
rect 251702 436170 281994 436226
rect 282050 436170 282118 436226
rect 282174 436170 282242 436226
rect 282298 436170 282366 436226
rect 282422 436170 312714 436226
rect 312770 436170 312838 436226
rect 312894 436170 312962 436226
rect 313018 436170 313086 436226
rect 313142 436170 343434 436226
rect 343490 436170 343558 436226
rect 343614 436170 343682 436226
rect 343738 436170 343806 436226
rect 343862 436170 374154 436226
rect 374210 436170 374278 436226
rect 374334 436170 374402 436226
rect 374458 436170 374526 436226
rect 374582 436170 404874 436226
rect 404930 436170 404998 436226
rect 405054 436170 405122 436226
rect 405178 436170 405246 436226
rect 405302 436170 435594 436226
rect 435650 436170 435718 436226
rect 435774 436170 435842 436226
rect 435898 436170 435966 436226
rect 436022 436170 466314 436226
rect 466370 436170 466438 436226
rect 466494 436170 466562 436226
rect 466618 436170 466686 436226
rect 466742 436170 497034 436226
rect 497090 436170 497158 436226
rect 497214 436170 497282 436226
rect 497338 436170 497406 436226
rect 497462 436170 527754 436226
rect 527810 436170 527878 436226
rect 527934 436170 528002 436226
rect 528058 436170 528126 436226
rect 528182 436170 558474 436226
rect 558530 436170 558598 436226
rect 558654 436170 558722 436226
rect 558778 436170 558846 436226
rect 558902 436170 589194 436226
rect 589250 436170 589318 436226
rect 589374 436170 589442 436226
rect 589498 436170 589566 436226
rect 589622 436170 596496 436226
rect 596552 436170 596620 436226
rect 596676 436170 596744 436226
rect 596800 436170 596868 436226
rect 596924 436170 597980 436226
rect -1916 436102 597980 436170
rect -1916 436046 -860 436102
rect -804 436046 -736 436102
rect -680 436046 -612 436102
rect -556 436046 -488 436102
rect -432 436046 5514 436102
rect 5570 436046 5638 436102
rect 5694 436046 5762 436102
rect 5818 436046 5886 436102
rect 5942 436046 36234 436102
rect 36290 436046 36358 436102
rect 36414 436046 36482 436102
rect 36538 436046 36606 436102
rect 36662 436046 66954 436102
rect 67010 436046 67078 436102
rect 67134 436046 67202 436102
rect 67258 436046 67326 436102
rect 67382 436046 97674 436102
rect 97730 436046 97798 436102
rect 97854 436046 97922 436102
rect 97978 436046 98046 436102
rect 98102 436046 128394 436102
rect 128450 436046 128518 436102
rect 128574 436046 128642 436102
rect 128698 436046 128766 436102
rect 128822 436046 159114 436102
rect 159170 436046 159238 436102
rect 159294 436046 159362 436102
rect 159418 436046 159486 436102
rect 159542 436046 189834 436102
rect 189890 436046 189958 436102
rect 190014 436046 190082 436102
rect 190138 436046 190206 436102
rect 190262 436046 220554 436102
rect 220610 436046 220678 436102
rect 220734 436046 220802 436102
rect 220858 436046 220926 436102
rect 220982 436046 251274 436102
rect 251330 436046 251398 436102
rect 251454 436046 251522 436102
rect 251578 436046 251646 436102
rect 251702 436046 281994 436102
rect 282050 436046 282118 436102
rect 282174 436046 282242 436102
rect 282298 436046 282366 436102
rect 282422 436046 312714 436102
rect 312770 436046 312838 436102
rect 312894 436046 312962 436102
rect 313018 436046 313086 436102
rect 313142 436046 343434 436102
rect 343490 436046 343558 436102
rect 343614 436046 343682 436102
rect 343738 436046 343806 436102
rect 343862 436046 374154 436102
rect 374210 436046 374278 436102
rect 374334 436046 374402 436102
rect 374458 436046 374526 436102
rect 374582 436046 404874 436102
rect 404930 436046 404998 436102
rect 405054 436046 405122 436102
rect 405178 436046 405246 436102
rect 405302 436046 435594 436102
rect 435650 436046 435718 436102
rect 435774 436046 435842 436102
rect 435898 436046 435966 436102
rect 436022 436046 466314 436102
rect 466370 436046 466438 436102
rect 466494 436046 466562 436102
rect 466618 436046 466686 436102
rect 466742 436046 497034 436102
rect 497090 436046 497158 436102
rect 497214 436046 497282 436102
rect 497338 436046 497406 436102
rect 497462 436046 527754 436102
rect 527810 436046 527878 436102
rect 527934 436046 528002 436102
rect 528058 436046 528126 436102
rect 528182 436046 558474 436102
rect 558530 436046 558598 436102
rect 558654 436046 558722 436102
rect 558778 436046 558846 436102
rect 558902 436046 589194 436102
rect 589250 436046 589318 436102
rect 589374 436046 589442 436102
rect 589498 436046 589566 436102
rect 589622 436046 596496 436102
rect 596552 436046 596620 436102
rect 596676 436046 596744 436102
rect 596800 436046 596868 436102
rect 596924 436046 597980 436102
rect -1916 435978 597980 436046
rect -1916 435922 -860 435978
rect -804 435922 -736 435978
rect -680 435922 -612 435978
rect -556 435922 -488 435978
rect -432 435922 5514 435978
rect 5570 435922 5638 435978
rect 5694 435922 5762 435978
rect 5818 435922 5886 435978
rect 5942 435922 36234 435978
rect 36290 435922 36358 435978
rect 36414 435922 36482 435978
rect 36538 435922 36606 435978
rect 36662 435922 66954 435978
rect 67010 435922 67078 435978
rect 67134 435922 67202 435978
rect 67258 435922 67326 435978
rect 67382 435922 97674 435978
rect 97730 435922 97798 435978
rect 97854 435922 97922 435978
rect 97978 435922 98046 435978
rect 98102 435922 128394 435978
rect 128450 435922 128518 435978
rect 128574 435922 128642 435978
rect 128698 435922 128766 435978
rect 128822 435922 159114 435978
rect 159170 435922 159238 435978
rect 159294 435922 159362 435978
rect 159418 435922 159486 435978
rect 159542 435922 189834 435978
rect 189890 435922 189958 435978
rect 190014 435922 190082 435978
rect 190138 435922 190206 435978
rect 190262 435922 220554 435978
rect 220610 435922 220678 435978
rect 220734 435922 220802 435978
rect 220858 435922 220926 435978
rect 220982 435922 251274 435978
rect 251330 435922 251398 435978
rect 251454 435922 251522 435978
rect 251578 435922 251646 435978
rect 251702 435922 281994 435978
rect 282050 435922 282118 435978
rect 282174 435922 282242 435978
rect 282298 435922 282366 435978
rect 282422 435922 312714 435978
rect 312770 435922 312838 435978
rect 312894 435922 312962 435978
rect 313018 435922 313086 435978
rect 313142 435922 343434 435978
rect 343490 435922 343558 435978
rect 343614 435922 343682 435978
rect 343738 435922 343806 435978
rect 343862 435922 374154 435978
rect 374210 435922 374278 435978
rect 374334 435922 374402 435978
rect 374458 435922 374526 435978
rect 374582 435922 404874 435978
rect 404930 435922 404998 435978
rect 405054 435922 405122 435978
rect 405178 435922 405246 435978
rect 405302 435922 435594 435978
rect 435650 435922 435718 435978
rect 435774 435922 435842 435978
rect 435898 435922 435966 435978
rect 436022 435922 466314 435978
rect 466370 435922 466438 435978
rect 466494 435922 466562 435978
rect 466618 435922 466686 435978
rect 466742 435922 497034 435978
rect 497090 435922 497158 435978
rect 497214 435922 497282 435978
rect 497338 435922 497406 435978
rect 497462 435922 527754 435978
rect 527810 435922 527878 435978
rect 527934 435922 528002 435978
rect 528058 435922 528126 435978
rect 528182 435922 558474 435978
rect 558530 435922 558598 435978
rect 558654 435922 558722 435978
rect 558778 435922 558846 435978
rect 558902 435922 589194 435978
rect 589250 435922 589318 435978
rect 589374 435922 589442 435978
rect 589498 435922 589566 435978
rect 589622 435922 596496 435978
rect 596552 435922 596620 435978
rect 596676 435922 596744 435978
rect 596800 435922 596868 435978
rect 596924 435922 597980 435978
rect -1916 435826 597980 435922
rect -1916 424350 597980 424446
rect -1916 424294 -1820 424350
rect -1764 424294 -1696 424350
rect -1640 424294 -1572 424350
rect -1516 424294 -1448 424350
rect -1392 424294 9234 424350
rect 9290 424294 9358 424350
rect 9414 424294 9482 424350
rect 9538 424294 9606 424350
rect 9662 424294 39954 424350
rect 40010 424294 40078 424350
rect 40134 424294 40202 424350
rect 40258 424294 40326 424350
rect 40382 424294 70674 424350
rect 70730 424294 70798 424350
rect 70854 424294 70922 424350
rect 70978 424294 71046 424350
rect 71102 424294 101394 424350
rect 101450 424294 101518 424350
rect 101574 424294 101642 424350
rect 101698 424294 101766 424350
rect 101822 424294 132114 424350
rect 132170 424294 132238 424350
rect 132294 424294 132362 424350
rect 132418 424294 132486 424350
rect 132542 424294 162834 424350
rect 162890 424294 162958 424350
rect 163014 424294 163082 424350
rect 163138 424294 163206 424350
rect 163262 424294 193554 424350
rect 193610 424294 193678 424350
rect 193734 424294 193802 424350
rect 193858 424294 193926 424350
rect 193982 424294 224274 424350
rect 224330 424294 224398 424350
rect 224454 424294 224522 424350
rect 224578 424294 224646 424350
rect 224702 424294 254994 424350
rect 255050 424294 255118 424350
rect 255174 424294 255242 424350
rect 255298 424294 255366 424350
rect 255422 424294 285714 424350
rect 285770 424294 285838 424350
rect 285894 424294 285962 424350
rect 286018 424294 286086 424350
rect 286142 424294 316434 424350
rect 316490 424294 316558 424350
rect 316614 424294 316682 424350
rect 316738 424294 316806 424350
rect 316862 424294 347154 424350
rect 347210 424294 347278 424350
rect 347334 424294 347402 424350
rect 347458 424294 347526 424350
rect 347582 424294 377874 424350
rect 377930 424294 377998 424350
rect 378054 424294 378122 424350
rect 378178 424294 378246 424350
rect 378302 424294 408594 424350
rect 408650 424294 408718 424350
rect 408774 424294 408842 424350
rect 408898 424294 408966 424350
rect 409022 424294 439314 424350
rect 439370 424294 439438 424350
rect 439494 424294 439562 424350
rect 439618 424294 439686 424350
rect 439742 424294 470034 424350
rect 470090 424294 470158 424350
rect 470214 424294 470282 424350
rect 470338 424294 470406 424350
rect 470462 424294 500754 424350
rect 500810 424294 500878 424350
rect 500934 424294 501002 424350
rect 501058 424294 501126 424350
rect 501182 424294 531474 424350
rect 531530 424294 531598 424350
rect 531654 424294 531722 424350
rect 531778 424294 531846 424350
rect 531902 424294 562194 424350
rect 562250 424294 562318 424350
rect 562374 424294 562442 424350
rect 562498 424294 562566 424350
rect 562622 424294 592914 424350
rect 592970 424294 593038 424350
rect 593094 424294 593162 424350
rect 593218 424294 593286 424350
rect 593342 424294 597456 424350
rect 597512 424294 597580 424350
rect 597636 424294 597704 424350
rect 597760 424294 597828 424350
rect 597884 424294 597980 424350
rect -1916 424226 597980 424294
rect -1916 424170 -1820 424226
rect -1764 424170 -1696 424226
rect -1640 424170 -1572 424226
rect -1516 424170 -1448 424226
rect -1392 424170 9234 424226
rect 9290 424170 9358 424226
rect 9414 424170 9482 424226
rect 9538 424170 9606 424226
rect 9662 424170 39954 424226
rect 40010 424170 40078 424226
rect 40134 424170 40202 424226
rect 40258 424170 40326 424226
rect 40382 424170 70674 424226
rect 70730 424170 70798 424226
rect 70854 424170 70922 424226
rect 70978 424170 71046 424226
rect 71102 424170 101394 424226
rect 101450 424170 101518 424226
rect 101574 424170 101642 424226
rect 101698 424170 101766 424226
rect 101822 424170 132114 424226
rect 132170 424170 132238 424226
rect 132294 424170 132362 424226
rect 132418 424170 132486 424226
rect 132542 424170 162834 424226
rect 162890 424170 162958 424226
rect 163014 424170 163082 424226
rect 163138 424170 163206 424226
rect 163262 424170 193554 424226
rect 193610 424170 193678 424226
rect 193734 424170 193802 424226
rect 193858 424170 193926 424226
rect 193982 424170 224274 424226
rect 224330 424170 224398 424226
rect 224454 424170 224522 424226
rect 224578 424170 224646 424226
rect 224702 424170 254994 424226
rect 255050 424170 255118 424226
rect 255174 424170 255242 424226
rect 255298 424170 255366 424226
rect 255422 424170 285714 424226
rect 285770 424170 285838 424226
rect 285894 424170 285962 424226
rect 286018 424170 286086 424226
rect 286142 424170 316434 424226
rect 316490 424170 316558 424226
rect 316614 424170 316682 424226
rect 316738 424170 316806 424226
rect 316862 424170 347154 424226
rect 347210 424170 347278 424226
rect 347334 424170 347402 424226
rect 347458 424170 347526 424226
rect 347582 424170 377874 424226
rect 377930 424170 377998 424226
rect 378054 424170 378122 424226
rect 378178 424170 378246 424226
rect 378302 424170 408594 424226
rect 408650 424170 408718 424226
rect 408774 424170 408842 424226
rect 408898 424170 408966 424226
rect 409022 424170 439314 424226
rect 439370 424170 439438 424226
rect 439494 424170 439562 424226
rect 439618 424170 439686 424226
rect 439742 424170 470034 424226
rect 470090 424170 470158 424226
rect 470214 424170 470282 424226
rect 470338 424170 470406 424226
rect 470462 424170 500754 424226
rect 500810 424170 500878 424226
rect 500934 424170 501002 424226
rect 501058 424170 501126 424226
rect 501182 424170 531474 424226
rect 531530 424170 531598 424226
rect 531654 424170 531722 424226
rect 531778 424170 531846 424226
rect 531902 424170 562194 424226
rect 562250 424170 562318 424226
rect 562374 424170 562442 424226
rect 562498 424170 562566 424226
rect 562622 424170 592914 424226
rect 592970 424170 593038 424226
rect 593094 424170 593162 424226
rect 593218 424170 593286 424226
rect 593342 424170 597456 424226
rect 597512 424170 597580 424226
rect 597636 424170 597704 424226
rect 597760 424170 597828 424226
rect 597884 424170 597980 424226
rect -1916 424102 597980 424170
rect -1916 424046 -1820 424102
rect -1764 424046 -1696 424102
rect -1640 424046 -1572 424102
rect -1516 424046 -1448 424102
rect -1392 424046 9234 424102
rect 9290 424046 9358 424102
rect 9414 424046 9482 424102
rect 9538 424046 9606 424102
rect 9662 424046 39954 424102
rect 40010 424046 40078 424102
rect 40134 424046 40202 424102
rect 40258 424046 40326 424102
rect 40382 424046 70674 424102
rect 70730 424046 70798 424102
rect 70854 424046 70922 424102
rect 70978 424046 71046 424102
rect 71102 424046 101394 424102
rect 101450 424046 101518 424102
rect 101574 424046 101642 424102
rect 101698 424046 101766 424102
rect 101822 424046 132114 424102
rect 132170 424046 132238 424102
rect 132294 424046 132362 424102
rect 132418 424046 132486 424102
rect 132542 424046 162834 424102
rect 162890 424046 162958 424102
rect 163014 424046 163082 424102
rect 163138 424046 163206 424102
rect 163262 424046 193554 424102
rect 193610 424046 193678 424102
rect 193734 424046 193802 424102
rect 193858 424046 193926 424102
rect 193982 424046 224274 424102
rect 224330 424046 224398 424102
rect 224454 424046 224522 424102
rect 224578 424046 224646 424102
rect 224702 424046 254994 424102
rect 255050 424046 255118 424102
rect 255174 424046 255242 424102
rect 255298 424046 255366 424102
rect 255422 424046 285714 424102
rect 285770 424046 285838 424102
rect 285894 424046 285962 424102
rect 286018 424046 286086 424102
rect 286142 424046 316434 424102
rect 316490 424046 316558 424102
rect 316614 424046 316682 424102
rect 316738 424046 316806 424102
rect 316862 424046 347154 424102
rect 347210 424046 347278 424102
rect 347334 424046 347402 424102
rect 347458 424046 347526 424102
rect 347582 424046 377874 424102
rect 377930 424046 377998 424102
rect 378054 424046 378122 424102
rect 378178 424046 378246 424102
rect 378302 424046 408594 424102
rect 408650 424046 408718 424102
rect 408774 424046 408842 424102
rect 408898 424046 408966 424102
rect 409022 424046 439314 424102
rect 439370 424046 439438 424102
rect 439494 424046 439562 424102
rect 439618 424046 439686 424102
rect 439742 424046 470034 424102
rect 470090 424046 470158 424102
rect 470214 424046 470282 424102
rect 470338 424046 470406 424102
rect 470462 424046 500754 424102
rect 500810 424046 500878 424102
rect 500934 424046 501002 424102
rect 501058 424046 501126 424102
rect 501182 424046 531474 424102
rect 531530 424046 531598 424102
rect 531654 424046 531722 424102
rect 531778 424046 531846 424102
rect 531902 424046 562194 424102
rect 562250 424046 562318 424102
rect 562374 424046 562442 424102
rect 562498 424046 562566 424102
rect 562622 424046 592914 424102
rect 592970 424046 593038 424102
rect 593094 424046 593162 424102
rect 593218 424046 593286 424102
rect 593342 424046 597456 424102
rect 597512 424046 597580 424102
rect 597636 424046 597704 424102
rect 597760 424046 597828 424102
rect 597884 424046 597980 424102
rect -1916 423978 597980 424046
rect -1916 423922 -1820 423978
rect -1764 423922 -1696 423978
rect -1640 423922 -1572 423978
rect -1516 423922 -1448 423978
rect -1392 423922 9234 423978
rect 9290 423922 9358 423978
rect 9414 423922 9482 423978
rect 9538 423922 9606 423978
rect 9662 423922 39954 423978
rect 40010 423922 40078 423978
rect 40134 423922 40202 423978
rect 40258 423922 40326 423978
rect 40382 423922 70674 423978
rect 70730 423922 70798 423978
rect 70854 423922 70922 423978
rect 70978 423922 71046 423978
rect 71102 423922 101394 423978
rect 101450 423922 101518 423978
rect 101574 423922 101642 423978
rect 101698 423922 101766 423978
rect 101822 423922 132114 423978
rect 132170 423922 132238 423978
rect 132294 423922 132362 423978
rect 132418 423922 132486 423978
rect 132542 423922 162834 423978
rect 162890 423922 162958 423978
rect 163014 423922 163082 423978
rect 163138 423922 163206 423978
rect 163262 423922 193554 423978
rect 193610 423922 193678 423978
rect 193734 423922 193802 423978
rect 193858 423922 193926 423978
rect 193982 423922 224274 423978
rect 224330 423922 224398 423978
rect 224454 423922 224522 423978
rect 224578 423922 224646 423978
rect 224702 423922 254994 423978
rect 255050 423922 255118 423978
rect 255174 423922 255242 423978
rect 255298 423922 255366 423978
rect 255422 423922 285714 423978
rect 285770 423922 285838 423978
rect 285894 423922 285962 423978
rect 286018 423922 286086 423978
rect 286142 423922 316434 423978
rect 316490 423922 316558 423978
rect 316614 423922 316682 423978
rect 316738 423922 316806 423978
rect 316862 423922 347154 423978
rect 347210 423922 347278 423978
rect 347334 423922 347402 423978
rect 347458 423922 347526 423978
rect 347582 423922 377874 423978
rect 377930 423922 377998 423978
rect 378054 423922 378122 423978
rect 378178 423922 378246 423978
rect 378302 423922 408594 423978
rect 408650 423922 408718 423978
rect 408774 423922 408842 423978
rect 408898 423922 408966 423978
rect 409022 423922 439314 423978
rect 439370 423922 439438 423978
rect 439494 423922 439562 423978
rect 439618 423922 439686 423978
rect 439742 423922 470034 423978
rect 470090 423922 470158 423978
rect 470214 423922 470282 423978
rect 470338 423922 470406 423978
rect 470462 423922 500754 423978
rect 500810 423922 500878 423978
rect 500934 423922 501002 423978
rect 501058 423922 501126 423978
rect 501182 423922 531474 423978
rect 531530 423922 531598 423978
rect 531654 423922 531722 423978
rect 531778 423922 531846 423978
rect 531902 423922 562194 423978
rect 562250 423922 562318 423978
rect 562374 423922 562442 423978
rect 562498 423922 562566 423978
rect 562622 423922 592914 423978
rect 592970 423922 593038 423978
rect 593094 423922 593162 423978
rect 593218 423922 593286 423978
rect 593342 423922 597456 423978
rect 597512 423922 597580 423978
rect 597636 423922 597704 423978
rect 597760 423922 597828 423978
rect 597884 423922 597980 423978
rect -1916 423826 597980 423922
rect -1916 418350 597980 418446
rect -1916 418294 -860 418350
rect -804 418294 -736 418350
rect -680 418294 -612 418350
rect -556 418294 -488 418350
rect -432 418294 5514 418350
rect 5570 418294 5638 418350
rect 5694 418294 5762 418350
rect 5818 418294 5886 418350
rect 5942 418294 36234 418350
rect 36290 418294 36358 418350
rect 36414 418294 36482 418350
rect 36538 418294 36606 418350
rect 36662 418294 66954 418350
rect 67010 418294 67078 418350
rect 67134 418294 67202 418350
rect 67258 418294 67326 418350
rect 67382 418294 97674 418350
rect 97730 418294 97798 418350
rect 97854 418294 97922 418350
rect 97978 418294 98046 418350
rect 98102 418294 128394 418350
rect 128450 418294 128518 418350
rect 128574 418294 128642 418350
rect 128698 418294 128766 418350
rect 128822 418294 159114 418350
rect 159170 418294 159238 418350
rect 159294 418294 159362 418350
rect 159418 418294 159486 418350
rect 159542 418294 189834 418350
rect 189890 418294 189958 418350
rect 190014 418294 190082 418350
rect 190138 418294 190206 418350
rect 190262 418294 220554 418350
rect 220610 418294 220678 418350
rect 220734 418294 220802 418350
rect 220858 418294 220926 418350
rect 220982 418294 251274 418350
rect 251330 418294 251398 418350
rect 251454 418294 251522 418350
rect 251578 418294 251646 418350
rect 251702 418294 281994 418350
rect 282050 418294 282118 418350
rect 282174 418294 282242 418350
rect 282298 418294 282366 418350
rect 282422 418294 312714 418350
rect 312770 418294 312838 418350
rect 312894 418294 312962 418350
rect 313018 418294 313086 418350
rect 313142 418294 343434 418350
rect 343490 418294 343558 418350
rect 343614 418294 343682 418350
rect 343738 418294 343806 418350
rect 343862 418294 374154 418350
rect 374210 418294 374278 418350
rect 374334 418294 374402 418350
rect 374458 418294 374526 418350
rect 374582 418294 404874 418350
rect 404930 418294 404998 418350
rect 405054 418294 405122 418350
rect 405178 418294 405246 418350
rect 405302 418294 435594 418350
rect 435650 418294 435718 418350
rect 435774 418294 435842 418350
rect 435898 418294 435966 418350
rect 436022 418294 466314 418350
rect 466370 418294 466438 418350
rect 466494 418294 466562 418350
rect 466618 418294 466686 418350
rect 466742 418294 497034 418350
rect 497090 418294 497158 418350
rect 497214 418294 497282 418350
rect 497338 418294 497406 418350
rect 497462 418294 527754 418350
rect 527810 418294 527878 418350
rect 527934 418294 528002 418350
rect 528058 418294 528126 418350
rect 528182 418294 558474 418350
rect 558530 418294 558598 418350
rect 558654 418294 558722 418350
rect 558778 418294 558846 418350
rect 558902 418294 589194 418350
rect 589250 418294 589318 418350
rect 589374 418294 589442 418350
rect 589498 418294 589566 418350
rect 589622 418294 596496 418350
rect 596552 418294 596620 418350
rect 596676 418294 596744 418350
rect 596800 418294 596868 418350
rect 596924 418294 597980 418350
rect -1916 418226 597980 418294
rect -1916 418170 -860 418226
rect -804 418170 -736 418226
rect -680 418170 -612 418226
rect -556 418170 -488 418226
rect -432 418170 5514 418226
rect 5570 418170 5638 418226
rect 5694 418170 5762 418226
rect 5818 418170 5886 418226
rect 5942 418170 36234 418226
rect 36290 418170 36358 418226
rect 36414 418170 36482 418226
rect 36538 418170 36606 418226
rect 36662 418170 66954 418226
rect 67010 418170 67078 418226
rect 67134 418170 67202 418226
rect 67258 418170 67326 418226
rect 67382 418170 97674 418226
rect 97730 418170 97798 418226
rect 97854 418170 97922 418226
rect 97978 418170 98046 418226
rect 98102 418170 128394 418226
rect 128450 418170 128518 418226
rect 128574 418170 128642 418226
rect 128698 418170 128766 418226
rect 128822 418170 159114 418226
rect 159170 418170 159238 418226
rect 159294 418170 159362 418226
rect 159418 418170 159486 418226
rect 159542 418170 189834 418226
rect 189890 418170 189958 418226
rect 190014 418170 190082 418226
rect 190138 418170 190206 418226
rect 190262 418170 220554 418226
rect 220610 418170 220678 418226
rect 220734 418170 220802 418226
rect 220858 418170 220926 418226
rect 220982 418170 251274 418226
rect 251330 418170 251398 418226
rect 251454 418170 251522 418226
rect 251578 418170 251646 418226
rect 251702 418170 281994 418226
rect 282050 418170 282118 418226
rect 282174 418170 282242 418226
rect 282298 418170 282366 418226
rect 282422 418170 312714 418226
rect 312770 418170 312838 418226
rect 312894 418170 312962 418226
rect 313018 418170 313086 418226
rect 313142 418170 343434 418226
rect 343490 418170 343558 418226
rect 343614 418170 343682 418226
rect 343738 418170 343806 418226
rect 343862 418170 374154 418226
rect 374210 418170 374278 418226
rect 374334 418170 374402 418226
rect 374458 418170 374526 418226
rect 374582 418170 404874 418226
rect 404930 418170 404998 418226
rect 405054 418170 405122 418226
rect 405178 418170 405246 418226
rect 405302 418170 435594 418226
rect 435650 418170 435718 418226
rect 435774 418170 435842 418226
rect 435898 418170 435966 418226
rect 436022 418170 466314 418226
rect 466370 418170 466438 418226
rect 466494 418170 466562 418226
rect 466618 418170 466686 418226
rect 466742 418170 497034 418226
rect 497090 418170 497158 418226
rect 497214 418170 497282 418226
rect 497338 418170 497406 418226
rect 497462 418170 527754 418226
rect 527810 418170 527878 418226
rect 527934 418170 528002 418226
rect 528058 418170 528126 418226
rect 528182 418170 558474 418226
rect 558530 418170 558598 418226
rect 558654 418170 558722 418226
rect 558778 418170 558846 418226
rect 558902 418170 589194 418226
rect 589250 418170 589318 418226
rect 589374 418170 589442 418226
rect 589498 418170 589566 418226
rect 589622 418170 596496 418226
rect 596552 418170 596620 418226
rect 596676 418170 596744 418226
rect 596800 418170 596868 418226
rect 596924 418170 597980 418226
rect -1916 418102 597980 418170
rect -1916 418046 -860 418102
rect -804 418046 -736 418102
rect -680 418046 -612 418102
rect -556 418046 -488 418102
rect -432 418046 5514 418102
rect 5570 418046 5638 418102
rect 5694 418046 5762 418102
rect 5818 418046 5886 418102
rect 5942 418046 36234 418102
rect 36290 418046 36358 418102
rect 36414 418046 36482 418102
rect 36538 418046 36606 418102
rect 36662 418046 66954 418102
rect 67010 418046 67078 418102
rect 67134 418046 67202 418102
rect 67258 418046 67326 418102
rect 67382 418046 97674 418102
rect 97730 418046 97798 418102
rect 97854 418046 97922 418102
rect 97978 418046 98046 418102
rect 98102 418046 128394 418102
rect 128450 418046 128518 418102
rect 128574 418046 128642 418102
rect 128698 418046 128766 418102
rect 128822 418046 159114 418102
rect 159170 418046 159238 418102
rect 159294 418046 159362 418102
rect 159418 418046 159486 418102
rect 159542 418046 189834 418102
rect 189890 418046 189958 418102
rect 190014 418046 190082 418102
rect 190138 418046 190206 418102
rect 190262 418046 220554 418102
rect 220610 418046 220678 418102
rect 220734 418046 220802 418102
rect 220858 418046 220926 418102
rect 220982 418046 251274 418102
rect 251330 418046 251398 418102
rect 251454 418046 251522 418102
rect 251578 418046 251646 418102
rect 251702 418046 281994 418102
rect 282050 418046 282118 418102
rect 282174 418046 282242 418102
rect 282298 418046 282366 418102
rect 282422 418046 312714 418102
rect 312770 418046 312838 418102
rect 312894 418046 312962 418102
rect 313018 418046 313086 418102
rect 313142 418046 343434 418102
rect 343490 418046 343558 418102
rect 343614 418046 343682 418102
rect 343738 418046 343806 418102
rect 343862 418046 374154 418102
rect 374210 418046 374278 418102
rect 374334 418046 374402 418102
rect 374458 418046 374526 418102
rect 374582 418046 404874 418102
rect 404930 418046 404998 418102
rect 405054 418046 405122 418102
rect 405178 418046 405246 418102
rect 405302 418046 435594 418102
rect 435650 418046 435718 418102
rect 435774 418046 435842 418102
rect 435898 418046 435966 418102
rect 436022 418046 466314 418102
rect 466370 418046 466438 418102
rect 466494 418046 466562 418102
rect 466618 418046 466686 418102
rect 466742 418046 497034 418102
rect 497090 418046 497158 418102
rect 497214 418046 497282 418102
rect 497338 418046 497406 418102
rect 497462 418046 527754 418102
rect 527810 418046 527878 418102
rect 527934 418046 528002 418102
rect 528058 418046 528126 418102
rect 528182 418046 558474 418102
rect 558530 418046 558598 418102
rect 558654 418046 558722 418102
rect 558778 418046 558846 418102
rect 558902 418046 589194 418102
rect 589250 418046 589318 418102
rect 589374 418046 589442 418102
rect 589498 418046 589566 418102
rect 589622 418046 596496 418102
rect 596552 418046 596620 418102
rect 596676 418046 596744 418102
rect 596800 418046 596868 418102
rect 596924 418046 597980 418102
rect -1916 417978 597980 418046
rect -1916 417922 -860 417978
rect -804 417922 -736 417978
rect -680 417922 -612 417978
rect -556 417922 -488 417978
rect -432 417922 5514 417978
rect 5570 417922 5638 417978
rect 5694 417922 5762 417978
rect 5818 417922 5886 417978
rect 5942 417922 36234 417978
rect 36290 417922 36358 417978
rect 36414 417922 36482 417978
rect 36538 417922 36606 417978
rect 36662 417922 66954 417978
rect 67010 417922 67078 417978
rect 67134 417922 67202 417978
rect 67258 417922 67326 417978
rect 67382 417922 97674 417978
rect 97730 417922 97798 417978
rect 97854 417922 97922 417978
rect 97978 417922 98046 417978
rect 98102 417922 128394 417978
rect 128450 417922 128518 417978
rect 128574 417922 128642 417978
rect 128698 417922 128766 417978
rect 128822 417922 159114 417978
rect 159170 417922 159238 417978
rect 159294 417922 159362 417978
rect 159418 417922 159486 417978
rect 159542 417922 189834 417978
rect 189890 417922 189958 417978
rect 190014 417922 190082 417978
rect 190138 417922 190206 417978
rect 190262 417922 220554 417978
rect 220610 417922 220678 417978
rect 220734 417922 220802 417978
rect 220858 417922 220926 417978
rect 220982 417922 251274 417978
rect 251330 417922 251398 417978
rect 251454 417922 251522 417978
rect 251578 417922 251646 417978
rect 251702 417922 281994 417978
rect 282050 417922 282118 417978
rect 282174 417922 282242 417978
rect 282298 417922 282366 417978
rect 282422 417922 312714 417978
rect 312770 417922 312838 417978
rect 312894 417922 312962 417978
rect 313018 417922 313086 417978
rect 313142 417922 343434 417978
rect 343490 417922 343558 417978
rect 343614 417922 343682 417978
rect 343738 417922 343806 417978
rect 343862 417922 374154 417978
rect 374210 417922 374278 417978
rect 374334 417922 374402 417978
rect 374458 417922 374526 417978
rect 374582 417922 404874 417978
rect 404930 417922 404998 417978
rect 405054 417922 405122 417978
rect 405178 417922 405246 417978
rect 405302 417922 435594 417978
rect 435650 417922 435718 417978
rect 435774 417922 435842 417978
rect 435898 417922 435966 417978
rect 436022 417922 466314 417978
rect 466370 417922 466438 417978
rect 466494 417922 466562 417978
rect 466618 417922 466686 417978
rect 466742 417922 497034 417978
rect 497090 417922 497158 417978
rect 497214 417922 497282 417978
rect 497338 417922 497406 417978
rect 497462 417922 527754 417978
rect 527810 417922 527878 417978
rect 527934 417922 528002 417978
rect 528058 417922 528126 417978
rect 528182 417922 558474 417978
rect 558530 417922 558598 417978
rect 558654 417922 558722 417978
rect 558778 417922 558846 417978
rect 558902 417922 589194 417978
rect 589250 417922 589318 417978
rect 589374 417922 589442 417978
rect 589498 417922 589566 417978
rect 589622 417922 596496 417978
rect 596552 417922 596620 417978
rect 596676 417922 596744 417978
rect 596800 417922 596868 417978
rect 596924 417922 597980 417978
rect -1916 417826 597980 417922
rect -1916 406350 597980 406446
rect -1916 406294 -1820 406350
rect -1764 406294 -1696 406350
rect -1640 406294 -1572 406350
rect -1516 406294 -1448 406350
rect -1392 406294 9234 406350
rect 9290 406294 9358 406350
rect 9414 406294 9482 406350
rect 9538 406294 9606 406350
rect 9662 406294 39954 406350
rect 40010 406294 40078 406350
rect 40134 406294 40202 406350
rect 40258 406294 40326 406350
rect 40382 406294 70674 406350
rect 70730 406294 70798 406350
rect 70854 406294 70922 406350
rect 70978 406294 71046 406350
rect 71102 406294 101394 406350
rect 101450 406294 101518 406350
rect 101574 406294 101642 406350
rect 101698 406294 101766 406350
rect 101822 406294 132114 406350
rect 132170 406294 132238 406350
rect 132294 406294 132362 406350
rect 132418 406294 132486 406350
rect 132542 406294 162834 406350
rect 162890 406294 162958 406350
rect 163014 406294 163082 406350
rect 163138 406294 163206 406350
rect 163262 406294 193554 406350
rect 193610 406294 193678 406350
rect 193734 406294 193802 406350
rect 193858 406294 193926 406350
rect 193982 406294 224274 406350
rect 224330 406294 224398 406350
rect 224454 406294 224522 406350
rect 224578 406294 224646 406350
rect 224702 406294 254994 406350
rect 255050 406294 255118 406350
rect 255174 406294 255242 406350
rect 255298 406294 255366 406350
rect 255422 406294 285714 406350
rect 285770 406294 285838 406350
rect 285894 406294 285962 406350
rect 286018 406294 286086 406350
rect 286142 406294 316434 406350
rect 316490 406294 316558 406350
rect 316614 406294 316682 406350
rect 316738 406294 316806 406350
rect 316862 406294 347154 406350
rect 347210 406294 347278 406350
rect 347334 406294 347402 406350
rect 347458 406294 347526 406350
rect 347582 406294 377874 406350
rect 377930 406294 377998 406350
rect 378054 406294 378122 406350
rect 378178 406294 378246 406350
rect 378302 406294 408594 406350
rect 408650 406294 408718 406350
rect 408774 406294 408842 406350
rect 408898 406294 408966 406350
rect 409022 406294 439314 406350
rect 439370 406294 439438 406350
rect 439494 406294 439562 406350
rect 439618 406294 439686 406350
rect 439742 406294 470034 406350
rect 470090 406294 470158 406350
rect 470214 406294 470282 406350
rect 470338 406294 470406 406350
rect 470462 406294 500754 406350
rect 500810 406294 500878 406350
rect 500934 406294 501002 406350
rect 501058 406294 501126 406350
rect 501182 406294 531474 406350
rect 531530 406294 531598 406350
rect 531654 406294 531722 406350
rect 531778 406294 531846 406350
rect 531902 406294 562194 406350
rect 562250 406294 562318 406350
rect 562374 406294 562442 406350
rect 562498 406294 562566 406350
rect 562622 406294 592914 406350
rect 592970 406294 593038 406350
rect 593094 406294 593162 406350
rect 593218 406294 593286 406350
rect 593342 406294 597456 406350
rect 597512 406294 597580 406350
rect 597636 406294 597704 406350
rect 597760 406294 597828 406350
rect 597884 406294 597980 406350
rect -1916 406226 597980 406294
rect -1916 406170 -1820 406226
rect -1764 406170 -1696 406226
rect -1640 406170 -1572 406226
rect -1516 406170 -1448 406226
rect -1392 406170 9234 406226
rect 9290 406170 9358 406226
rect 9414 406170 9482 406226
rect 9538 406170 9606 406226
rect 9662 406170 39954 406226
rect 40010 406170 40078 406226
rect 40134 406170 40202 406226
rect 40258 406170 40326 406226
rect 40382 406170 70674 406226
rect 70730 406170 70798 406226
rect 70854 406170 70922 406226
rect 70978 406170 71046 406226
rect 71102 406170 101394 406226
rect 101450 406170 101518 406226
rect 101574 406170 101642 406226
rect 101698 406170 101766 406226
rect 101822 406170 132114 406226
rect 132170 406170 132238 406226
rect 132294 406170 132362 406226
rect 132418 406170 132486 406226
rect 132542 406170 162834 406226
rect 162890 406170 162958 406226
rect 163014 406170 163082 406226
rect 163138 406170 163206 406226
rect 163262 406170 193554 406226
rect 193610 406170 193678 406226
rect 193734 406170 193802 406226
rect 193858 406170 193926 406226
rect 193982 406170 224274 406226
rect 224330 406170 224398 406226
rect 224454 406170 224522 406226
rect 224578 406170 224646 406226
rect 224702 406170 254994 406226
rect 255050 406170 255118 406226
rect 255174 406170 255242 406226
rect 255298 406170 255366 406226
rect 255422 406170 285714 406226
rect 285770 406170 285838 406226
rect 285894 406170 285962 406226
rect 286018 406170 286086 406226
rect 286142 406170 316434 406226
rect 316490 406170 316558 406226
rect 316614 406170 316682 406226
rect 316738 406170 316806 406226
rect 316862 406170 347154 406226
rect 347210 406170 347278 406226
rect 347334 406170 347402 406226
rect 347458 406170 347526 406226
rect 347582 406170 377874 406226
rect 377930 406170 377998 406226
rect 378054 406170 378122 406226
rect 378178 406170 378246 406226
rect 378302 406170 408594 406226
rect 408650 406170 408718 406226
rect 408774 406170 408842 406226
rect 408898 406170 408966 406226
rect 409022 406170 439314 406226
rect 439370 406170 439438 406226
rect 439494 406170 439562 406226
rect 439618 406170 439686 406226
rect 439742 406170 470034 406226
rect 470090 406170 470158 406226
rect 470214 406170 470282 406226
rect 470338 406170 470406 406226
rect 470462 406170 500754 406226
rect 500810 406170 500878 406226
rect 500934 406170 501002 406226
rect 501058 406170 501126 406226
rect 501182 406170 531474 406226
rect 531530 406170 531598 406226
rect 531654 406170 531722 406226
rect 531778 406170 531846 406226
rect 531902 406170 562194 406226
rect 562250 406170 562318 406226
rect 562374 406170 562442 406226
rect 562498 406170 562566 406226
rect 562622 406170 592914 406226
rect 592970 406170 593038 406226
rect 593094 406170 593162 406226
rect 593218 406170 593286 406226
rect 593342 406170 597456 406226
rect 597512 406170 597580 406226
rect 597636 406170 597704 406226
rect 597760 406170 597828 406226
rect 597884 406170 597980 406226
rect -1916 406102 597980 406170
rect -1916 406046 -1820 406102
rect -1764 406046 -1696 406102
rect -1640 406046 -1572 406102
rect -1516 406046 -1448 406102
rect -1392 406046 9234 406102
rect 9290 406046 9358 406102
rect 9414 406046 9482 406102
rect 9538 406046 9606 406102
rect 9662 406046 39954 406102
rect 40010 406046 40078 406102
rect 40134 406046 40202 406102
rect 40258 406046 40326 406102
rect 40382 406046 70674 406102
rect 70730 406046 70798 406102
rect 70854 406046 70922 406102
rect 70978 406046 71046 406102
rect 71102 406046 101394 406102
rect 101450 406046 101518 406102
rect 101574 406046 101642 406102
rect 101698 406046 101766 406102
rect 101822 406046 132114 406102
rect 132170 406046 132238 406102
rect 132294 406046 132362 406102
rect 132418 406046 132486 406102
rect 132542 406046 162834 406102
rect 162890 406046 162958 406102
rect 163014 406046 163082 406102
rect 163138 406046 163206 406102
rect 163262 406046 193554 406102
rect 193610 406046 193678 406102
rect 193734 406046 193802 406102
rect 193858 406046 193926 406102
rect 193982 406046 224274 406102
rect 224330 406046 224398 406102
rect 224454 406046 224522 406102
rect 224578 406046 224646 406102
rect 224702 406046 254994 406102
rect 255050 406046 255118 406102
rect 255174 406046 255242 406102
rect 255298 406046 255366 406102
rect 255422 406046 285714 406102
rect 285770 406046 285838 406102
rect 285894 406046 285962 406102
rect 286018 406046 286086 406102
rect 286142 406046 316434 406102
rect 316490 406046 316558 406102
rect 316614 406046 316682 406102
rect 316738 406046 316806 406102
rect 316862 406046 347154 406102
rect 347210 406046 347278 406102
rect 347334 406046 347402 406102
rect 347458 406046 347526 406102
rect 347582 406046 377874 406102
rect 377930 406046 377998 406102
rect 378054 406046 378122 406102
rect 378178 406046 378246 406102
rect 378302 406046 408594 406102
rect 408650 406046 408718 406102
rect 408774 406046 408842 406102
rect 408898 406046 408966 406102
rect 409022 406046 439314 406102
rect 439370 406046 439438 406102
rect 439494 406046 439562 406102
rect 439618 406046 439686 406102
rect 439742 406046 470034 406102
rect 470090 406046 470158 406102
rect 470214 406046 470282 406102
rect 470338 406046 470406 406102
rect 470462 406046 500754 406102
rect 500810 406046 500878 406102
rect 500934 406046 501002 406102
rect 501058 406046 501126 406102
rect 501182 406046 531474 406102
rect 531530 406046 531598 406102
rect 531654 406046 531722 406102
rect 531778 406046 531846 406102
rect 531902 406046 562194 406102
rect 562250 406046 562318 406102
rect 562374 406046 562442 406102
rect 562498 406046 562566 406102
rect 562622 406046 592914 406102
rect 592970 406046 593038 406102
rect 593094 406046 593162 406102
rect 593218 406046 593286 406102
rect 593342 406046 597456 406102
rect 597512 406046 597580 406102
rect 597636 406046 597704 406102
rect 597760 406046 597828 406102
rect 597884 406046 597980 406102
rect -1916 405978 597980 406046
rect -1916 405922 -1820 405978
rect -1764 405922 -1696 405978
rect -1640 405922 -1572 405978
rect -1516 405922 -1448 405978
rect -1392 405922 9234 405978
rect 9290 405922 9358 405978
rect 9414 405922 9482 405978
rect 9538 405922 9606 405978
rect 9662 405922 39954 405978
rect 40010 405922 40078 405978
rect 40134 405922 40202 405978
rect 40258 405922 40326 405978
rect 40382 405922 70674 405978
rect 70730 405922 70798 405978
rect 70854 405922 70922 405978
rect 70978 405922 71046 405978
rect 71102 405922 101394 405978
rect 101450 405922 101518 405978
rect 101574 405922 101642 405978
rect 101698 405922 101766 405978
rect 101822 405922 132114 405978
rect 132170 405922 132238 405978
rect 132294 405922 132362 405978
rect 132418 405922 132486 405978
rect 132542 405922 162834 405978
rect 162890 405922 162958 405978
rect 163014 405922 163082 405978
rect 163138 405922 163206 405978
rect 163262 405922 193554 405978
rect 193610 405922 193678 405978
rect 193734 405922 193802 405978
rect 193858 405922 193926 405978
rect 193982 405922 224274 405978
rect 224330 405922 224398 405978
rect 224454 405922 224522 405978
rect 224578 405922 224646 405978
rect 224702 405922 254994 405978
rect 255050 405922 255118 405978
rect 255174 405922 255242 405978
rect 255298 405922 255366 405978
rect 255422 405922 285714 405978
rect 285770 405922 285838 405978
rect 285894 405922 285962 405978
rect 286018 405922 286086 405978
rect 286142 405922 316434 405978
rect 316490 405922 316558 405978
rect 316614 405922 316682 405978
rect 316738 405922 316806 405978
rect 316862 405922 347154 405978
rect 347210 405922 347278 405978
rect 347334 405922 347402 405978
rect 347458 405922 347526 405978
rect 347582 405922 377874 405978
rect 377930 405922 377998 405978
rect 378054 405922 378122 405978
rect 378178 405922 378246 405978
rect 378302 405922 408594 405978
rect 408650 405922 408718 405978
rect 408774 405922 408842 405978
rect 408898 405922 408966 405978
rect 409022 405922 439314 405978
rect 439370 405922 439438 405978
rect 439494 405922 439562 405978
rect 439618 405922 439686 405978
rect 439742 405922 470034 405978
rect 470090 405922 470158 405978
rect 470214 405922 470282 405978
rect 470338 405922 470406 405978
rect 470462 405922 500754 405978
rect 500810 405922 500878 405978
rect 500934 405922 501002 405978
rect 501058 405922 501126 405978
rect 501182 405922 531474 405978
rect 531530 405922 531598 405978
rect 531654 405922 531722 405978
rect 531778 405922 531846 405978
rect 531902 405922 562194 405978
rect 562250 405922 562318 405978
rect 562374 405922 562442 405978
rect 562498 405922 562566 405978
rect 562622 405922 592914 405978
rect 592970 405922 593038 405978
rect 593094 405922 593162 405978
rect 593218 405922 593286 405978
rect 593342 405922 597456 405978
rect 597512 405922 597580 405978
rect 597636 405922 597704 405978
rect 597760 405922 597828 405978
rect 597884 405922 597980 405978
rect -1916 405826 597980 405922
rect -1916 400350 597980 400446
rect -1916 400294 -860 400350
rect -804 400294 -736 400350
rect -680 400294 -612 400350
rect -556 400294 -488 400350
rect -432 400294 5514 400350
rect 5570 400294 5638 400350
rect 5694 400294 5762 400350
rect 5818 400294 5886 400350
rect 5942 400294 36234 400350
rect 36290 400294 36358 400350
rect 36414 400294 36482 400350
rect 36538 400294 36606 400350
rect 36662 400294 66954 400350
rect 67010 400294 67078 400350
rect 67134 400294 67202 400350
rect 67258 400294 67326 400350
rect 67382 400294 97674 400350
rect 97730 400294 97798 400350
rect 97854 400294 97922 400350
rect 97978 400294 98046 400350
rect 98102 400294 128394 400350
rect 128450 400294 128518 400350
rect 128574 400294 128642 400350
rect 128698 400294 128766 400350
rect 128822 400294 159114 400350
rect 159170 400294 159238 400350
rect 159294 400294 159362 400350
rect 159418 400294 159486 400350
rect 159542 400294 189834 400350
rect 189890 400294 189958 400350
rect 190014 400294 190082 400350
rect 190138 400294 190206 400350
rect 190262 400294 220554 400350
rect 220610 400294 220678 400350
rect 220734 400294 220802 400350
rect 220858 400294 220926 400350
rect 220982 400294 251274 400350
rect 251330 400294 251398 400350
rect 251454 400294 251522 400350
rect 251578 400294 251646 400350
rect 251702 400294 281994 400350
rect 282050 400294 282118 400350
rect 282174 400294 282242 400350
rect 282298 400294 282366 400350
rect 282422 400294 312714 400350
rect 312770 400294 312838 400350
rect 312894 400294 312962 400350
rect 313018 400294 313086 400350
rect 313142 400294 343434 400350
rect 343490 400294 343558 400350
rect 343614 400294 343682 400350
rect 343738 400294 343806 400350
rect 343862 400294 374154 400350
rect 374210 400294 374278 400350
rect 374334 400294 374402 400350
rect 374458 400294 374526 400350
rect 374582 400294 404874 400350
rect 404930 400294 404998 400350
rect 405054 400294 405122 400350
rect 405178 400294 405246 400350
rect 405302 400294 435594 400350
rect 435650 400294 435718 400350
rect 435774 400294 435842 400350
rect 435898 400294 435966 400350
rect 436022 400294 466314 400350
rect 466370 400294 466438 400350
rect 466494 400294 466562 400350
rect 466618 400294 466686 400350
rect 466742 400294 497034 400350
rect 497090 400294 497158 400350
rect 497214 400294 497282 400350
rect 497338 400294 497406 400350
rect 497462 400294 527754 400350
rect 527810 400294 527878 400350
rect 527934 400294 528002 400350
rect 528058 400294 528126 400350
rect 528182 400294 558474 400350
rect 558530 400294 558598 400350
rect 558654 400294 558722 400350
rect 558778 400294 558846 400350
rect 558902 400294 589194 400350
rect 589250 400294 589318 400350
rect 589374 400294 589442 400350
rect 589498 400294 589566 400350
rect 589622 400294 596496 400350
rect 596552 400294 596620 400350
rect 596676 400294 596744 400350
rect 596800 400294 596868 400350
rect 596924 400294 597980 400350
rect -1916 400226 597980 400294
rect -1916 400170 -860 400226
rect -804 400170 -736 400226
rect -680 400170 -612 400226
rect -556 400170 -488 400226
rect -432 400170 5514 400226
rect 5570 400170 5638 400226
rect 5694 400170 5762 400226
rect 5818 400170 5886 400226
rect 5942 400170 36234 400226
rect 36290 400170 36358 400226
rect 36414 400170 36482 400226
rect 36538 400170 36606 400226
rect 36662 400170 66954 400226
rect 67010 400170 67078 400226
rect 67134 400170 67202 400226
rect 67258 400170 67326 400226
rect 67382 400170 97674 400226
rect 97730 400170 97798 400226
rect 97854 400170 97922 400226
rect 97978 400170 98046 400226
rect 98102 400170 128394 400226
rect 128450 400170 128518 400226
rect 128574 400170 128642 400226
rect 128698 400170 128766 400226
rect 128822 400170 159114 400226
rect 159170 400170 159238 400226
rect 159294 400170 159362 400226
rect 159418 400170 159486 400226
rect 159542 400170 189834 400226
rect 189890 400170 189958 400226
rect 190014 400170 190082 400226
rect 190138 400170 190206 400226
rect 190262 400170 220554 400226
rect 220610 400170 220678 400226
rect 220734 400170 220802 400226
rect 220858 400170 220926 400226
rect 220982 400170 251274 400226
rect 251330 400170 251398 400226
rect 251454 400170 251522 400226
rect 251578 400170 251646 400226
rect 251702 400170 281994 400226
rect 282050 400170 282118 400226
rect 282174 400170 282242 400226
rect 282298 400170 282366 400226
rect 282422 400170 312714 400226
rect 312770 400170 312838 400226
rect 312894 400170 312962 400226
rect 313018 400170 313086 400226
rect 313142 400170 343434 400226
rect 343490 400170 343558 400226
rect 343614 400170 343682 400226
rect 343738 400170 343806 400226
rect 343862 400170 374154 400226
rect 374210 400170 374278 400226
rect 374334 400170 374402 400226
rect 374458 400170 374526 400226
rect 374582 400170 404874 400226
rect 404930 400170 404998 400226
rect 405054 400170 405122 400226
rect 405178 400170 405246 400226
rect 405302 400170 435594 400226
rect 435650 400170 435718 400226
rect 435774 400170 435842 400226
rect 435898 400170 435966 400226
rect 436022 400170 466314 400226
rect 466370 400170 466438 400226
rect 466494 400170 466562 400226
rect 466618 400170 466686 400226
rect 466742 400170 497034 400226
rect 497090 400170 497158 400226
rect 497214 400170 497282 400226
rect 497338 400170 497406 400226
rect 497462 400170 527754 400226
rect 527810 400170 527878 400226
rect 527934 400170 528002 400226
rect 528058 400170 528126 400226
rect 528182 400170 558474 400226
rect 558530 400170 558598 400226
rect 558654 400170 558722 400226
rect 558778 400170 558846 400226
rect 558902 400170 589194 400226
rect 589250 400170 589318 400226
rect 589374 400170 589442 400226
rect 589498 400170 589566 400226
rect 589622 400170 596496 400226
rect 596552 400170 596620 400226
rect 596676 400170 596744 400226
rect 596800 400170 596868 400226
rect 596924 400170 597980 400226
rect -1916 400102 597980 400170
rect -1916 400046 -860 400102
rect -804 400046 -736 400102
rect -680 400046 -612 400102
rect -556 400046 -488 400102
rect -432 400046 5514 400102
rect 5570 400046 5638 400102
rect 5694 400046 5762 400102
rect 5818 400046 5886 400102
rect 5942 400046 36234 400102
rect 36290 400046 36358 400102
rect 36414 400046 36482 400102
rect 36538 400046 36606 400102
rect 36662 400046 66954 400102
rect 67010 400046 67078 400102
rect 67134 400046 67202 400102
rect 67258 400046 67326 400102
rect 67382 400046 97674 400102
rect 97730 400046 97798 400102
rect 97854 400046 97922 400102
rect 97978 400046 98046 400102
rect 98102 400046 128394 400102
rect 128450 400046 128518 400102
rect 128574 400046 128642 400102
rect 128698 400046 128766 400102
rect 128822 400046 159114 400102
rect 159170 400046 159238 400102
rect 159294 400046 159362 400102
rect 159418 400046 159486 400102
rect 159542 400046 189834 400102
rect 189890 400046 189958 400102
rect 190014 400046 190082 400102
rect 190138 400046 190206 400102
rect 190262 400046 220554 400102
rect 220610 400046 220678 400102
rect 220734 400046 220802 400102
rect 220858 400046 220926 400102
rect 220982 400046 251274 400102
rect 251330 400046 251398 400102
rect 251454 400046 251522 400102
rect 251578 400046 251646 400102
rect 251702 400046 281994 400102
rect 282050 400046 282118 400102
rect 282174 400046 282242 400102
rect 282298 400046 282366 400102
rect 282422 400046 312714 400102
rect 312770 400046 312838 400102
rect 312894 400046 312962 400102
rect 313018 400046 313086 400102
rect 313142 400046 343434 400102
rect 343490 400046 343558 400102
rect 343614 400046 343682 400102
rect 343738 400046 343806 400102
rect 343862 400046 374154 400102
rect 374210 400046 374278 400102
rect 374334 400046 374402 400102
rect 374458 400046 374526 400102
rect 374582 400046 404874 400102
rect 404930 400046 404998 400102
rect 405054 400046 405122 400102
rect 405178 400046 405246 400102
rect 405302 400046 435594 400102
rect 435650 400046 435718 400102
rect 435774 400046 435842 400102
rect 435898 400046 435966 400102
rect 436022 400046 466314 400102
rect 466370 400046 466438 400102
rect 466494 400046 466562 400102
rect 466618 400046 466686 400102
rect 466742 400046 497034 400102
rect 497090 400046 497158 400102
rect 497214 400046 497282 400102
rect 497338 400046 497406 400102
rect 497462 400046 527754 400102
rect 527810 400046 527878 400102
rect 527934 400046 528002 400102
rect 528058 400046 528126 400102
rect 528182 400046 558474 400102
rect 558530 400046 558598 400102
rect 558654 400046 558722 400102
rect 558778 400046 558846 400102
rect 558902 400046 589194 400102
rect 589250 400046 589318 400102
rect 589374 400046 589442 400102
rect 589498 400046 589566 400102
rect 589622 400046 596496 400102
rect 596552 400046 596620 400102
rect 596676 400046 596744 400102
rect 596800 400046 596868 400102
rect 596924 400046 597980 400102
rect -1916 399978 597980 400046
rect -1916 399922 -860 399978
rect -804 399922 -736 399978
rect -680 399922 -612 399978
rect -556 399922 -488 399978
rect -432 399922 5514 399978
rect 5570 399922 5638 399978
rect 5694 399922 5762 399978
rect 5818 399922 5886 399978
rect 5942 399922 36234 399978
rect 36290 399922 36358 399978
rect 36414 399922 36482 399978
rect 36538 399922 36606 399978
rect 36662 399922 66954 399978
rect 67010 399922 67078 399978
rect 67134 399922 67202 399978
rect 67258 399922 67326 399978
rect 67382 399922 97674 399978
rect 97730 399922 97798 399978
rect 97854 399922 97922 399978
rect 97978 399922 98046 399978
rect 98102 399922 128394 399978
rect 128450 399922 128518 399978
rect 128574 399922 128642 399978
rect 128698 399922 128766 399978
rect 128822 399922 159114 399978
rect 159170 399922 159238 399978
rect 159294 399922 159362 399978
rect 159418 399922 159486 399978
rect 159542 399922 189834 399978
rect 189890 399922 189958 399978
rect 190014 399922 190082 399978
rect 190138 399922 190206 399978
rect 190262 399922 220554 399978
rect 220610 399922 220678 399978
rect 220734 399922 220802 399978
rect 220858 399922 220926 399978
rect 220982 399922 251274 399978
rect 251330 399922 251398 399978
rect 251454 399922 251522 399978
rect 251578 399922 251646 399978
rect 251702 399922 281994 399978
rect 282050 399922 282118 399978
rect 282174 399922 282242 399978
rect 282298 399922 282366 399978
rect 282422 399922 312714 399978
rect 312770 399922 312838 399978
rect 312894 399922 312962 399978
rect 313018 399922 313086 399978
rect 313142 399922 343434 399978
rect 343490 399922 343558 399978
rect 343614 399922 343682 399978
rect 343738 399922 343806 399978
rect 343862 399922 374154 399978
rect 374210 399922 374278 399978
rect 374334 399922 374402 399978
rect 374458 399922 374526 399978
rect 374582 399922 404874 399978
rect 404930 399922 404998 399978
rect 405054 399922 405122 399978
rect 405178 399922 405246 399978
rect 405302 399922 435594 399978
rect 435650 399922 435718 399978
rect 435774 399922 435842 399978
rect 435898 399922 435966 399978
rect 436022 399922 466314 399978
rect 466370 399922 466438 399978
rect 466494 399922 466562 399978
rect 466618 399922 466686 399978
rect 466742 399922 497034 399978
rect 497090 399922 497158 399978
rect 497214 399922 497282 399978
rect 497338 399922 497406 399978
rect 497462 399922 527754 399978
rect 527810 399922 527878 399978
rect 527934 399922 528002 399978
rect 528058 399922 528126 399978
rect 528182 399922 558474 399978
rect 558530 399922 558598 399978
rect 558654 399922 558722 399978
rect 558778 399922 558846 399978
rect 558902 399922 589194 399978
rect 589250 399922 589318 399978
rect 589374 399922 589442 399978
rect 589498 399922 589566 399978
rect 589622 399922 596496 399978
rect 596552 399922 596620 399978
rect 596676 399922 596744 399978
rect 596800 399922 596868 399978
rect 596924 399922 597980 399978
rect -1916 399826 597980 399922
rect -1916 388350 597980 388446
rect -1916 388294 -1820 388350
rect -1764 388294 -1696 388350
rect -1640 388294 -1572 388350
rect -1516 388294 -1448 388350
rect -1392 388294 9234 388350
rect 9290 388294 9358 388350
rect 9414 388294 9482 388350
rect 9538 388294 9606 388350
rect 9662 388294 39954 388350
rect 40010 388294 40078 388350
rect 40134 388294 40202 388350
rect 40258 388294 40326 388350
rect 40382 388294 70674 388350
rect 70730 388294 70798 388350
rect 70854 388294 70922 388350
rect 70978 388294 71046 388350
rect 71102 388294 101394 388350
rect 101450 388294 101518 388350
rect 101574 388294 101642 388350
rect 101698 388294 101766 388350
rect 101822 388294 132114 388350
rect 132170 388294 132238 388350
rect 132294 388294 132362 388350
rect 132418 388294 132486 388350
rect 132542 388294 162834 388350
rect 162890 388294 162958 388350
rect 163014 388294 163082 388350
rect 163138 388294 163206 388350
rect 163262 388294 193554 388350
rect 193610 388294 193678 388350
rect 193734 388294 193802 388350
rect 193858 388294 193926 388350
rect 193982 388294 224274 388350
rect 224330 388294 224398 388350
rect 224454 388294 224522 388350
rect 224578 388294 224646 388350
rect 224702 388294 254994 388350
rect 255050 388294 255118 388350
rect 255174 388294 255242 388350
rect 255298 388294 255366 388350
rect 255422 388294 285714 388350
rect 285770 388294 285838 388350
rect 285894 388294 285962 388350
rect 286018 388294 286086 388350
rect 286142 388294 316434 388350
rect 316490 388294 316558 388350
rect 316614 388294 316682 388350
rect 316738 388294 316806 388350
rect 316862 388294 347154 388350
rect 347210 388294 347278 388350
rect 347334 388294 347402 388350
rect 347458 388294 347526 388350
rect 347582 388294 377874 388350
rect 377930 388294 377998 388350
rect 378054 388294 378122 388350
rect 378178 388294 378246 388350
rect 378302 388294 408594 388350
rect 408650 388294 408718 388350
rect 408774 388294 408842 388350
rect 408898 388294 408966 388350
rect 409022 388294 439314 388350
rect 439370 388294 439438 388350
rect 439494 388294 439562 388350
rect 439618 388294 439686 388350
rect 439742 388294 470034 388350
rect 470090 388294 470158 388350
rect 470214 388294 470282 388350
rect 470338 388294 470406 388350
rect 470462 388294 500754 388350
rect 500810 388294 500878 388350
rect 500934 388294 501002 388350
rect 501058 388294 501126 388350
rect 501182 388294 531474 388350
rect 531530 388294 531598 388350
rect 531654 388294 531722 388350
rect 531778 388294 531846 388350
rect 531902 388294 562194 388350
rect 562250 388294 562318 388350
rect 562374 388294 562442 388350
rect 562498 388294 562566 388350
rect 562622 388294 592914 388350
rect 592970 388294 593038 388350
rect 593094 388294 593162 388350
rect 593218 388294 593286 388350
rect 593342 388294 597456 388350
rect 597512 388294 597580 388350
rect 597636 388294 597704 388350
rect 597760 388294 597828 388350
rect 597884 388294 597980 388350
rect -1916 388226 597980 388294
rect -1916 388170 -1820 388226
rect -1764 388170 -1696 388226
rect -1640 388170 -1572 388226
rect -1516 388170 -1448 388226
rect -1392 388170 9234 388226
rect 9290 388170 9358 388226
rect 9414 388170 9482 388226
rect 9538 388170 9606 388226
rect 9662 388170 39954 388226
rect 40010 388170 40078 388226
rect 40134 388170 40202 388226
rect 40258 388170 40326 388226
rect 40382 388170 70674 388226
rect 70730 388170 70798 388226
rect 70854 388170 70922 388226
rect 70978 388170 71046 388226
rect 71102 388170 101394 388226
rect 101450 388170 101518 388226
rect 101574 388170 101642 388226
rect 101698 388170 101766 388226
rect 101822 388170 132114 388226
rect 132170 388170 132238 388226
rect 132294 388170 132362 388226
rect 132418 388170 132486 388226
rect 132542 388170 162834 388226
rect 162890 388170 162958 388226
rect 163014 388170 163082 388226
rect 163138 388170 163206 388226
rect 163262 388170 193554 388226
rect 193610 388170 193678 388226
rect 193734 388170 193802 388226
rect 193858 388170 193926 388226
rect 193982 388170 224274 388226
rect 224330 388170 224398 388226
rect 224454 388170 224522 388226
rect 224578 388170 224646 388226
rect 224702 388170 254994 388226
rect 255050 388170 255118 388226
rect 255174 388170 255242 388226
rect 255298 388170 255366 388226
rect 255422 388170 285714 388226
rect 285770 388170 285838 388226
rect 285894 388170 285962 388226
rect 286018 388170 286086 388226
rect 286142 388170 316434 388226
rect 316490 388170 316558 388226
rect 316614 388170 316682 388226
rect 316738 388170 316806 388226
rect 316862 388170 347154 388226
rect 347210 388170 347278 388226
rect 347334 388170 347402 388226
rect 347458 388170 347526 388226
rect 347582 388170 377874 388226
rect 377930 388170 377998 388226
rect 378054 388170 378122 388226
rect 378178 388170 378246 388226
rect 378302 388170 408594 388226
rect 408650 388170 408718 388226
rect 408774 388170 408842 388226
rect 408898 388170 408966 388226
rect 409022 388170 439314 388226
rect 439370 388170 439438 388226
rect 439494 388170 439562 388226
rect 439618 388170 439686 388226
rect 439742 388170 470034 388226
rect 470090 388170 470158 388226
rect 470214 388170 470282 388226
rect 470338 388170 470406 388226
rect 470462 388170 500754 388226
rect 500810 388170 500878 388226
rect 500934 388170 501002 388226
rect 501058 388170 501126 388226
rect 501182 388170 531474 388226
rect 531530 388170 531598 388226
rect 531654 388170 531722 388226
rect 531778 388170 531846 388226
rect 531902 388170 562194 388226
rect 562250 388170 562318 388226
rect 562374 388170 562442 388226
rect 562498 388170 562566 388226
rect 562622 388170 592914 388226
rect 592970 388170 593038 388226
rect 593094 388170 593162 388226
rect 593218 388170 593286 388226
rect 593342 388170 597456 388226
rect 597512 388170 597580 388226
rect 597636 388170 597704 388226
rect 597760 388170 597828 388226
rect 597884 388170 597980 388226
rect -1916 388102 597980 388170
rect -1916 388046 -1820 388102
rect -1764 388046 -1696 388102
rect -1640 388046 -1572 388102
rect -1516 388046 -1448 388102
rect -1392 388046 9234 388102
rect 9290 388046 9358 388102
rect 9414 388046 9482 388102
rect 9538 388046 9606 388102
rect 9662 388046 39954 388102
rect 40010 388046 40078 388102
rect 40134 388046 40202 388102
rect 40258 388046 40326 388102
rect 40382 388046 70674 388102
rect 70730 388046 70798 388102
rect 70854 388046 70922 388102
rect 70978 388046 71046 388102
rect 71102 388046 101394 388102
rect 101450 388046 101518 388102
rect 101574 388046 101642 388102
rect 101698 388046 101766 388102
rect 101822 388046 132114 388102
rect 132170 388046 132238 388102
rect 132294 388046 132362 388102
rect 132418 388046 132486 388102
rect 132542 388046 162834 388102
rect 162890 388046 162958 388102
rect 163014 388046 163082 388102
rect 163138 388046 163206 388102
rect 163262 388046 193554 388102
rect 193610 388046 193678 388102
rect 193734 388046 193802 388102
rect 193858 388046 193926 388102
rect 193982 388046 224274 388102
rect 224330 388046 224398 388102
rect 224454 388046 224522 388102
rect 224578 388046 224646 388102
rect 224702 388046 254994 388102
rect 255050 388046 255118 388102
rect 255174 388046 255242 388102
rect 255298 388046 255366 388102
rect 255422 388046 285714 388102
rect 285770 388046 285838 388102
rect 285894 388046 285962 388102
rect 286018 388046 286086 388102
rect 286142 388046 316434 388102
rect 316490 388046 316558 388102
rect 316614 388046 316682 388102
rect 316738 388046 316806 388102
rect 316862 388046 347154 388102
rect 347210 388046 347278 388102
rect 347334 388046 347402 388102
rect 347458 388046 347526 388102
rect 347582 388046 377874 388102
rect 377930 388046 377998 388102
rect 378054 388046 378122 388102
rect 378178 388046 378246 388102
rect 378302 388046 408594 388102
rect 408650 388046 408718 388102
rect 408774 388046 408842 388102
rect 408898 388046 408966 388102
rect 409022 388046 439314 388102
rect 439370 388046 439438 388102
rect 439494 388046 439562 388102
rect 439618 388046 439686 388102
rect 439742 388046 470034 388102
rect 470090 388046 470158 388102
rect 470214 388046 470282 388102
rect 470338 388046 470406 388102
rect 470462 388046 500754 388102
rect 500810 388046 500878 388102
rect 500934 388046 501002 388102
rect 501058 388046 501126 388102
rect 501182 388046 531474 388102
rect 531530 388046 531598 388102
rect 531654 388046 531722 388102
rect 531778 388046 531846 388102
rect 531902 388046 562194 388102
rect 562250 388046 562318 388102
rect 562374 388046 562442 388102
rect 562498 388046 562566 388102
rect 562622 388046 592914 388102
rect 592970 388046 593038 388102
rect 593094 388046 593162 388102
rect 593218 388046 593286 388102
rect 593342 388046 597456 388102
rect 597512 388046 597580 388102
rect 597636 388046 597704 388102
rect 597760 388046 597828 388102
rect 597884 388046 597980 388102
rect -1916 387978 597980 388046
rect -1916 387922 -1820 387978
rect -1764 387922 -1696 387978
rect -1640 387922 -1572 387978
rect -1516 387922 -1448 387978
rect -1392 387922 9234 387978
rect 9290 387922 9358 387978
rect 9414 387922 9482 387978
rect 9538 387922 9606 387978
rect 9662 387922 39954 387978
rect 40010 387922 40078 387978
rect 40134 387922 40202 387978
rect 40258 387922 40326 387978
rect 40382 387922 70674 387978
rect 70730 387922 70798 387978
rect 70854 387922 70922 387978
rect 70978 387922 71046 387978
rect 71102 387922 101394 387978
rect 101450 387922 101518 387978
rect 101574 387922 101642 387978
rect 101698 387922 101766 387978
rect 101822 387922 132114 387978
rect 132170 387922 132238 387978
rect 132294 387922 132362 387978
rect 132418 387922 132486 387978
rect 132542 387922 162834 387978
rect 162890 387922 162958 387978
rect 163014 387922 163082 387978
rect 163138 387922 163206 387978
rect 163262 387922 193554 387978
rect 193610 387922 193678 387978
rect 193734 387922 193802 387978
rect 193858 387922 193926 387978
rect 193982 387922 224274 387978
rect 224330 387922 224398 387978
rect 224454 387922 224522 387978
rect 224578 387922 224646 387978
rect 224702 387922 254994 387978
rect 255050 387922 255118 387978
rect 255174 387922 255242 387978
rect 255298 387922 255366 387978
rect 255422 387922 285714 387978
rect 285770 387922 285838 387978
rect 285894 387922 285962 387978
rect 286018 387922 286086 387978
rect 286142 387922 316434 387978
rect 316490 387922 316558 387978
rect 316614 387922 316682 387978
rect 316738 387922 316806 387978
rect 316862 387922 347154 387978
rect 347210 387922 347278 387978
rect 347334 387922 347402 387978
rect 347458 387922 347526 387978
rect 347582 387922 377874 387978
rect 377930 387922 377998 387978
rect 378054 387922 378122 387978
rect 378178 387922 378246 387978
rect 378302 387922 408594 387978
rect 408650 387922 408718 387978
rect 408774 387922 408842 387978
rect 408898 387922 408966 387978
rect 409022 387922 439314 387978
rect 439370 387922 439438 387978
rect 439494 387922 439562 387978
rect 439618 387922 439686 387978
rect 439742 387922 470034 387978
rect 470090 387922 470158 387978
rect 470214 387922 470282 387978
rect 470338 387922 470406 387978
rect 470462 387922 500754 387978
rect 500810 387922 500878 387978
rect 500934 387922 501002 387978
rect 501058 387922 501126 387978
rect 501182 387922 531474 387978
rect 531530 387922 531598 387978
rect 531654 387922 531722 387978
rect 531778 387922 531846 387978
rect 531902 387922 562194 387978
rect 562250 387922 562318 387978
rect 562374 387922 562442 387978
rect 562498 387922 562566 387978
rect 562622 387922 592914 387978
rect 592970 387922 593038 387978
rect 593094 387922 593162 387978
rect 593218 387922 593286 387978
rect 593342 387922 597456 387978
rect 597512 387922 597580 387978
rect 597636 387922 597704 387978
rect 597760 387922 597828 387978
rect 597884 387922 597980 387978
rect -1916 387826 597980 387922
rect -1916 382350 597980 382446
rect -1916 382294 -860 382350
rect -804 382294 -736 382350
rect -680 382294 -612 382350
rect -556 382294 -488 382350
rect -432 382294 5514 382350
rect 5570 382294 5638 382350
rect 5694 382294 5762 382350
rect 5818 382294 5886 382350
rect 5942 382294 36234 382350
rect 36290 382294 36358 382350
rect 36414 382294 36482 382350
rect 36538 382294 36606 382350
rect 36662 382294 66954 382350
rect 67010 382294 67078 382350
rect 67134 382294 67202 382350
rect 67258 382294 67326 382350
rect 67382 382294 97674 382350
rect 97730 382294 97798 382350
rect 97854 382294 97922 382350
rect 97978 382294 98046 382350
rect 98102 382294 128394 382350
rect 128450 382294 128518 382350
rect 128574 382294 128642 382350
rect 128698 382294 128766 382350
rect 128822 382294 159114 382350
rect 159170 382294 159238 382350
rect 159294 382294 159362 382350
rect 159418 382294 159486 382350
rect 159542 382294 189834 382350
rect 189890 382294 189958 382350
rect 190014 382294 190082 382350
rect 190138 382294 190206 382350
rect 190262 382294 220554 382350
rect 220610 382294 220678 382350
rect 220734 382294 220802 382350
rect 220858 382294 220926 382350
rect 220982 382294 251274 382350
rect 251330 382294 251398 382350
rect 251454 382294 251522 382350
rect 251578 382294 251646 382350
rect 251702 382294 281994 382350
rect 282050 382294 282118 382350
rect 282174 382294 282242 382350
rect 282298 382294 282366 382350
rect 282422 382294 312714 382350
rect 312770 382294 312838 382350
rect 312894 382294 312962 382350
rect 313018 382294 313086 382350
rect 313142 382294 343434 382350
rect 343490 382294 343558 382350
rect 343614 382294 343682 382350
rect 343738 382294 343806 382350
rect 343862 382294 374154 382350
rect 374210 382294 374278 382350
rect 374334 382294 374402 382350
rect 374458 382294 374526 382350
rect 374582 382294 404874 382350
rect 404930 382294 404998 382350
rect 405054 382294 405122 382350
rect 405178 382294 405246 382350
rect 405302 382294 435594 382350
rect 435650 382294 435718 382350
rect 435774 382294 435842 382350
rect 435898 382294 435966 382350
rect 436022 382294 466314 382350
rect 466370 382294 466438 382350
rect 466494 382294 466562 382350
rect 466618 382294 466686 382350
rect 466742 382294 497034 382350
rect 497090 382294 497158 382350
rect 497214 382294 497282 382350
rect 497338 382294 497406 382350
rect 497462 382294 527754 382350
rect 527810 382294 527878 382350
rect 527934 382294 528002 382350
rect 528058 382294 528126 382350
rect 528182 382294 558474 382350
rect 558530 382294 558598 382350
rect 558654 382294 558722 382350
rect 558778 382294 558846 382350
rect 558902 382294 589194 382350
rect 589250 382294 589318 382350
rect 589374 382294 589442 382350
rect 589498 382294 589566 382350
rect 589622 382294 596496 382350
rect 596552 382294 596620 382350
rect 596676 382294 596744 382350
rect 596800 382294 596868 382350
rect 596924 382294 597980 382350
rect -1916 382226 597980 382294
rect -1916 382170 -860 382226
rect -804 382170 -736 382226
rect -680 382170 -612 382226
rect -556 382170 -488 382226
rect -432 382170 5514 382226
rect 5570 382170 5638 382226
rect 5694 382170 5762 382226
rect 5818 382170 5886 382226
rect 5942 382170 36234 382226
rect 36290 382170 36358 382226
rect 36414 382170 36482 382226
rect 36538 382170 36606 382226
rect 36662 382170 66954 382226
rect 67010 382170 67078 382226
rect 67134 382170 67202 382226
rect 67258 382170 67326 382226
rect 67382 382170 97674 382226
rect 97730 382170 97798 382226
rect 97854 382170 97922 382226
rect 97978 382170 98046 382226
rect 98102 382170 128394 382226
rect 128450 382170 128518 382226
rect 128574 382170 128642 382226
rect 128698 382170 128766 382226
rect 128822 382170 159114 382226
rect 159170 382170 159238 382226
rect 159294 382170 159362 382226
rect 159418 382170 159486 382226
rect 159542 382170 189834 382226
rect 189890 382170 189958 382226
rect 190014 382170 190082 382226
rect 190138 382170 190206 382226
rect 190262 382170 220554 382226
rect 220610 382170 220678 382226
rect 220734 382170 220802 382226
rect 220858 382170 220926 382226
rect 220982 382170 251274 382226
rect 251330 382170 251398 382226
rect 251454 382170 251522 382226
rect 251578 382170 251646 382226
rect 251702 382170 281994 382226
rect 282050 382170 282118 382226
rect 282174 382170 282242 382226
rect 282298 382170 282366 382226
rect 282422 382170 312714 382226
rect 312770 382170 312838 382226
rect 312894 382170 312962 382226
rect 313018 382170 313086 382226
rect 313142 382170 343434 382226
rect 343490 382170 343558 382226
rect 343614 382170 343682 382226
rect 343738 382170 343806 382226
rect 343862 382170 374154 382226
rect 374210 382170 374278 382226
rect 374334 382170 374402 382226
rect 374458 382170 374526 382226
rect 374582 382170 404874 382226
rect 404930 382170 404998 382226
rect 405054 382170 405122 382226
rect 405178 382170 405246 382226
rect 405302 382170 435594 382226
rect 435650 382170 435718 382226
rect 435774 382170 435842 382226
rect 435898 382170 435966 382226
rect 436022 382170 466314 382226
rect 466370 382170 466438 382226
rect 466494 382170 466562 382226
rect 466618 382170 466686 382226
rect 466742 382170 497034 382226
rect 497090 382170 497158 382226
rect 497214 382170 497282 382226
rect 497338 382170 497406 382226
rect 497462 382170 527754 382226
rect 527810 382170 527878 382226
rect 527934 382170 528002 382226
rect 528058 382170 528126 382226
rect 528182 382170 558474 382226
rect 558530 382170 558598 382226
rect 558654 382170 558722 382226
rect 558778 382170 558846 382226
rect 558902 382170 589194 382226
rect 589250 382170 589318 382226
rect 589374 382170 589442 382226
rect 589498 382170 589566 382226
rect 589622 382170 596496 382226
rect 596552 382170 596620 382226
rect 596676 382170 596744 382226
rect 596800 382170 596868 382226
rect 596924 382170 597980 382226
rect -1916 382102 597980 382170
rect -1916 382046 -860 382102
rect -804 382046 -736 382102
rect -680 382046 -612 382102
rect -556 382046 -488 382102
rect -432 382046 5514 382102
rect 5570 382046 5638 382102
rect 5694 382046 5762 382102
rect 5818 382046 5886 382102
rect 5942 382046 36234 382102
rect 36290 382046 36358 382102
rect 36414 382046 36482 382102
rect 36538 382046 36606 382102
rect 36662 382046 66954 382102
rect 67010 382046 67078 382102
rect 67134 382046 67202 382102
rect 67258 382046 67326 382102
rect 67382 382046 97674 382102
rect 97730 382046 97798 382102
rect 97854 382046 97922 382102
rect 97978 382046 98046 382102
rect 98102 382046 128394 382102
rect 128450 382046 128518 382102
rect 128574 382046 128642 382102
rect 128698 382046 128766 382102
rect 128822 382046 159114 382102
rect 159170 382046 159238 382102
rect 159294 382046 159362 382102
rect 159418 382046 159486 382102
rect 159542 382046 189834 382102
rect 189890 382046 189958 382102
rect 190014 382046 190082 382102
rect 190138 382046 190206 382102
rect 190262 382046 220554 382102
rect 220610 382046 220678 382102
rect 220734 382046 220802 382102
rect 220858 382046 220926 382102
rect 220982 382046 251274 382102
rect 251330 382046 251398 382102
rect 251454 382046 251522 382102
rect 251578 382046 251646 382102
rect 251702 382046 281994 382102
rect 282050 382046 282118 382102
rect 282174 382046 282242 382102
rect 282298 382046 282366 382102
rect 282422 382046 312714 382102
rect 312770 382046 312838 382102
rect 312894 382046 312962 382102
rect 313018 382046 313086 382102
rect 313142 382046 343434 382102
rect 343490 382046 343558 382102
rect 343614 382046 343682 382102
rect 343738 382046 343806 382102
rect 343862 382046 374154 382102
rect 374210 382046 374278 382102
rect 374334 382046 374402 382102
rect 374458 382046 374526 382102
rect 374582 382046 404874 382102
rect 404930 382046 404998 382102
rect 405054 382046 405122 382102
rect 405178 382046 405246 382102
rect 405302 382046 435594 382102
rect 435650 382046 435718 382102
rect 435774 382046 435842 382102
rect 435898 382046 435966 382102
rect 436022 382046 466314 382102
rect 466370 382046 466438 382102
rect 466494 382046 466562 382102
rect 466618 382046 466686 382102
rect 466742 382046 497034 382102
rect 497090 382046 497158 382102
rect 497214 382046 497282 382102
rect 497338 382046 497406 382102
rect 497462 382046 527754 382102
rect 527810 382046 527878 382102
rect 527934 382046 528002 382102
rect 528058 382046 528126 382102
rect 528182 382046 558474 382102
rect 558530 382046 558598 382102
rect 558654 382046 558722 382102
rect 558778 382046 558846 382102
rect 558902 382046 589194 382102
rect 589250 382046 589318 382102
rect 589374 382046 589442 382102
rect 589498 382046 589566 382102
rect 589622 382046 596496 382102
rect 596552 382046 596620 382102
rect 596676 382046 596744 382102
rect 596800 382046 596868 382102
rect 596924 382046 597980 382102
rect -1916 381978 597980 382046
rect -1916 381922 -860 381978
rect -804 381922 -736 381978
rect -680 381922 -612 381978
rect -556 381922 -488 381978
rect -432 381922 5514 381978
rect 5570 381922 5638 381978
rect 5694 381922 5762 381978
rect 5818 381922 5886 381978
rect 5942 381922 36234 381978
rect 36290 381922 36358 381978
rect 36414 381922 36482 381978
rect 36538 381922 36606 381978
rect 36662 381922 66954 381978
rect 67010 381922 67078 381978
rect 67134 381922 67202 381978
rect 67258 381922 67326 381978
rect 67382 381922 97674 381978
rect 97730 381922 97798 381978
rect 97854 381922 97922 381978
rect 97978 381922 98046 381978
rect 98102 381922 128394 381978
rect 128450 381922 128518 381978
rect 128574 381922 128642 381978
rect 128698 381922 128766 381978
rect 128822 381922 159114 381978
rect 159170 381922 159238 381978
rect 159294 381922 159362 381978
rect 159418 381922 159486 381978
rect 159542 381922 189834 381978
rect 189890 381922 189958 381978
rect 190014 381922 190082 381978
rect 190138 381922 190206 381978
rect 190262 381922 220554 381978
rect 220610 381922 220678 381978
rect 220734 381922 220802 381978
rect 220858 381922 220926 381978
rect 220982 381922 251274 381978
rect 251330 381922 251398 381978
rect 251454 381922 251522 381978
rect 251578 381922 251646 381978
rect 251702 381922 281994 381978
rect 282050 381922 282118 381978
rect 282174 381922 282242 381978
rect 282298 381922 282366 381978
rect 282422 381922 312714 381978
rect 312770 381922 312838 381978
rect 312894 381922 312962 381978
rect 313018 381922 313086 381978
rect 313142 381922 343434 381978
rect 343490 381922 343558 381978
rect 343614 381922 343682 381978
rect 343738 381922 343806 381978
rect 343862 381922 374154 381978
rect 374210 381922 374278 381978
rect 374334 381922 374402 381978
rect 374458 381922 374526 381978
rect 374582 381922 404874 381978
rect 404930 381922 404998 381978
rect 405054 381922 405122 381978
rect 405178 381922 405246 381978
rect 405302 381922 435594 381978
rect 435650 381922 435718 381978
rect 435774 381922 435842 381978
rect 435898 381922 435966 381978
rect 436022 381922 466314 381978
rect 466370 381922 466438 381978
rect 466494 381922 466562 381978
rect 466618 381922 466686 381978
rect 466742 381922 497034 381978
rect 497090 381922 497158 381978
rect 497214 381922 497282 381978
rect 497338 381922 497406 381978
rect 497462 381922 527754 381978
rect 527810 381922 527878 381978
rect 527934 381922 528002 381978
rect 528058 381922 528126 381978
rect 528182 381922 558474 381978
rect 558530 381922 558598 381978
rect 558654 381922 558722 381978
rect 558778 381922 558846 381978
rect 558902 381922 589194 381978
rect 589250 381922 589318 381978
rect 589374 381922 589442 381978
rect 589498 381922 589566 381978
rect 589622 381922 596496 381978
rect 596552 381922 596620 381978
rect 596676 381922 596744 381978
rect 596800 381922 596868 381978
rect 596924 381922 597980 381978
rect -1916 381826 597980 381922
rect -1916 370350 597980 370446
rect -1916 370294 -1820 370350
rect -1764 370294 -1696 370350
rect -1640 370294 -1572 370350
rect -1516 370294 -1448 370350
rect -1392 370294 9234 370350
rect 9290 370294 9358 370350
rect 9414 370294 9482 370350
rect 9538 370294 9606 370350
rect 9662 370294 39954 370350
rect 40010 370294 40078 370350
rect 40134 370294 40202 370350
rect 40258 370294 40326 370350
rect 40382 370294 70674 370350
rect 70730 370294 70798 370350
rect 70854 370294 70922 370350
rect 70978 370294 71046 370350
rect 71102 370294 101394 370350
rect 101450 370294 101518 370350
rect 101574 370294 101642 370350
rect 101698 370294 101766 370350
rect 101822 370294 132114 370350
rect 132170 370294 132238 370350
rect 132294 370294 132362 370350
rect 132418 370294 132486 370350
rect 132542 370294 162834 370350
rect 162890 370294 162958 370350
rect 163014 370294 163082 370350
rect 163138 370294 163206 370350
rect 163262 370294 193554 370350
rect 193610 370294 193678 370350
rect 193734 370294 193802 370350
rect 193858 370294 193926 370350
rect 193982 370294 224274 370350
rect 224330 370294 224398 370350
rect 224454 370294 224522 370350
rect 224578 370294 224646 370350
rect 224702 370294 254994 370350
rect 255050 370294 255118 370350
rect 255174 370294 255242 370350
rect 255298 370294 255366 370350
rect 255422 370294 285714 370350
rect 285770 370294 285838 370350
rect 285894 370294 285962 370350
rect 286018 370294 286086 370350
rect 286142 370294 316434 370350
rect 316490 370294 316558 370350
rect 316614 370294 316682 370350
rect 316738 370294 316806 370350
rect 316862 370294 347154 370350
rect 347210 370294 347278 370350
rect 347334 370294 347402 370350
rect 347458 370294 347526 370350
rect 347582 370294 377874 370350
rect 377930 370294 377998 370350
rect 378054 370294 378122 370350
rect 378178 370294 378246 370350
rect 378302 370294 408594 370350
rect 408650 370294 408718 370350
rect 408774 370294 408842 370350
rect 408898 370294 408966 370350
rect 409022 370294 439314 370350
rect 439370 370294 439438 370350
rect 439494 370294 439562 370350
rect 439618 370294 439686 370350
rect 439742 370294 470034 370350
rect 470090 370294 470158 370350
rect 470214 370294 470282 370350
rect 470338 370294 470406 370350
rect 470462 370294 500754 370350
rect 500810 370294 500878 370350
rect 500934 370294 501002 370350
rect 501058 370294 501126 370350
rect 501182 370294 531474 370350
rect 531530 370294 531598 370350
rect 531654 370294 531722 370350
rect 531778 370294 531846 370350
rect 531902 370294 562194 370350
rect 562250 370294 562318 370350
rect 562374 370294 562442 370350
rect 562498 370294 562566 370350
rect 562622 370294 592914 370350
rect 592970 370294 593038 370350
rect 593094 370294 593162 370350
rect 593218 370294 593286 370350
rect 593342 370294 597456 370350
rect 597512 370294 597580 370350
rect 597636 370294 597704 370350
rect 597760 370294 597828 370350
rect 597884 370294 597980 370350
rect -1916 370226 597980 370294
rect -1916 370170 -1820 370226
rect -1764 370170 -1696 370226
rect -1640 370170 -1572 370226
rect -1516 370170 -1448 370226
rect -1392 370170 9234 370226
rect 9290 370170 9358 370226
rect 9414 370170 9482 370226
rect 9538 370170 9606 370226
rect 9662 370170 39954 370226
rect 40010 370170 40078 370226
rect 40134 370170 40202 370226
rect 40258 370170 40326 370226
rect 40382 370170 70674 370226
rect 70730 370170 70798 370226
rect 70854 370170 70922 370226
rect 70978 370170 71046 370226
rect 71102 370170 101394 370226
rect 101450 370170 101518 370226
rect 101574 370170 101642 370226
rect 101698 370170 101766 370226
rect 101822 370170 132114 370226
rect 132170 370170 132238 370226
rect 132294 370170 132362 370226
rect 132418 370170 132486 370226
rect 132542 370170 162834 370226
rect 162890 370170 162958 370226
rect 163014 370170 163082 370226
rect 163138 370170 163206 370226
rect 163262 370170 193554 370226
rect 193610 370170 193678 370226
rect 193734 370170 193802 370226
rect 193858 370170 193926 370226
rect 193982 370170 224274 370226
rect 224330 370170 224398 370226
rect 224454 370170 224522 370226
rect 224578 370170 224646 370226
rect 224702 370170 254994 370226
rect 255050 370170 255118 370226
rect 255174 370170 255242 370226
rect 255298 370170 255366 370226
rect 255422 370170 285714 370226
rect 285770 370170 285838 370226
rect 285894 370170 285962 370226
rect 286018 370170 286086 370226
rect 286142 370170 316434 370226
rect 316490 370170 316558 370226
rect 316614 370170 316682 370226
rect 316738 370170 316806 370226
rect 316862 370170 347154 370226
rect 347210 370170 347278 370226
rect 347334 370170 347402 370226
rect 347458 370170 347526 370226
rect 347582 370170 377874 370226
rect 377930 370170 377998 370226
rect 378054 370170 378122 370226
rect 378178 370170 378246 370226
rect 378302 370170 408594 370226
rect 408650 370170 408718 370226
rect 408774 370170 408842 370226
rect 408898 370170 408966 370226
rect 409022 370170 439314 370226
rect 439370 370170 439438 370226
rect 439494 370170 439562 370226
rect 439618 370170 439686 370226
rect 439742 370170 470034 370226
rect 470090 370170 470158 370226
rect 470214 370170 470282 370226
rect 470338 370170 470406 370226
rect 470462 370170 500754 370226
rect 500810 370170 500878 370226
rect 500934 370170 501002 370226
rect 501058 370170 501126 370226
rect 501182 370170 531474 370226
rect 531530 370170 531598 370226
rect 531654 370170 531722 370226
rect 531778 370170 531846 370226
rect 531902 370170 562194 370226
rect 562250 370170 562318 370226
rect 562374 370170 562442 370226
rect 562498 370170 562566 370226
rect 562622 370170 592914 370226
rect 592970 370170 593038 370226
rect 593094 370170 593162 370226
rect 593218 370170 593286 370226
rect 593342 370170 597456 370226
rect 597512 370170 597580 370226
rect 597636 370170 597704 370226
rect 597760 370170 597828 370226
rect 597884 370170 597980 370226
rect -1916 370102 597980 370170
rect -1916 370046 -1820 370102
rect -1764 370046 -1696 370102
rect -1640 370046 -1572 370102
rect -1516 370046 -1448 370102
rect -1392 370046 9234 370102
rect 9290 370046 9358 370102
rect 9414 370046 9482 370102
rect 9538 370046 9606 370102
rect 9662 370046 39954 370102
rect 40010 370046 40078 370102
rect 40134 370046 40202 370102
rect 40258 370046 40326 370102
rect 40382 370046 70674 370102
rect 70730 370046 70798 370102
rect 70854 370046 70922 370102
rect 70978 370046 71046 370102
rect 71102 370046 101394 370102
rect 101450 370046 101518 370102
rect 101574 370046 101642 370102
rect 101698 370046 101766 370102
rect 101822 370046 132114 370102
rect 132170 370046 132238 370102
rect 132294 370046 132362 370102
rect 132418 370046 132486 370102
rect 132542 370046 162834 370102
rect 162890 370046 162958 370102
rect 163014 370046 163082 370102
rect 163138 370046 163206 370102
rect 163262 370046 193554 370102
rect 193610 370046 193678 370102
rect 193734 370046 193802 370102
rect 193858 370046 193926 370102
rect 193982 370046 224274 370102
rect 224330 370046 224398 370102
rect 224454 370046 224522 370102
rect 224578 370046 224646 370102
rect 224702 370046 254994 370102
rect 255050 370046 255118 370102
rect 255174 370046 255242 370102
rect 255298 370046 255366 370102
rect 255422 370046 285714 370102
rect 285770 370046 285838 370102
rect 285894 370046 285962 370102
rect 286018 370046 286086 370102
rect 286142 370046 316434 370102
rect 316490 370046 316558 370102
rect 316614 370046 316682 370102
rect 316738 370046 316806 370102
rect 316862 370046 347154 370102
rect 347210 370046 347278 370102
rect 347334 370046 347402 370102
rect 347458 370046 347526 370102
rect 347582 370046 377874 370102
rect 377930 370046 377998 370102
rect 378054 370046 378122 370102
rect 378178 370046 378246 370102
rect 378302 370046 408594 370102
rect 408650 370046 408718 370102
rect 408774 370046 408842 370102
rect 408898 370046 408966 370102
rect 409022 370046 439314 370102
rect 439370 370046 439438 370102
rect 439494 370046 439562 370102
rect 439618 370046 439686 370102
rect 439742 370046 470034 370102
rect 470090 370046 470158 370102
rect 470214 370046 470282 370102
rect 470338 370046 470406 370102
rect 470462 370046 500754 370102
rect 500810 370046 500878 370102
rect 500934 370046 501002 370102
rect 501058 370046 501126 370102
rect 501182 370046 531474 370102
rect 531530 370046 531598 370102
rect 531654 370046 531722 370102
rect 531778 370046 531846 370102
rect 531902 370046 562194 370102
rect 562250 370046 562318 370102
rect 562374 370046 562442 370102
rect 562498 370046 562566 370102
rect 562622 370046 592914 370102
rect 592970 370046 593038 370102
rect 593094 370046 593162 370102
rect 593218 370046 593286 370102
rect 593342 370046 597456 370102
rect 597512 370046 597580 370102
rect 597636 370046 597704 370102
rect 597760 370046 597828 370102
rect 597884 370046 597980 370102
rect -1916 369978 597980 370046
rect -1916 369922 -1820 369978
rect -1764 369922 -1696 369978
rect -1640 369922 -1572 369978
rect -1516 369922 -1448 369978
rect -1392 369922 9234 369978
rect 9290 369922 9358 369978
rect 9414 369922 9482 369978
rect 9538 369922 9606 369978
rect 9662 369922 39954 369978
rect 40010 369922 40078 369978
rect 40134 369922 40202 369978
rect 40258 369922 40326 369978
rect 40382 369922 70674 369978
rect 70730 369922 70798 369978
rect 70854 369922 70922 369978
rect 70978 369922 71046 369978
rect 71102 369922 101394 369978
rect 101450 369922 101518 369978
rect 101574 369922 101642 369978
rect 101698 369922 101766 369978
rect 101822 369922 132114 369978
rect 132170 369922 132238 369978
rect 132294 369922 132362 369978
rect 132418 369922 132486 369978
rect 132542 369922 162834 369978
rect 162890 369922 162958 369978
rect 163014 369922 163082 369978
rect 163138 369922 163206 369978
rect 163262 369922 193554 369978
rect 193610 369922 193678 369978
rect 193734 369922 193802 369978
rect 193858 369922 193926 369978
rect 193982 369922 224274 369978
rect 224330 369922 224398 369978
rect 224454 369922 224522 369978
rect 224578 369922 224646 369978
rect 224702 369922 254994 369978
rect 255050 369922 255118 369978
rect 255174 369922 255242 369978
rect 255298 369922 255366 369978
rect 255422 369922 285714 369978
rect 285770 369922 285838 369978
rect 285894 369922 285962 369978
rect 286018 369922 286086 369978
rect 286142 369922 316434 369978
rect 316490 369922 316558 369978
rect 316614 369922 316682 369978
rect 316738 369922 316806 369978
rect 316862 369922 347154 369978
rect 347210 369922 347278 369978
rect 347334 369922 347402 369978
rect 347458 369922 347526 369978
rect 347582 369922 377874 369978
rect 377930 369922 377998 369978
rect 378054 369922 378122 369978
rect 378178 369922 378246 369978
rect 378302 369922 408594 369978
rect 408650 369922 408718 369978
rect 408774 369922 408842 369978
rect 408898 369922 408966 369978
rect 409022 369922 439314 369978
rect 439370 369922 439438 369978
rect 439494 369922 439562 369978
rect 439618 369922 439686 369978
rect 439742 369922 470034 369978
rect 470090 369922 470158 369978
rect 470214 369922 470282 369978
rect 470338 369922 470406 369978
rect 470462 369922 500754 369978
rect 500810 369922 500878 369978
rect 500934 369922 501002 369978
rect 501058 369922 501126 369978
rect 501182 369922 531474 369978
rect 531530 369922 531598 369978
rect 531654 369922 531722 369978
rect 531778 369922 531846 369978
rect 531902 369922 562194 369978
rect 562250 369922 562318 369978
rect 562374 369922 562442 369978
rect 562498 369922 562566 369978
rect 562622 369922 592914 369978
rect 592970 369922 593038 369978
rect 593094 369922 593162 369978
rect 593218 369922 593286 369978
rect 593342 369922 597456 369978
rect 597512 369922 597580 369978
rect 597636 369922 597704 369978
rect 597760 369922 597828 369978
rect 597884 369922 597980 369978
rect -1916 369826 597980 369922
rect -1916 364350 597980 364446
rect -1916 364294 -860 364350
rect -804 364294 -736 364350
rect -680 364294 -612 364350
rect -556 364294 -488 364350
rect -432 364294 5514 364350
rect 5570 364294 5638 364350
rect 5694 364294 5762 364350
rect 5818 364294 5886 364350
rect 5942 364294 36234 364350
rect 36290 364294 36358 364350
rect 36414 364294 36482 364350
rect 36538 364294 36606 364350
rect 36662 364294 66954 364350
rect 67010 364294 67078 364350
rect 67134 364294 67202 364350
rect 67258 364294 67326 364350
rect 67382 364294 97674 364350
rect 97730 364294 97798 364350
rect 97854 364294 97922 364350
rect 97978 364294 98046 364350
rect 98102 364294 128394 364350
rect 128450 364294 128518 364350
rect 128574 364294 128642 364350
rect 128698 364294 128766 364350
rect 128822 364294 159114 364350
rect 159170 364294 159238 364350
rect 159294 364294 159362 364350
rect 159418 364294 159486 364350
rect 159542 364294 189834 364350
rect 189890 364294 189958 364350
rect 190014 364294 190082 364350
rect 190138 364294 190206 364350
rect 190262 364294 220554 364350
rect 220610 364294 220678 364350
rect 220734 364294 220802 364350
rect 220858 364294 220926 364350
rect 220982 364294 251274 364350
rect 251330 364294 251398 364350
rect 251454 364294 251522 364350
rect 251578 364294 251646 364350
rect 251702 364294 281994 364350
rect 282050 364294 282118 364350
rect 282174 364294 282242 364350
rect 282298 364294 282366 364350
rect 282422 364294 312714 364350
rect 312770 364294 312838 364350
rect 312894 364294 312962 364350
rect 313018 364294 313086 364350
rect 313142 364294 343434 364350
rect 343490 364294 343558 364350
rect 343614 364294 343682 364350
rect 343738 364294 343806 364350
rect 343862 364294 374154 364350
rect 374210 364294 374278 364350
rect 374334 364294 374402 364350
rect 374458 364294 374526 364350
rect 374582 364294 404874 364350
rect 404930 364294 404998 364350
rect 405054 364294 405122 364350
rect 405178 364294 405246 364350
rect 405302 364294 435594 364350
rect 435650 364294 435718 364350
rect 435774 364294 435842 364350
rect 435898 364294 435966 364350
rect 436022 364294 466314 364350
rect 466370 364294 466438 364350
rect 466494 364294 466562 364350
rect 466618 364294 466686 364350
rect 466742 364294 497034 364350
rect 497090 364294 497158 364350
rect 497214 364294 497282 364350
rect 497338 364294 497406 364350
rect 497462 364294 527754 364350
rect 527810 364294 527878 364350
rect 527934 364294 528002 364350
rect 528058 364294 528126 364350
rect 528182 364294 558474 364350
rect 558530 364294 558598 364350
rect 558654 364294 558722 364350
rect 558778 364294 558846 364350
rect 558902 364294 589194 364350
rect 589250 364294 589318 364350
rect 589374 364294 589442 364350
rect 589498 364294 589566 364350
rect 589622 364294 596496 364350
rect 596552 364294 596620 364350
rect 596676 364294 596744 364350
rect 596800 364294 596868 364350
rect 596924 364294 597980 364350
rect -1916 364226 597980 364294
rect -1916 364170 -860 364226
rect -804 364170 -736 364226
rect -680 364170 -612 364226
rect -556 364170 -488 364226
rect -432 364170 5514 364226
rect 5570 364170 5638 364226
rect 5694 364170 5762 364226
rect 5818 364170 5886 364226
rect 5942 364170 36234 364226
rect 36290 364170 36358 364226
rect 36414 364170 36482 364226
rect 36538 364170 36606 364226
rect 36662 364170 66954 364226
rect 67010 364170 67078 364226
rect 67134 364170 67202 364226
rect 67258 364170 67326 364226
rect 67382 364170 97674 364226
rect 97730 364170 97798 364226
rect 97854 364170 97922 364226
rect 97978 364170 98046 364226
rect 98102 364170 128394 364226
rect 128450 364170 128518 364226
rect 128574 364170 128642 364226
rect 128698 364170 128766 364226
rect 128822 364170 159114 364226
rect 159170 364170 159238 364226
rect 159294 364170 159362 364226
rect 159418 364170 159486 364226
rect 159542 364170 189834 364226
rect 189890 364170 189958 364226
rect 190014 364170 190082 364226
rect 190138 364170 190206 364226
rect 190262 364170 220554 364226
rect 220610 364170 220678 364226
rect 220734 364170 220802 364226
rect 220858 364170 220926 364226
rect 220982 364170 251274 364226
rect 251330 364170 251398 364226
rect 251454 364170 251522 364226
rect 251578 364170 251646 364226
rect 251702 364170 281994 364226
rect 282050 364170 282118 364226
rect 282174 364170 282242 364226
rect 282298 364170 282366 364226
rect 282422 364170 312714 364226
rect 312770 364170 312838 364226
rect 312894 364170 312962 364226
rect 313018 364170 313086 364226
rect 313142 364170 343434 364226
rect 343490 364170 343558 364226
rect 343614 364170 343682 364226
rect 343738 364170 343806 364226
rect 343862 364170 374154 364226
rect 374210 364170 374278 364226
rect 374334 364170 374402 364226
rect 374458 364170 374526 364226
rect 374582 364170 404874 364226
rect 404930 364170 404998 364226
rect 405054 364170 405122 364226
rect 405178 364170 405246 364226
rect 405302 364170 435594 364226
rect 435650 364170 435718 364226
rect 435774 364170 435842 364226
rect 435898 364170 435966 364226
rect 436022 364170 466314 364226
rect 466370 364170 466438 364226
rect 466494 364170 466562 364226
rect 466618 364170 466686 364226
rect 466742 364170 497034 364226
rect 497090 364170 497158 364226
rect 497214 364170 497282 364226
rect 497338 364170 497406 364226
rect 497462 364170 527754 364226
rect 527810 364170 527878 364226
rect 527934 364170 528002 364226
rect 528058 364170 528126 364226
rect 528182 364170 558474 364226
rect 558530 364170 558598 364226
rect 558654 364170 558722 364226
rect 558778 364170 558846 364226
rect 558902 364170 589194 364226
rect 589250 364170 589318 364226
rect 589374 364170 589442 364226
rect 589498 364170 589566 364226
rect 589622 364170 596496 364226
rect 596552 364170 596620 364226
rect 596676 364170 596744 364226
rect 596800 364170 596868 364226
rect 596924 364170 597980 364226
rect -1916 364102 597980 364170
rect -1916 364046 -860 364102
rect -804 364046 -736 364102
rect -680 364046 -612 364102
rect -556 364046 -488 364102
rect -432 364046 5514 364102
rect 5570 364046 5638 364102
rect 5694 364046 5762 364102
rect 5818 364046 5886 364102
rect 5942 364046 36234 364102
rect 36290 364046 36358 364102
rect 36414 364046 36482 364102
rect 36538 364046 36606 364102
rect 36662 364046 66954 364102
rect 67010 364046 67078 364102
rect 67134 364046 67202 364102
rect 67258 364046 67326 364102
rect 67382 364046 97674 364102
rect 97730 364046 97798 364102
rect 97854 364046 97922 364102
rect 97978 364046 98046 364102
rect 98102 364046 128394 364102
rect 128450 364046 128518 364102
rect 128574 364046 128642 364102
rect 128698 364046 128766 364102
rect 128822 364046 159114 364102
rect 159170 364046 159238 364102
rect 159294 364046 159362 364102
rect 159418 364046 159486 364102
rect 159542 364046 189834 364102
rect 189890 364046 189958 364102
rect 190014 364046 190082 364102
rect 190138 364046 190206 364102
rect 190262 364046 220554 364102
rect 220610 364046 220678 364102
rect 220734 364046 220802 364102
rect 220858 364046 220926 364102
rect 220982 364046 251274 364102
rect 251330 364046 251398 364102
rect 251454 364046 251522 364102
rect 251578 364046 251646 364102
rect 251702 364046 281994 364102
rect 282050 364046 282118 364102
rect 282174 364046 282242 364102
rect 282298 364046 282366 364102
rect 282422 364046 312714 364102
rect 312770 364046 312838 364102
rect 312894 364046 312962 364102
rect 313018 364046 313086 364102
rect 313142 364046 343434 364102
rect 343490 364046 343558 364102
rect 343614 364046 343682 364102
rect 343738 364046 343806 364102
rect 343862 364046 374154 364102
rect 374210 364046 374278 364102
rect 374334 364046 374402 364102
rect 374458 364046 374526 364102
rect 374582 364046 404874 364102
rect 404930 364046 404998 364102
rect 405054 364046 405122 364102
rect 405178 364046 405246 364102
rect 405302 364046 435594 364102
rect 435650 364046 435718 364102
rect 435774 364046 435842 364102
rect 435898 364046 435966 364102
rect 436022 364046 466314 364102
rect 466370 364046 466438 364102
rect 466494 364046 466562 364102
rect 466618 364046 466686 364102
rect 466742 364046 497034 364102
rect 497090 364046 497158 364102
rect 497214 364046 497282 364102
rect 497338 364046 497406 364102
rect 497462 364046 527754 364102
rect 527810 364046 527878 364102
rect 527934 364046 528002 364102
rect 528058 364046 528126 364102
rect 528182 364046 558474 364102
rect 558530 364046 558598 364102
rect 558654 364046 558722 364102
rect 558778 364046 558846 364102
rect 558902 364046 589194 364102
rect 589250 364046 589318 364102
rect 589374 364046 589442 364102
rect 589498 364046 589566 364102
rect 589622 364046 596496 364102
rect 596552 364046 596620 364102
rect 596676 364046 596744 364102
rect 596800 364046 596868 364102
rect 596924 364046 597980 364102
rect -1916 363978 597980 364046
rect -1916 363922 -860 363978
rect -804 363922 -736 363978
rect -680 363922 -612 363978
rect -556 363922 -488 363978
rect -432 363922 5514 363978
rect 5570 363922 5638 363978
rect 5694 363922 5762 363978
rect 5818 363922 5886 363978
rect 5942 363922 36234 363978
rect 36290 363922 36358 363978
rect 36414 363922 36482 363978
rect 36538 363922 36606 363978
rect 36662 363922 66954 363978
rect 67010 363922 67078 363978
rect 67134 363922 67202 363978
rect 67258 363922 67326 363978
rect 67382 363922 97674 363978
rect 97730 363922 97798 363978
rect 97854 363922 97922 363978
rect 97978 363922 98046 363978
rect 98102 363922 128394 363978
rect 128450 363922 128518 363978
rect 128574 363922 128642 363978
rect 128698 363922 128766 363978
rect 128822 363922 159114 363978
rect 159170 363922 159238 363978
rect 159294 363922 159362 363978
rect 159418 363922 159486 363978
rect 159542 363922 189834 363978
rect 189890 363922 189958 363978
rect 190014 363922 190082 363978
rect 190138 363922 190206 363978
rect 190262 363922 220554 363978
rect 220610 363922 220678 363978
rect 220734 363922 220802 363978
rect 220858 363922 220926 363978
rect 220982 363922 251274 363978
rect 251330 363922 251398 363978
rect 251454 363922 251522 363978
rect 251578 363922 251646 363978
rect 251702 363922 281994 363978
rect 282050 363922 282118 363978
rect 282174 363922 282242 363978
rect 282298 363922 282366 363978
rect 282422 363922 312714 363978
rect 312770 363922 312838 363978
rect 312894 363922 312962 363978
rect 313018 363922 313086 363978
rect 313142 363922 343434 363978
rect 343490 363922 343558 363978
rect 343614 363922 343682 363978
rect 343738 363922 343806 363978
rect 343862 363922 374154 363978
rect 374210 363922 374278 363978
rect 374334 363922 374402 363978
rect 374458 363922 374526 363978
rect 374582 363922 404874 363978
rect 404930 363922 404998 363978
rect 405054 363922 405122 363978
rect 405178 363922 405246 363978
rect 405302 363922 435594 363978
rect 435650 363922 435718 363978
rect 435774 363922 435842 363978
rect 435898 363922 435966 363978
rect 436022 363922 466314 363978
rect 466370 363922 466438 363978
rect 466494 363922 466562 363978
rect 466618 363922 466686 363978
rect 466742 363922 497034 363978
rect 497090 363922 497158 363978
rect 497214 363922 497282 363978
rect 497338 363922 497406 363978
rect 497462 363922 527754 363978
rect 527810 363922 527878 363978
rect 527934 363922 528002 363978
rect 528058 363922 528126 363978
rect 528182 363922 558474 363978
rect 558530 363922 558598 363978
rect 558654 363922 558722 363978
rect 558778 363922 558846 363978
rect 558902 363922 589194 363978
rect 589250 363922 589318 363978
rect 589374 363922 589442 363978
rect 589498 363922 589566 363978
rect 589622 363922 596496 363978
rect 596552 363922 596620 363978
rect 596676 363922 596744 363978
rect 596800 363922 596868 363978
rect 596924 363922 597980 363978
rect -1916 363826 597980 363922
rect -1916 352350 597980 352446
rect -1916 352294 -1820 352350
rect -1764 352294 -1696 352350
rect -1640 352294 -1572 352350
rect -1516 352294 -1448 352350
rect -1392 352294 9234 352350
rect 9290 352294 9358 352350
rect 9414 352294 9482 352350
rect 9538 352294 9606 352350
rect 9662 352294 39954 352350
rect 40010 352294 40078 352350
rect 40134 352294 40202 352350
rect 40258 352294 40326 352350
rect 40382 352294 70674 352350
rect 70730 352294 70798 352350
rect 70854 352294 70922 352350
rect 70978 352294 71046 352350
rect 71102 352294 101394 352350
rect 101450 352294 101518 352350
rect 101574 352294 101642 352350
rect 101698 352294 101766 352350
rect 101822 352294 132114 352350
rect 132170 352294 132238 352350
rect 132294 352294 132362 352350
rect 132418 352294 132486 352350
rect 132542 352294 162834 352350
rect 162890 352294 162958 352350
rect 163014 352294 163082 352350
rect 163138 352294 163206 352350
rect 163262 352294 193554 352350
rect 193610 352294 193678 352350
rect 193734 352294 193802 352350
rect 193858 352294 193926 352350
rect 193982 352294 224274 352350
rect 224330 352294 224398 352350
rect 224454 352294 224522 352350
rect 224578 352294 224646 352350
rect 224702 352294 254994 352350
rect 255050 352294 255118 352350
rect 255174 352294 255242 352350
rect 255298 352294 255366 352350
rect 255422 352294 285714 352350
rect 285770 352294 285838 352350
rect 285894 352294 285962 352350
rect 286018 352294 286086 352350
rect 286142 352294 316434 352350
rect 316490 352294 316558 352350
rect 316614 352294 316682 352350
rect 316738 352294 316806 352350
rect 316862 352294 347154 352350
rect 347210 352294 347278 352350
rect 347334 352294 347402 352350
rect 347458 352294 347526 352350
rect 347582 352294 377874 352350
rect 377930 352294 377998 352350
rect 378054 352294 378122 352350
rect 378178 352294 378246 352350
rect 378302 352294 408594 352350
rect 408650 352294 408718 352350
rect 408774 352294 408842 352350
rect 408898 352294 408966 352350
rect 409022 352294 439314 352350
rect 439370 352294 439438 352350
rect 439494 352294 439562 352350
rect 439618 352294 439686 352350
rect 439742 352294 470034 352350
rect 470090 352294 470158 352350
rect 470214 352294 470282 352350
rect 470338 352294 470406 352350
rect 470462 352294 500754 352350
rect 500810 352294 500878 352350
rect 500934 352294 501002 352350
rect 501058 352294 501126 352350
rect 501182 352294 531474 352350
rect 531530 352294 531598 352350
rect 531654 352294 531722 352350
rect 531778 352294 531846 352350
rect 531902 352294 562194 352350
rect 562250 352294 562318 352350
rect 562374 352294 562442 352350
rect 562498 352294 562566 352350
rect 562622 352294 592914 352350
rect 592970 352294 593038 352350
rect 593094 352294 593162 352350
rect 593218 352294 593286 352350
rect 593342 352294 597456 352350
rect 597512 352294 597580 352350
rect 597636 352294 597704 352350
rect 597760 352294 597828 352350
rect 597884 352294 597980 352350
rect -1916 352226 597980 352294
rect -1916 352170 -1820 352226
rect -1764 352170 -1696 352226
rect -1640 352170 -1572 352226
rect -1516 352170 -1448 352226
rect -1392 352170 9234 352226
rect 9290 352170 9358 352226
rect 9414 352170 9482 352226
rect 9538 352170 9606 352226
rect 9662 352170 39954 352226
rect 40010 352170 40078 352226
rect 40134 352170 40202 352226
rect 40258 352170 40326 352226
rect 40382 352170 70674 352226
rect 70730 352170 70798 352226
rect 70854 352170 70922 352226
rect 70978 352170 71046 352226
rect 71102 352170 101394 352226
rect 101450 352170 101518 352226
rect 101574 352170 101642 352226
rect 101698 352170 101766 352226
rect 101822 352170 132114 352226
rect 132170 352170 132238 352226
rect 132294 352170 132362 352226
rect 132418 352170 132486 352226
rect 132542 352170 162834 352226
rect 162890 352170 162958 352226
rect 163014 352170 163082 352226
rect 163138 352170 163206 352226
rect 163262 352170 193554 352226
rect 193610 352170 193678 352226
rect 193734 352170 193802 352226
rect 193858 352170 193926 352226
rect 193982 352170 224274 352226
rect 224330 352170 224398 352226
rect 224454 352170 224522 352226
rect 224578 352170 224646 352226
rect 224702 352170 254994 352226
rect 255050 352170 255118 352226
rect 255174 352170 255242 352226
rect 255298 352170 255366 352226
rect 255422 352170 285714 352226
rect 285770 352170 285838 352226
rect 285894 352170 285962 352226
rect 286018 352170 286086 352226
rect 286142 352170 316434 352226
rect 316490 352170 316558 352226
rect 316614 352170 316682 352226
rect 316738 352170 316806 352226
rect 316862 352170 347154 352226
rect 347210 352170 347278 352226
rect 347334 352170 347402 352226
rect 347458 352170 347526 352226
rect 347582 352170 377874 352226
rect 377930 352170 377998 352226
rect 378054 352170 378122 352226
rect 378178 352170 378246 352226
rect 378302 352170 408594 352226
rect 408650 352170 408718 352226
rect 408774 352170 408842 352226
rect 408898 352170 408966 352226
rect 409022 352170 439314 352226
rect 439370 352170 439438 352226
rect 439494 352170 439562 352226
rect 439618 352170 439686 352226
rect 439742 352170 470034 352226
rect 470090 352170 470158 352226
rect 470214 352170 470282 352226
rect 470338 352170 470406 352226
rect 470462 352170 500754 352226
rect 500810 352170 500878 352226
rect 500934 352170 501002 352226
rect 501058 352170 501126 352226
rect 501182 352170 531474 352226
rect 531530 352170 531598 352226
rect 531654 352170 531722 352226
rect 531778 352170 531846 352226
rect 531902 352170 562194 352226
rect 562250 352170 562318 352226
rect 562374 352170 562442 352226
rect 562498 352170 562566 352226
rect 562622 352170 592914 352226
rect 592970 352170 593038 352226
rect 593094 352170 593162 352226
rect 593218 352170 593286 352226
rect 593342 352170 597456 352226
rect 597512 352170 597580 352226
rect 597636 352170 597704 352226
rect 597760 352170 597828 352226
rect 597884 352170 597980 352226
rect -1916 352102 597980 352170
rect -1916 352046 -1820 352102
rect -1764 352046 -1696 352102
rect -1640 352046 -1572 352102
rect -1516 352046 -1448 352102
rect -1392 352046 9234 352102
rect 9290 352046 9358 352102
rect 9414 352046 9482 352102
rect 9538 352046 9606 352102
rect 9662 352046 39954 352102
rect 40010 352046 40078 352102
rect 40134 352046 40202 352102
rect 40258 352046 40326 352102
rect 40382 352046 70674 352102
rect 70730 352046 70798 352102
rect 70854 352046 70922 352102
rect 70978 352046 71046 352102
rect 71102 352046 101394 352102
rect 101450 352046 101518 352102
rect 101574 352046 101642 352102
rect 101698 352046 101766 352102
rect 101822 352046 132114 352102
rect 132170 352046 132238 352102
rect 132294 352046 132362 352102
rect 132418 352046 132486 352102
rect 132542 352046 162834 352102
rect 162890 352046 162958 352102
rect 163014 352046 163082 352102
rect 163138 352046 163206 352102
rect 163262 352046 193554 352102
rect 193610 352046 193678 352102
rect 193734 352046 193802 352102
rect 193858 352046 193926 352102
rect 193982 352046 224274 352102
rect 224330 352046 224398 352102
rect 224454 352046 224522 352102
rect 224578 352046 224646 352102
rect 224702 352046 254994 352102
rect 255050 352046 255118 352102
rect 255174 352046 255242 352102
rect 255298 352046 255366 352102
rect 255422 352046 285714 352102
rect 285770 352046 285838 352102
rect 285894 352046 285962 352102
rect 286018 352046 286086 352102
rect 286142 352046 316434 352102
rect 316490 352046 316558 352102
rect 316614 352046 316682 352102
rect 316738 352046 316806 352102
rect 316862 352046 347154 352102
rect 347210 352046 347278 352102
rect 347334 352046 347402 352102
rect 347458 352046 347526 352102
rect 347582 352046 377874 352102
rect 377930 352046 377998 352102
rect 378054 352046 378122 352102
rect 378178 352046 378246 352102
rect 378302 352046 408594 352102
rect 408650 352046 408718 352102
rect 408774 352046 408842 352102
rect 408898 352046 408966 352102
rect 409022 352046 439314 352102
rect 439370 352046 439438 352102
rect 439494 352046 439562 352102
rect 439618 352046 439686 352102
rect 439742 352046 470034 352102
rect 470090 352046 470158 352102
rect 470214 352046 470282 352102
rect 470338 352046 470406 352102
rect 470462 352046 500754 352102
rect 500810 352046 500878 352102
rect 500934 352046 501002 352102
rect 501058 352046 501126 352102
rect 501182 352046 531474 352102
rect 531530 352046 531598 352102
rect 531654 352046 531722 352102
rect 531778 352046 531846 352102
rect 531902 352046 562194 352102
rect 562250 352046 562318 352102
rect 562374 352046 562442 352102
rect 562498 352046 562566 352102
rect 562622 352046 592914 352102
rect 592970 352046 593038 352102
rect 593094 352046 593162 352102
rect 593218 352046 593286 352102
rect 593342 352046 597456 352102
rect 597512 352046 597580 352102
rect 597636 352046 597704 352102
rect 597760 352046 597828 352102
rect 597884 352046 597980 352102
rect -1916 351978 597980 352046
rect -1916 351922 -1820 351978
rect -1764 351922 -1696 351978
rect -1640 351922 -1572 351978
rect -1516 351922 -1448 351978
rect -1392 351922 9234 351978
rect 9290 351922 9358 351978
rect 9414 351922 9482 351978
rect 9538 351922 9606 351978
rect 9662 351922 39954 351978
rect 40010 351922 40078 351978
rect 40134 351922 40202 351978
rect 40258 351922 40326 351978
rect 40382 351922 70674 351978
rect 70730 351922 70798 351978
rect 70854 351922 70922 351978
rect 70978 351922 71046 351978
rect 71102 351922 101394 351978
rect 101450 351922 101518 351978
rect 101574 351922 101642 351978
rect 101698 351922 101766 351978
rect 101822 351922 132114 351978
rect 132170 351922 132238 351978
rect 132294 351922 132362 351978
rect 132418 351922 132486 351978
rect 132542 351922 162834 351978
rect 162890 351922 162958 351978
rect 163014 351922 163082 351978
rect 163138 351922 163206 351978
rect 163262 351922 193554 351978
rect 193610 351922 193678 351978
rect 193734 351922 193802 351978
rect 193858 351922 193926 351978
rect 193982 351922 224274 351978
rect 224330 351922 224398 351978
rect 224454 351922 224522 351978
rect 224578 351922 224646 351978
rect 224702 351922 254994 351978
rect 255050 351922 255118 351978
rect 255174 351922 255242 351978
rect 255298 351922 255366 351978
rect 255422 351922 285714 351978
rect 285770 351922 285838 351978
rect 285894 351922 285962 351978
rect 286018 351922 286086 351978
rect 286142 351922 316434 351978
rect 316490 351922 316558 351978
rect 316614 351922 316682 351978
rect 316738 351922 316806 351978
rect 316862 351922 347154 351978
rect 347210 351922 347278 351978
rect 347334 351922 347402 351978
rect 347458 351922 347526 351978
rect 347582 351922 377874 351978
rect 377930 351922 377998 351978
rect 378054 351922 378122 351978
rect 378178 351922 378246 351978
rect 378302 351922 408594 351978
rect 408650 351922 408718 351978
rect 408774 351922 408842 351978
rect 408898 351922 408966 351978
rect 409022 351922 439314 351978
rect 439370 351922 439438 351978
rect 439494 351922 439562 351978
rect 439618 351922 439686 351978
rect 439742 351922 470034 351978
rect 470090 351922 470158 351978
rect 470214 351922 470282 351978
rect 470338 351922 470406 351978
rect 470462 351922 500754 351978
rect 500810 351922 500878 351978
rect 500934 351922 501002 351978
rect 501058 351922 501126 351978
rect 501182 351922 531474 351978
rect 531530 351922 531598 351978
rect 531654 351922 531722 351978
rect 531778 351922 531846 351978
rect 531902 351922 562194 351978
rect 562250 351922 562318 351978
rect 562374 351922 562442 351978
rect 562498 351922 562566 351978
rect 562622 351922 592914 351978
rect 592970 351922 593038 351978
rect 593094 351922 593162 351978
rect 593218 351922 593286 351978
rect 593342 351922 597456 351978
rect 597512 351922 597580 351978
rect 597636 351922 597704 351978
rect 597760 351922 597828 351978
rect 597884 351922 597980 351978
rect -1916 351826 597980 351922
rect -1916 346350 597980 346446
rect -1916 346294 -860 346350
rect -804 346294 -736 346350
rect -680 346294 -612 346350
rect -556 346294 -488 346350
rect -432 346294 5514 346350
rect 5570 346294 5638 346350
rect 5694 346294 5762 346350
rect 5818 346294 5886 346350
rect 5942 346294 36234 346350
rect 36290 346294 36358 346350
rect 36414 346294 36482 346350
rect 36538 346294 36606 346350
rect 36662 346294 66954 346350
rect 67010 346294 67078 346350
rect 67134 346294 67202 346350
rect 67258 346294 67326 346350
rect 67382 346294 97674 346350
rect 97730 346294 97798 346350
rect 97854 346294 97922 346350
rect 97978 346294 98046 346350
rect 98102 346294 128394 346350
rect 128450 346294 128518 346350
rect 128574 346294 128642 346350
rect 128698 346294 128766 346350
rect 128822 346294 159114 346350
rect 159170 346294 159238 346350
rect 159294 346294 159362 346350
rect 159418 346294 159486 346350
rect 159542 346294 189834 346350
rect 189890 346294 189958 346350
rect 190014 346294 190082 346350
rect 190138 346294 190206 346350
rect 190262 346294 220554 346350
rect 220610 346294 220678 346350
rect 220734 346294 220802 346350
rect 220858 346294 220926 346350
rect 220982 346294 251274 346350
rect 251330 346294 251398 346350
rect 251454 346294 251522 346350
rect 251578 346294 251646 346350
rect 251702 346294 281994 346350
rect 282050 346294 282118 346350
rect 282174 346294 282242 346350
rect 282298 346294 282366 346350
rect 282422 346294 312714 346350
rect 312770 346294 312838 346350
rect 312894 346294 312962 346350
rect 313018 346294 313086 346350
rect 313142 346294 343434 346350
rect 343490 346294 343558 346350
rect 343614 346294 343682 346350
rect 343738 346294 343806 346350
rect 343862 346294 374154 346350
rect 374210 346294 374278 346350
rect 374334 346294 374402 346350
rect 374458 346294 374526 346350
rect 374582 346294 404874 346350
rect 404930 346294 404998 346350
rect 405054 346294 405122 346350
rect 405178 346294 405246 346350
rect 405302 346294 435594 346350
rect 435650 346294 435718 346350
rect 435774 346294 435842 346350
rect 435898 346294 435966 346350
rect 436022 346294 466314 346350
rect 466370 346294 466438 346350
rect 466494 346294 466562 346350
rect 466618 346294 466686 346350
rect 466742 346294 497034 346350
rect 497090 346294 497158 346350
rect 497214 346294 497282 346350
rect 497338 346294 497406 346350
rect 497462 346294 527754 346350
rect 527810 346294 527878 346350
rect 527934 346294 528002 346350
rect 528058 346294 528126 346350
rect 528182 346294 558474 346350
rect 558530 346294 558598 346350
rect 558654 346294 558722 346350
rect 558778 346294 558846 346350
rect 558902 346294 589194 346350
rect 589250 346294 589318 346350
rect 589374 346294 589442 346350
rect 589498 346294 589566 346350
rect 589622 346294 596496 346350
rect 596552 346294 596620 346350
rect 596676 346294 596744 346350
rect 596800 346294 596868 346350
rect 596924 346294 597980 346350
rect -1916 346226 597980 346294
rect -1916 346170 -860 346226
rect -804 346170 -736 346226
rect -680 346170 -612 346226
rect -556 346170 -488 346226
rect -432 346170 5514 346226
rect 5570 346170 5638 346226
rect 5694 346170 5762 346226
rect 5818 346170 5886 346226
rect 5942 346170 36234 346226
rect 36290 346170 36358 346226
rect 36414 346170 36482 346226
rect 36538 346170 36606 346226
rect 36662 346170 66954 346226
rect 67010 346170 67078 346226
rect 67134 346170 67202 346226
rect 67258 346170 67326 346226
rect 67382 346170 97674 346226
rect 97730 346170 97798 346226
rect 97854 346170 97922 346226
rect 97978 346170 98046 346226
rect 98102 346170 128394 346226
rect 128450 346170 128518 346226
rect 128574 346170 128642 346226
rect 128698 346170 128766 346226
rect 128822 346170 159114 346226
rect 159170 346170 159238 346226
rect 159294 346170 159362 346226
rect 159418 346170 159486 346226
rect 159542 346170 189834 346226
rect 189890 346170 189958 346226
rect 190014 346170 190082 346226
rect 190138 346170 190206 346226
rect 190262 346170 220554 346226
rect 220610 346170 220678 346226
rect 220734 346170 220802 346226
rect 220858 346170 220926 346226
rect 220982 346170 251274 346226
rect 251330 346170 251398 346226
rect 251454 346170 251522 346226
rect 251578 346170 251646 346226
rect 251702 346170 281994 346226
rect 282050 346170 282118 346226
rect 282174 346170 282242 346226
rect 282298 346170 282366 346226
rect 282422 346170 312714 346226
rect 312770 346170 312838 346226
rect 312894 346170 312962 346226
rect 313018 346170 313086 346226
rect 313142 346170 343434 346226
rect 343490 346170 343558 346226
rect 343614 346170 343682 346226
rect 343738 346170 343806 346226
rect 343862 346170 374154 346226
rect 374210 346170 374278 346226
rect 374334 346170 374402 346226
rect 374458 346170 374526 346226
rect 374582 346170 404874 346226
rect 404930 346170 404998 346226
rect 405054 346170 405122 346226
rect 405178 346170 405246 346226
rect 405302 346170 435594 346226
rect 435650 346170 435718 346226
rect 435774 346170 435842 346226
rect 435898 346170 435966 346226
rect 436022 346170 466314 346226
rect 466370 346170 466438 346226
rect 466494 346170 466562 346226
rect 466618 346170 466686 346226
rect 466742 346170 497034 346226
rect 497090 346170 497158 346226
rect 497214 346170 497282 346226
rect 497338 346170 497406 346226
rect 497462 346170 527754 346226
rect 527810 346170 527878 346226
rect 527934 346170 528002 346226
rect 528058 346170 528126 346226
rect 528182 346170 558474 346226
rect 558530 346170 558598 346226
rect 558654 346170 558722 346226
rect 558778 346170 558846 346226
rect 558902 346170 589194 346226
rect 589250 346170 589318 346226
rect 589374 346170 589442 346226
rect 589498 346170 589566 346226
rect 589622 346170 596496 346226
rect 596552 346170 596620 346226
rect 596676 346170 596744 346226
rect 596800 346170 596868 346226
rect 596924 346170 597980 346226
rect -1916 346102 597980 346170
rect -1916 346046 -860 346102
rect -804 346046 -736 346102
rect -680 346046 -612 346102
rect -556 346046 -488 346102
rect -432 346046 5514 346102
rect 5570 346046 5638 346102
rect 5694 346046 5762 346102
rect 5818 346046 5886 346102
rect 5942 346046 36234 346102
rect 36290 346046 36358 346102
rect 36414 346046 36482 346102
rect 36538 346046 36606 346102
rect 36662 346046 66954 346102
rect 67010 346046 67078 346102
rect 67134 346046 67202 346102
rect 67258 346046 67326 346102
rect 67382 346046 97674 346102
rect 97730 346046 97798 346102
rect 97854 346046 97922 346102
rect 97978 346046 98046 346102
rect 98102 346046 128394 346102
rect 128450 346046 128518 346102
rect 128574 346046 128642 346102
rect 128698 346046 128766 346102
rect 128822 346046 159114 346102
rect 159170 346046 159238 346102
rect 159294 346046 159362 346102
rect 159418 346046 159486 346102
rect 159542 346046 189834 346102
rect 189890 346046 189958 346102
rect 190014 346046 190082 346102
rect 190138 346046 190206 346102
rect 190262 346046 220554 346102
rect 220610 346046 220678 346102
rect 220734 346046 220802 346102
rect 220858 346046 220926 346102
rect 220982 346046 251274 346102
rect 251330 346046 251398 346102
rect 251454 346046 251522 346102
rect 251578 346046 251646 346102
rect 251702 346046 281994 346102
rect 282050 346046 282118 346102
rect 282174 346046 282242 346102
rect 282298 346046 282366 346102
rect 282422 346046 312714 346102
rect 312770 346046 312838 346102
rect 312894 346046 312962 346102
rect 313018 346046 313086 346102
rect 313142 346046 343434 346102
rect 343490 346046 343558 346102
rect 343614 346046 343682 346102
rect 343738 346046 343806 346102
rect 343862 346046 374154 346102
rect 374210 346046 374278 346102
rect 374334 346046 374402 346102
rect 374458 346046 374526 346102
rect 374582 346046 404874 346102
rect 404930 346046 404998 346102
rect 405054 346046 405122 346102
rect 405178 346046 405246 346102
rect 405302 346046 435594 346102
rect 435650 346046 435718 346102
rect 435774 346046 435842 346102
rect 435898 346046 435966 346102
rect 436022 346046 466314 346102
rect 466370 346046 466438 346102
rect 466494 346046 466562 346102
rect 466618 346046 466686 346102
rect 466742 346046 497034 346102
rect 497090 346046 497158 346102
rect 497214 346046 497282 346102
rect 497338 346046 497406 346102
rect 497462 346046 527754 346102
rect 527810 346046 527878 346102
rect 527934 346046 528002 346102
rect 528058 346046 528126 346102
rect 528182 346046 558474 346102
rect 558530 346046 558598 346102
rect 558654 346046 558722 346102
rect 558778 346046 558846 346102
rect 558902 346046 589194 346102
rect 589250 346046 589318 346102
rect 589374 346046 589442 346102
rect 589498 346046 589566 346102
rect 589622 346046 596496 346102
rect 596552 346046 596620 346102
rect 596676 346046 596744 346102
rect 596800 346046 596868 346102
rect 596924 346046 597980 346102
rect -1916 345978 597980 346046
rect -1916 345922 -860 345978
rect -804 345922 -736 345978
rect -680 345922 -612 345978
rect -556 345922 -488 345978
rect -432 345922 5514 345978
rect 5570 345922 5638 345978
rect 5694 345922 5762 345978
rect 5818 345922 5886 345978
rect 5942 345922 36234 345978
rect 36290 345922 36358 345978
rect 36414 345922 36482 345978
rect 36538 345922 36606 345978
rect 36662 345922 66954 345978
rect 67010 345922 67078 345978
rect 67134 345922 67202 345978
rect 67258 345922 67326 345978
rect 67382 345922 97674 345978
rect 97730 345922 97798 345978
rect 97854 345922 97922 345978
rect 97978 345922 98046 345978
rect 98102 345922 128394 345978
rect 128450 345922 128518 345978
rect 128574 345922 128642 345978
rect 128698 345922 128766 345978
rect 128822 345922 159114 345978
rect 159170 345922 159238 345978
rect 159294 345922 159362 345978
rect 159418 345922 159486 345978
rect 159542 345922 189834 345978
rect 189890 345922 189958 345978
rect 190014 345922 190082 345978
rect 190138 345922 190206 345978
rect 190262 345922 220554 345978
rect 220610 345922 220678 345978
rect 220734 345922 220802 345978
rect 220858 345922 220926 345978
rect 220982 345922 251274 345978
rect 251330 345922 251398 345978
rect 251454 345922 251522 345978
rect 251578 345922 251646 345978
rect 251702 345922 281994 345978
rect 282050 345922 282118 345978
rect 282174 345922 282242 345978
rect 282298 345922 282366 345978
rect 282422 345922 312714 345978
rect 312770 345922 312838 345978
rect 312894 345922 312962 345978
rect 313018 345922 313086 345978
rect 313142 345922 343434 345978
rect 343490 345922 343558 345978
rect 343614 345922 343682 345978
rect 343738 345922 343806 345978
rect 343862 345922 374154 345978
rect 374210 345922 374278 345978
rect 374334 345922 374402 345978
rect 374458 345922 374526 345978
rect 374582 345922 404874 345978
rect 404930 345922 404998 345978
rect 405054 345922 405122 345978
rect 405178 345922 405246 345978
rect 405302 345922 435594 345978
rect 435650 345922 435718 345978
rect 435774 345922 435842 345978
rect 435898 345922 435966 345978
rect 436022 345922 466314 345978
rect 466370 345922 466438 345978
rect 466494 345922 466562 345978
rect 466618 345922 466686 345978
rect 466742 345922 497034 345978
rect 497090 345922 497158 345978
rect 497214 345922 497282 345978
rect 497338 345922 497406 345978
rect 497462 345922 527754 345978
rect 527810 345922 527878 345978
rect 527934 345922 528002 345978
rect 528058 345922 528126 345978
rect 528182 345922 558474 345978
rect 558530 345922 558598 345978
rect 558654 345922 558722 345978
rect 558778 345922 558846 345978
rect 558902 345922 589194 345978
rect 589250 345922 589318 345978
rect 589374 345922 589442 345978
rect 589498 345922 589566 345978
rect 589622 345922 596496 345978
rect 596552 345922 596620 345978
rect 596676 345922 596744 345978
rect 596800 345922 596868 345978
rect 596924 345922 597980 345978
rect -1916 345826 597980 345922
rect -1916 334350 597980 334446
rect -1916 334294 -1820 334350
rect -1764 334294 -1696 334350
rect -1640 334294 -1572 334350
rect -1516 334294 -1448 334350
rect -1392 334294 9234 334350
rect 9290 334294 9358 334350
rect 9414 334294 9482 334350
rect 9538 334294 9606 334350
rect 9662 334294 39954 334350
rect 40010 334294 40078 334350
rect 40134 334294 40202 334350
rect 40258 334294 40326 334350
rect 40382 334294 70674 334350
rect 70730 334294 70798 334350
rect 70854 334294 70922 334350
rect 70978 334294 71046 334350
rect 71102 334294 101394 334350
rect 101450 334294 101518 334350
rect 101574 334294 101642 334350
rect 101698 334294 101766 334350
rect 101822 334294 132114 334350
rect 132170 334294 132238 334350
rect 132294 334294 132362 334350
rect 132418 334294 132486 334350
rect 132542 334294 162834 334350
rect 162890 334294 162958 334350
rect 163014 334294 163082 334350
rect 163138 334294 163206 334350
rect 163262 334294 193554 334350
rect 193610 334294 193678 334350
rect 193734 334294 193802 334350
rect 193858 334294 193926 334350
rect 193982 334294 224274 334350
rect 224330 334294 224398 334350
rect 224454 334294 224522 334350
rect 224578 334294 224646 334350
rect 224702 334294 254994 334350
rect 255050 334294 255118 334350
rect 255174 334294 255242 334350
rect 255298 334294 255366 334350
rect 255422 334294 285714 334350
rect 285770 334294 285838 334350
rect 285894 334294 285962 334350
rect 286018 334294 286086 334350
rect 286142 334294 316434 334350
rect 316490 334294 316558 334350
rect 316614 334294 316682 334350
rect 316738 334294 316806 334350
rect 316862 334294 347154 334350
rect 347210 334294 347278 334350
rect 347334 334294 347402 334350
rect 347458 334294 347526 334350
rect 347582 334294 377874 334350
rect 377930 334294 377998 334350
rect 378054 334294 378122 334350
rect 378178 334294 378246 334350
rect 378302 334294 408594 334350
rect 408650 334294 408718 334350
rect 408774 334294 408842 334350
rect 408898 334294 408966 334350
rect 409022 334294 439314 334350
rect 439370 334294 439438 334350
rect 439494 334294 439562 334350
rect 439618 334294 439686 334350
rect 439742 334294 470034 334350
rect 470090 334294 470158 334350
rect 470214 334294 470282 334350
rect 470338 334294 470406 334350
rect 470462 334294 500754 334350
rect 500810 334294 500878 334350
rect 500934 334294 501002 334350
rect 501058 334294 501126 334350
rect 501182 334294 531474 334350
rect 531530 334294 531598 334350
rect 531654 334294 531722 334350
rect 531778 334294 531846 334350
rect 531902 334294 562194 334350
rect 562250 334294 562318 334350
rect 562374 334294 562442 334350
rect 562498 334294 562566 334350
rect 562622 334294 592914 334350
rect 592970 334294 593038 334350
rect 593094 334294 593162 334350
rect 593218 334294 593286 334350
rect 593342 334294 597456 334350
rect 597512 334294 597580 334350
rect 597636 334294 597704 334350
rect 597760 334294 597828 334350
rect 597884 334294 597980 334350
rect -1916 334226 597980 334294
rect -1916 334170 -1820 334226
rect -1764 334170 -1696 334226
rect -1640 334170 -1572 334226
rect -1516 334170 -1448 334226
rect -1392 334170 9234 334226
rect 9290 334170 9358 334226
rect 9414 334170 9482 334226
rect 9538 334170 9606 334226
rect 9662 334170 39954 334226
rect 40010 334170 40078 334226
rect 40134 334170 40202 334226
rect 40258 334170 40326 334226
rect 40382 334170 70674 334226
rect 70730 334170 70798 334226
rect 70854 334170 70922 334226
rect 70978 334170 71046 334226
rect 71102 334170 101394 334226
rect 101450 334170 101518 334226
rect 101574 334170 101642 334226
rect 101698 334170 101766 334226
rect 101822 334170 132114 334226
rect 132170 334170 132238 334226
rect 132294 334170 132362 334226
rect 132418 334170 132486 334226
rect 132542 334170 162834 334226
rect 162890 334170 162958 334226
rect 163014 334170 163082 334226
rect 163138 334170 163206 334226
rect 163262 334170 193554 334226
rect 193610 334170 193678 334226
rect 193734 334170 193802 334226
rect 193858 334170 193926 334226
rect 193982 334170 224274 334226
rect 224330 334170 224398 334226
rect 224454 334170 224522 334226
rect 224578 334170 224646 334226
rect 224702 334170 254994 334226
rect 255050 334170 255118 334226
rect 255174 334170 255242 334226
rect 255298 334170 255366 334226
rect 255422 334170 285714 334226
rect 285770 334170 285838 334226
rect 285894 334170 285962 334226
rect 286018 334170 286086 334226
rect 286142 334170 316434 334226
rect 316490 334170 316558 334226
rect 316614 334170 316682 334226
rect 316738 334170 316806 334226
rect 316862 334170 347154 334226
rect 347210 334170 347278 334226
rect 347334 334170 347402 334226
rect 347458 334170 347526 334226
rect 347582 334170 377874 334226
rect 377930 334170 377998 334226
rect 378054 334170 378122 334226
rect 378178 334170 378246 334226
rect 378302 334170 408594 334226
rect 408650 334170 408718 334226
rect 408774 334170 408842 334226
rect 408898 334170 408966 334226
rect 409022 334170 439314 334226
rect 439370 334170 439438 334226
rect 439494 334170 439562 334226
rect 439618 334170 439686 334226
rect 439742 334170 470034 334226
rect 470090 334170 470158 334226
rect 470214 334170 470282 334226
rect 470338 334170 470406 334226
rect 470462 334170 500754 334226
rect 500810 334170 500878 334226
rect 500934 334170 501002 334226
rect 501058 334170 501126 334226
rect 501182 334170 531474 334226
rect 531530 334170 531598 334226
rect 531654 334170 531722 334226
rect 531778 334170 531846 334226
rect 531902 334170 562194 334226
rect 562250 334170 562318 334226
rect 562374 334170 562442 334226
rect 562498 334170 562566 334226
rect 562622 334170 592914 334226
rect 592970 334170 593038 334226
rect 593094 334170 593162 334226
rect 593218 334170 593286 334226
rect 593342 334170 597456 334226
rect 597512 334170 597580 334226
rect 597636 334170 597704 334226
rect 597760 334170 597828 334226
rect 597884 334170 597980 334226
rect -1916 334102 597980 334170
rect -1916 334046 -1820 334102
rect -1764 334046 -1696 334102
rect -1640 334046 -1572 334102
rect -1516 334046 -1448 334102
rect -1392 334046 9234 334102
rect 9290 334046 9358 334102
rect 9414 334046 9482 334102
rect 9538 334046 9606 334102
rect 9662 334046 39954 334102
rect 40010 334046 40078 334102
rect 40134 334046 40202 334102
rect 40258 334046 40326 334102
rect 40382 334046 70674 334102
rect 70730 334046 70798 334102
rect 70854 334046 70922 334102
rect 70978 334046 71046 334102
rect 71102 334046 101394 334102
rect 101450 334046 101518 334102
rect 101574 334046 101642 334102
rect 101698 334046 101766 334102
rect 101822 334046 132114 334102
rect 132170 334046 132238 334102
rect 132294 334046 132362 334102
rect 132418 334046 132486 334102
rect 132542 334046 162834 334102
rect 162890 334046 162958 334102
rect 163014 334046 163082 334102
rect 163138 334046 163206 334102
rect 163262 334046 193554 334102
rect 193610 334046 193678 334102
rect 193734 334046 193802 334102
rect 193858 334046 193926 334102
rect 193982 334046 224274 334102
rect 224330 334046 224398 334102
rect 224454 334046 224522 334102
rect 224578 334046 224646 334102
rect 224702 334046 254994 334102
rect 255050 334046 255118 334102
rect 255174 334046 255242 334102
rect 255298 334046 255366 334102
rect 255422 334046 285714 334102
rect 285770 334046 285838 334102
rect 285894 334046 285962 334102
rect 286018 334046 286086 334102
rect 286142 334046 316434 334102
rect 316490 334046 316558 334102
rect 316614 334046 316682 334102
rect 316738 334046 316806 334102
rect 316862 334046 347154 334102
rect 347210 334046 347278 334102
rect 347334 334046 347402 334102
rect 347458 334046 347526 334102
rect 347582 334046 377874 334102
rect 377930 334046 377998 334102
rect 378054 334046 378122 334102
rect 378178 334046 378246 334102
rect 378302 334046 408594 334102
rect 408650 334046 408718 334102
rect 408774 334046 408842 334102
rect 408898 334046 408966 334102
rect 409022 334046 439314 334102
rect 439370 334046 439438 334102
rect 439494 334046 439562 334102
rect 439618 334046 439686 334102
rect 439742 334046 470034 334102
rect 470090 334046 470158 334102
rect 470214 334046 470282 334102
rect 470338 334046 470406 334102
rect 470462 334046 500754 334102
rect 500810 334046 500878 334102
rect 500934 334046 501002 334102
rect 501058 334046 501126 334102
rect 501182 334046 531474 334102
rect 531530 334046 531598 334102
rect 531654 334046 531722 334102
rect 531778 334046 531846 334102
rect 531902 334046 562194 334102
rect 562250 334046 562318 334102
rect 562374 334046 562442 334102
rect 562498 334046 562566 334102
rect 562622 334046 592914 334102
rect 592970 334046 593038 334102
rect 593094 334046 593162 334102
rect 593218 334046 593286 334102
rect 593342 334046 597456 334102
rect 597512 334046 597580 334102
rect 597636 334046 597704 334102
rect 597760 334046 597828 334102
rect 597884 334046 597980 334102
rect -1916 333978 597980 334046
rect -1916 333922 -1820 333978
rect -1764 333922 -1696 333978
rect -1640 333922 -1572 333978
rect -1516 333922 -1448 333978
rect -1392 333922 9234 333978
rect 9290 333922 9358 333978
rect 9414 333922 9482 333978
rect 9538 333922 9606 333978
rect 9662 333922 39954 333978
rect 40010 333922 40078 333978
rect 40134 333922 40202 333978
rect 40258 333922 40326 333978
rect 40382 333922 70674 333978
rect 70730 333922 70798 333978
rect 70854 333922 70922 333978
rect 70978 333922 71046 333978
rect 71102 333922 101394 333978
rect 101450 333922 101518 333978
rect 101574 333922 101642 333978
rect 101698 333922 101766 333978
rect 101822 333922 132114 333978
rect 132170 333922 132238 333978
rect 132294 333922 132362 333978
rect 132418 333922 132486 333978
rect 132542 333922 162834 333978
rect 162890 333922 162958 333978
rect 163014 333922 163082 333978
rect 163138 333922 163206 333978
rect 163262 333922 193554 333978
rect 193610 333922 193678 333978
rect 193734 333922 193802 333978
rect 193858 333922 193926 333978
rect 193982 333922 224274 333978
rect 224330 333922 224398 333978
rect 224454 333922 224522 333978
rect 224578 333922 224646 333978
rect 224702 333922 254994 333978
rect 255050 333922 255118 333978
rect 255174 333922 255242 333978
rect 255298 333922 255366 333978
rect 255422 333922 285714 333978
rect 285770 333922 285838 333978
rect 285894 333922 285962 333978
rect 286018 333922 286086 333978
rect 286142 333922 316434 333978
rect 316490 333922 316558 333978
rect 316614 333922 316682 333978
rect 316738 333922 316806 333978
rect 316862 333922 347154 333978
rect 347210 333922 347278 333978
rect 347334 333922 347402 333978
rect 347458 333922 347526 333978
rect 347582 333922 377874 333978
rect 377930 333922 377998 333978
rect 378054 333922 378122 333978
rect 378178 333922 378246 333978
rect 378302 333922 408594 333978
rect 408650 333922 408718 333978
rect 408774 333922 408842 333978
rect 408898 333922 408966 333978
rect 409022 333922 439314 333978
rect 439370 333922 439438 333978
rect 439494 333922 439562 333978
rect 439618 333922 439686 333978
rect 439742 333922 470034 333978
rect 470090 333922 470158 333978
rect 470214 333922 470282 333978
rect 470338 333922 470406 333978
rect 470462 333922 500754 333978
rect 500810 333922 500878 333978
rect 500934 333922 501002 333978
rect 501058 333922 501126 333978
rect 501182 333922 531474 333978
rect 531530 333922 531598 333978
rect 531654 333922 531722 333978
rect 531778 333922 531846 333978
rect 531902 333922 562194 333978
rect 562250 333922 562318 333978
rect 562374 333922 562442 333978
rect 562498 333922 562566 333978
rect 562622 333922 592914 333978
rect 592970 333922 593038 333978
rect 593094 333922 593162 333978
rect 593218 333922 593286 333978
rect 593342 333922 597456 333978
rect 597512 333922 597580 333978
rect 597636 333922 597704 333978
rect 597760 333922 597828 333978
rect 597884 333922 597980 333978
rect -1916 333826 597980 333922
rect -1916 328350 597980 328446
rect -1916 328294 -860 328350
rect -804 328294 -736 328350
rect -680 328294 -612 328350
rect -556 328294 -488 328350
rect -432 328294 5514 328350
rect 5570 328294 5638 328350
rect 5694 328294 5762 328350
rect 5818 328294 5886 328350
rect 5942 328294 36234 328350
rect 36290 328294 36358 328350
rect 36414 328294 36482 328350
rect 36538 328294 36606 328350
rect 36662 328294 66954 328350
rect 67010 328294 67078 328350
rect 67134 328294 67202 328350
rect 67258 328294 67326 328350
rect 67382 328294 97674 328350
rect 97730 328294 97798 328350
rect 97854 328294 97922 328350
rect 97978 328294 98046 328350
rect 98102 328294 128394 328350
rect 128450 328294 128518 328350
rect 128574 328294 128642 328350
rect 128698 328294 128766 328350
rect 128822 328294 159114 328350
rect 159170 328294 159238 328350
rect 159294 328294 159362 328350
rect 159418 328294 159486 328350
rect 159542 328294 189834 328350
rect 189890 328294 189958 328350
rect 190014 328294 190082 328350
rect 190138 328294 190206 328350
rect 190262 328294 220554 328350
rect 220610 328294 220678 328350
rect 220734 328294 220802 328350
rect 220858 328294 220926 328350
rect 220982 328294 251274 328350
rect 251330 328294 251398 328350
rect 251454 328294 251522 328350
rect 251578 328294 251646 328350
rect 251702 328294 281994 328350
rect 282050 328294 282118 328350
rect 282174 328294 282242 328350
rect 282298 328294 282366 328350
rect 282422 328294 312714 328350
rect 312770 328294 312838 328350
rect 312894 328294 312962 328350
rect 313018 328294 313086 328350
rect 313142 328294 343434 328350
rect 343490 328294 343558 328350
rect 343614 328294 343682 328350
rect 343738 328294 343806 328350
rect 343862 328294 374154 328350
rect 374210 328294 374278 328350
rect 374334 328294 374402 328350
rect 374458 328294 374526 328350
rect 374582 328294 404874 328350
rect 404930 328294 404998 328350
rect 405054 328294 405122 328350
rect 405178 328294 405246 328350
rect 405302 328294 435594 328350
rect 435650 328294 435718 328350
rect 435774 328294 435842 328350
rect 435898 328294 435966 328350
rect 436022 328294 466314 328350
rect 466370 328294 466438 328350
rect 466494 328294 466562 328350
rect 466618 328294 466686 328350
rect 466742 328294 497034 328350
rect 497090 328294 497158 328350
rect 497214 328294 497282 328350
rect 497338 328294 497406 328350
rect 497462 328294 527754 328350
rect 527810 328294 527878 328350
rect 527934 328294 528002 328350
rect 528058 328294 528126 328350
rect 528182 328294 558474 328350
rect 558530 328294 558598 328350
rect 558654 328294 558722 328350
rect 558778 328294 558846 328350
rect 558902 328294 589194 328350
rect 589250 328294 589318 328350
rect 589374 328294 589442 328350
rect 589498 328294 589566 328350
rect 589622 328294 596496 328350
rect 596552 328294 596620 328350
rect 596676 328294 596744 328350
rect 596800 328294 596868 328350
rect 596924 328294 597980 328350
rect -1916 328226 597980 328294
rect -1916 328170 -860 328226
rect -804 328170 -736 328226
rect -680 328170 -612 328226
rect -556 328170 -488 328226
rect -432 328170 5514 328226
rect 5570 328170 5638 328226
rect 5694 328170 5762 328226
rect 5818 328170 5886 328226
rect 5942 328170 36234 328226
rect 36290 328170 36358 328226
rect 36414 328170 36482 328226
rect 36538 328170 36606 328226
rect 36662 328170 66954 328226
rect 67010 328170 67078 328226
rect 67134 328170 67202 328226
rect 67258 328170 67326 328226
rect 67382 328170 97674 328226
rect 97730 328170 97798 328226
rect 97854 328170 97922 328226
rect 97978 328170 98046 328226
rect 98102 328170 128394 328226
rect 128450 328170 128518 328226
rect 128574 328170 128642 328226
rect 128698 328170 128766 328226
rect 128822 328170 159114 328226
rect 159170 328170 159238 328226
rect 159294 328170 159362 328226
rect 159418 328170 159486 328226
rect 159542 328170 189834 328226
rect 189890 328170 189958 328226
rect 190014 328170 190082 328226
rect 190138 328170 190206 328226
rect 190262 328170 220554 328226
rect 220610 328170 220678 328226
rect 220734 328170 220802 328226
rect 220858 328170 220926 328226
rect 220982 328170 251274 328226
rect 251330 328170 251398 328226
rect 251454 328170 251522 328226
rect 251578 328170 251646 328226
rect 251702 328170 281994 328226
rect 282050 328170 282118 328226
rect 282174 328170 282242 328226
rect 282298 328170 282366 328226
rect 282422 328170 312714 328226
rect 312770 328170 312838 328226
rect 312894 328170 312962 328226
rect 313018 328170 313086 328226
rect 313142 328170 343434 328226
rect 343490 328170 343558 328226
rect 343614 328170 343682 328226
rect 343738 328170 343806 328226
rect 343862 328170 374154 328226
rect 374210 328170 374278 328226
rect 374334 328170 374402 328226
rect 374458 328170 374526 328226
rect 374582 328170 404874 328226
rect 404930 328170 404998 328226
rect 405054 328170 405122 328226
rect 405178 328170 405246 328226
rect 405302 328170 435594 328226
rect 435650 328170 435718 328226
rect 435774 328170 435842 328226
rect 435898 328170 435966 328226
rect 436022 328170 466314 328226
rect 466370 328170 466438 328226
rect 466494 328170 466562 328226
rect 466618 328170 466686 328226
rect 466742 328170 497034 328226
rect 497090 328170 497158 328226
rect 497214 328170 497282 328226
rect 497338 328170 497406 328226
rect 497462 328170 527754 328226
rect 527810 328170 527878 328226
rect 527934 328170 528002 328226
rect 528058 328170 528126 328226
rect 528182 328170 558474 328226
rect 558530 328170 558598 328226
rect 558654 328170 558722 328226
rect 558778 328170 558846 328226
rect 558902 328170 589194 328226
rect 589250 328170 589318 328226
rect 589374 328170 589442 328226
rect 589498 328170 589566 328226
rect 589622 328170 596496 328226
rect 596552 328170 596620 328226
rect 596676 328170 596744 328226
rect 596800 328170 596868 328226
rect 596924 328170 597980 328226
rect -1916 328102 597980 328170
rect -1916 328046 -860 328102
rect -804 328046 -736 328102
rect -680 328046 -612 328102
rect -556 328046 -488 328102
rect -432 328046 5514 328102
rect 5570 328046 5638 328102
rect 5694 328046 5762 328102
rect 5818 328046 5886 328102
rect 5942 328046 36234 328102
rect 36290 328046 36358 328102
rect 36414 328046 36482 328102
rect 36538 328046 36606 328102
rect 36662 328046 66954 328102
rect 67010 328046 67078 328102
rect 67134 328046 67202 328102
rect 67258 328046 67326 328102
rect 67382 328046 97674 328102
rect 97730 328046 97798 328102
rect 97854 328046 97922 328102
rect 97978 328046 98046 328102
rect 98102 328046 128394 328102
rect 128450 328046 128518 328102
rect 128574 328046 128642 328102
rect 128698 328046 128766 328102
rect 128822 328046 159114 328102
rect 159170 328046 159238 328102
rect 159294 328046 159362 328102
rect 159418 328046 159486 328102
rect 159542 328046 189834 328102
rect 189890 328046 189958 328102
rect 190014 328046 190082 328102
rect 190138 328046 190206 328102
rect 190262 328046 220554 328102
rect 220610 328046 220678 328102
rect 220734 328046 220802 328102
rect 220858 328046 220926 328102
rect 220982 328046 251274 328102
rect 251330 328046 251398 328102
rect 251454 328046 251522 328102
rect 251578 328046 251646 328102
rect 251702 328046 281994 328102
rect 282050 328046 282118 328102
rect 282174 328046 282242 328102
rect 282298 328046 282366 328102
rect 282422 328046 312714 328102
rect 312770 328046 312838 328102
rect 312894 328046 312962 328102
rect 313018 328046 313086 328102
rect 313142 328046 343434 328102
rect 343490 328046 343558 328102
rect 343614 328046 343682 328102
rect 343738 328046 343806 328102
rect 343862 328046 374154 328102
rect 374210 328046 374278 328102
rect 374334 328046 374402 328102
rect 374458 328046 374526 328102
rect 374582 328046 404874 328102
rect 404930 328046 404998 328102
rect 405054 328046 405122 328102
rect 405178 328046 405246 328102
rect 405302 328046 435594 328102
rect 435650 328046 435718 328102
rect 435774 328046 435842 328102
rect 435898 328046 435966 328102
rect 436022 328046 466314 328102
rect 466370 328046 466438 328102
rect 466494 328046 466562 328102
rect 466618 328046 466686 328102
rect 466742 328046 497034 328102
rect 497090 328046 497158 328102
rect 497214 328046 497282 328102
rect 497338 328046 497406 328102
rect 497462 328046 527754 328102
rect 527810 328046 527878 328102
rect 527934 328046 528002 328102
rect 528058 328046 528126 328102
rect 528182 328046 558474 328102
rect 558530 328046 558598 328102
rect 558654 328046 558722 328102
rect 558778 328046 558846 328102
rect 558902 328046 589194 328102
rect 589250 328046 589318 328102
rect 589374 328046 589442 328102
rect 589498 328046 589566 328102
rect 589622 328046 596496 328102
rect 596552 328046 596620 328102
rect 596676 328046 596744 328102
rect 596800 328046 596868 328102
rect 596924 328046 597980 328102
rect -1916 327978 597980 328046
rect -1916 327922 -860 327978
rect -804 327922 -736 327978
rect -680 327922 -612 327978
rect -556 327922 -488 327978
rect -432 327922 5514 327978
rect 5570 327922 5638 327978
rect 5694 327922 5762 327978
rect 5818 327922 5886 327978
rect 5942 327922 36234 327978
rect 36290 327922 36358 327978
rect 36414 327922 36482 327978
rect 36538 327922 36606 327978
rect 36662 327922 66954 327978
rect 67010 327922 67078 327978
rect 67134 327922 67202 327978
rect 67258 327922 67326 327978
rect 67382 327922 97674 327978
rect 97730 327922 97798 327978
rect 97854 327922 97922 327978
rect 97978 327922 98046 327978
rect 98102 327922 128394 327978
rect 128450 327922 128518 327978
rect 128574 327922 128642 327978
rect 128698 327922 128766 327978
rect 128822 327922 159114 327978
rect 159170 327922 159238 327978
rect 159294 327922 159362 327978
rect 159418 327922 159486 327978
rect 159542 327922 189834 327978
rect 189890 327922 189958 327978
rect 190014 327922 190082 327978
rect 190138 327922 190206 327978
rect 190262 327922 220554 327978
rect 220610 327922 220678 327978
rect 220734 327922 220802 327978
rect 220858 327922 220926 327978
rect 220982 327922 251274 327978
rect 251330 327922 251398 327978
rect 251454 327922 251522 327978
rect 251578 327922 251646 327978
rect 251702 327922 281994 327978
rect 282050 327922 282118 327978
rect 282174 327922 282242 327978
rect 282298 327922 282366 327978
rect 282422 327922 312714 327978
rect 312770 327922 312838 327978
rect 312894 327922 312962 327978
rect 313018 327922 313086 327978
rect 313142 327922 343434 327978
rect 343490 327922 343558 327978
rect 343614 327922 343682 327978
rect 343738 327922 343806 327978
rect 343862 327922 374154 327978
rect 374210 327922 374278 327978
rect 374334 327922 374402 327978
rect 374458 327922 374526 327978
rect 374582 327922 404874 327978
rect 404930 327922 404998 327978
rect 405054 327922 405122 327978
rect 405178 327922 405246 327978
rect 405302 327922 435594 327978
rect 435650 327922 435718 327978
rect 435774 327922 435842 327978
rect 435898 327922 435966 327978
rect 436022 327922 466314 327978
rect 466370 327922 466438 327978
rect 466494 327922 466562 327978
rect 466618 327922 466686 327978
rect 466742 327922 497034 327978
rect 497090 327922 497158 327978
rect 497214 327922 497282 327978
rect 497338 327922 497406 327978
rect 497462 327922 527754 327978
rect 527810 327922 527878 327978
rect 527934 327922 528002 327978
rect 528058 327922 528126 327978
rect 528182 327922 558474 327978
rect 558530 327922 558598 327978
rect 558654 327922 558722 327978
rect 558778 327922 558846 327978
rect 558902 327922 589194 327978
rect 589250 327922 589318 327978
rect 589374 327922 589442 327978
rect 589498 327922 589566 327978
rect 589622 327922 596496 327978
rect 596552 327922 596620 327978
rect 596676 327922 596744 327978
rect 596800 327922 596868 327978
rect 596924 327922 597980 327978
rect -1916 327826 597980 327922
rect -1916 316350 597980 316446
rect -1916 316294 -1820 316350
rect -1764 316294 -1696 316350
rect -1640 316294 -1572 316350
rect -1516 316294 -1448 316350
rect -1392 316294 9234 316350
rect 9290 316294 9358 316350
rect 9414 316294 9482 316350
rect 9538 316294 9606 316350
rect 9662 316294 39954 316350
rect 40010 316294 40078 316350
rect 40134 316294 40202 316350
rect 40258 316294 40326 316350
rect 40382 316294 70674 316350
rect 70730 316294 70798 316350
rect 70854 316294 70922 316350
rect 70978 316294 71046 316350
rect 71102 316294 101394 316350
rect 101450 316294 101518 316350
rect 101574 316294 101642 316350
rect 101698 316294 101766 316350
rect 101822 316294 132114 316350
rect 132170 316294 132238 316350
rect 132294 316294 132362 316350
rect 132418 316294 132486 316350
rect 132542 316294 162834 316350
rect 162890 316294 162958 316350
rect 163014 316294 163082 316350
rect 163138 316294 163206 316350
rect 163262 316294 193554 316350
rect 193610 316294 193678 316350
rect 193734 316294 193802 316350
rect 193858 316294 193926 316350
rect 193982 316294 224274 316350
rect 224330 316294 224398 316350
rect 224454 316294 224522 316350
rect 224578 316294 224646 316350
rect 224702 316294 254994 316350
rect 255050 316294 255118 316350
rect 255174 316294 255242 316350
rect 255298 316294 255366 316350
rect 255422 316294 285714 316350
rect 285770 316294 285838 316350
rect 285894 316294 285962 316350
rect 286018 316294 286086 316350
rect 286142 316294 316434 316350
rect 316490 316294 316558 316350
rect 316614 316294 316682 316350
rect 316738 316294 316806 316350
rect 316862 316294 347154 316350
rect 347210 316294 347278 316350
rect 347334 316294 347402 316350
rect 347458 316294 347526 316350
rect 347582 316294 377874 316350
rect 377930 316294 377998 316350
rect 378054 316294 378122 316350
rect 378178 316294 378246 316350
rect 378302 316294 408594 316350
rect 408650 316294 408718 316350
rect 408774 316294 408842 316350
rect 408898 316294 408966 316350
rect 409022 316294 439314 316350
rect 439370 316294 439438 316350
rect 439494 316294 439562 316350
rect 439618 316294 439686 316350
rect 439742 316294 470034 316350
rect 470090 316294 470158 316350
rect 470214 316294 470282 316350
rect 470338 316294 470406 316350
rect 470462 316294 500754 316350
rect 500810 316294 500878 316350
rect 500934 316294 501002 316350
rect 501058 316294 501126 316350
rect 501182 316294 531474 316350
rect 531530 316294 531598 316350
rect 531654 316294 531722 316350
rect 531778 316294 531846 316350
rect 531902 316294 562194 316350
rect 562250 316294 562318 316350
rect 562374 316294 562442 316350
rect 562498 316294 562566 316350
rect 562622 316294 592914 316350
rect 592970 316294 593038 316350
rect 593094 316294 593162 316350
rect 593218 316294 593286 316350
rect 593342 316294 597456 316350
rect 597512 316294 597580 316350
rect 597636 316294 597704 316350
rect 597760 316294 597828 316350
rect 597884 316294 597980 316350
rect -1916 316226 597980 316294
rect -1916 316170 -1820 316226
rect -1764 316170 -1696 316226
rect -1640 316170 -1572 316226
rect -1516 316170 -1448 316226
rect -1392 316170 9234 316226
rect 9290 316170 9358 316226
rect 9414 316170 9482 316226
rect 9538 316170 9606 316226
rect 9662 316170 39954 316226
rect 40010 316170 40078 316226
rect 40134 316170 40202 316226
rect 40258 316170 40326 316226
rect 40382 316170 70674 316226
rect 70730 316170 70798 316226
rect 70854 316170 70922 316226
rect 70978 316170 71046 316226
rect 71102 316170 101394 316226
rect 101450 316170 101518 316226
rect 101574 316170 101642 316226
rect 101698 316170 101766 316226
rect 101822 316170 132114 316226
rect 132170 316170 132238 316226
rect 132294 316170 132362 316226
rect 132418 316170 132486 316226
rect 132542 316170 162834 316226
rect 162890 316170 162958 316226
rect 163014 316170 163082 316226
rect 163138 316170 163206 316226
rect 163262 316170 193554 316226
rect 193610 316170 193678 316226
rect 193734 316170 193802 316226
rect 193858 316170 193926 316226
rect 193982 316170 224274 316226
rect 224330 316170 224398 316226
rect 224454 316170 224522 316226
rect 224578 316170 224646 316226
rect 224702 316170 254994 316226
rect 255050 316170 255118 316226
rect 255174 316170 255242 316226
rect 255298 316170 255366 316226
rect 255422 316170 285714 316226
rect 285770 316170 285838 316226
rect 285894 316170 285962 316226
rect 286018 316170 286086 316226
rect 286142 316170 316434 316226
rect 316490 316170 316558 316226
rect 316614 316170 316682 316226
rect 316738 316170 316806 316226
rect 316862 316170 347154 316226
rect 347210 316170 347278 316226
rect 347334 316170 347402 316226
rect 347458 316170 347526 316226
rect 347582 316170 377874 316226
rect 377930 316170 377998 316226
rect 378054 316170 378122 316226
rect 378178 316170 378246 316226
rect 378302 316170 408594 316226
rect 408650 316170 408718 316226
rect 408774 316170 408842 316226
rect 408898 316170 408966 316226
rect 409022 316170 439314 316226
rect 439370 316170 439438 316226
rect 439494 316170 439562 316226
rect 439618 316170 439686 316226
rect 439742 316170 470034 316226
rect 470090 316170 470158 316226
rect 470214 316170 470282 316226
rect 470338 316170 470406 316226
rect 470462 316170 500754 316226
rect 500810 316170 500878 316226
rect 500934 316170 501002 316226
rect 501058 316170 501126 316226
rect 501182 316170 531474 316226
rect 531530 316170 531598 316226
rect 531654 316170 531722 316226
rect 531778 316170 531846 316226
rect 531902 316170 562194 316226
rect 562250 316170 562318 316226
rect 562374 316170 562442 316226
rect 562498 316170 562566 316226
rect 562622 316170 592914 316226
rect 592970 316170 593038 316226
rect 593094 316170 593162 316226
rect 593218 316170 593286 316226
rect 593342 316170 597456 316226
rect 597512 316170 597580 316226
rect 597636 316170 597704 316226
rect 597760 316170 597828 316226
rect 597884 316170 597980 316226
rect -1916 316102 597980 316170
rect -1916 316046 -1820 316102
rect -1764 316046 -1696 316102
rect -1640 316046 -1572 316102
rect -1516 316046 -1448 316102
rect -1392 316046 9234 316102
rect 9290 316046 9358 316102
rect 9414 316046 9482 316102
rect 9538 316046 9606 316102
rect 9662 316046 39954 316102
rect 40010 316046 40078 316102
rect 40134 316046 40202 316102
rect 40258 316046 40326 316102
rect 40382 316046 70674 316102
rect 70730 316046 70798 316102
rect 70854 316046 70922 316102
rect 70978 316046 71046 316102
rect 71102 316046 101394 316102
rect 101450 316046 101518 316102
rect 101574 316046 101642 316102
rect 101698 316046 101766 316102
rect 101822 316046 132114 316102
rect 132170 316046 132238 316102
rect 132294 316046 132362 316102
rect 132418 316046 132486 316102
rect 132542 316046 162834 316102
rect 162890 316046 162958 316102
rect 163014 316046 163082 316102
rect 163138 316046 163206 316102
rect 163262 316046 193554 316102
rect 193610 316046 193678 316102
rect 193734 316046 193802 316102
rect 193858 316046 193926 316102
rect 193982 316046 224274 316102
rect 224330 316046 224398 316102
rect 224454 316046 224522 316102
rect 224578 316046 224646 316102
rect 224702 316046 254994 316102
rect 255050 316046 255118 316102
rect 255174 316046 255242 316102
rect 255298 316046 255366 316102
rect 255422 316046 285714 316102
rect 285770 316046 285838 316102
rect 285894 316046 285962 316102
rect 286018 316046 286086 316102
rect 286142 316046 316434 316102
rect 316490 316046 316558 316102
rect 316614 316046 316682 316102
rect 316738 316046 316806 316102
rect 316862 316046 347154 316102
rect 347210 316046 347278 316102
rect 347334 316046 347402 316102
rect 347458 316046 347526 316102
rect 347582 316046 377874 316102
rect 377930 316046 377998 316102
rect 378054 316046 378122 316102
rect 378178 316046 378246 316102
rect 378302 316046 408594 316102
rect 408650 316046 408718 316102
rect 408774 316046 408842 316102
rect 408898 316046 408966 316102
rect 409022 316046 439314 316102
rect 439370 316046 439438 316102
rect 439494 316046 439562 316102
rect 439618 316046 439686 316102
rect 439742 316046 470034 316102
rect 470090 316046 470158 316102
rect 470214 316046 470282 316102
rect 470338 316046 470406 316102
rect 470462 316046 500754 316102
rect 500810 316046 500878 316102
rect 500934 316046 501002 316102
rect 501058 316046 501126 316102
rect 501182 316046 531474 316102
rect 531530 316046 531598 316102
rect 531654 316046 531722 316102
rect 531778 316046 531846 316102
rect 531902 316046 562194 316102
rect 562250 316046 562318 316102
rect 562374 316046 562442 316102
rect 562498 316046 562566 316102
rect 562622 316046 592914 316102
rect 592970 316046 593038 316102
rect 593094 316046 593162 316102
rect 593218 316046 593286 316102
rect 593342 316046 597456 316102
rect 597512 316046 597580 316102
rect 597636 316046 597704 316102
rect 597760 316046 597828 316102
rect 597884 316046 597980 316102
rect -1916 315978 597980 316046
rect -1916 315922 -1820 315978
rect -1764 315922 -1696 315978
rect -1640 315922 -1572 315978
rect -1516 315922 -1448 315978
rect -1392 315922 9234 315978
rect 9290 315922 9358 315978
rect 9414 315922 9482 315978
rect 9538 315922 9606 315978
rect 9662 315922 39954 315978
rect 40010 315922 40078 315978
rect 40134 315922 40202 315978
rect 40258 315922 40326 315978
rect 40382 315922 70674 315978
rect 70730 315922 70798 315978
rect 70854 315922 70922 315978
rect 70978 315922 71046 315978
rect 71102 315922 101394 315978
rect 101450 315922 101518 315978
rect 101574 315922 101642 315978
rect 101698 315922 101766 315978
rect 101822 315922 132114 315978
rect 132170 315922 132238 315978
rect 132294 315922 132362 315978
rect 132418 315922 132486 315978
rect 132542 315922 162834 315978
rect 162890 315922 162958 315978
rect 163014 315922 163082 315978
rect 163138 315922 163206 315978
rect 163262 315922 193554 315978
rect 193610 315922 193678 315978
rect 193734 315922 193802 315978
rect 193858 315922 193926 315978
rect 193982 315922 224274 315978
rect 224330 315922 224398 315978
rect 224454 315922 224522 315978
rect 224578 315922 224646 315978
rect 224702 315922 254994 315978
rect 255050 315922 255118 315978
rect 255174 315922 255242 315978
rect 255298 315922 255366 315978
rect 255422 315922 285714 315978
rect 285770 315922 285838 315978
rect 285894 315922 285962 315978
rect 286018 315922 286086 315978
rect 286142 315922 316434 315978
rect 316490 315922 316558 315978
rect 316614 315922 316682 315978
rect 316738 315922 316806 315978
rect 316862 315922 347154 315978
rect 347210 315922 347278 315978
rect 347334 315922 347402 315978
rect 347458 315922 347526 315978
rect 347582 315922 377874 315978
rect 377930 315922 377998 315978
rect 378054 315922 378122 315978
rect 378178 315922 378246 315978
rect 378302 315922 408594 315978
rect 408650 315922 408718 315978
rect 408774 315922 408842 315978
rect 408898 315922 408966 315978
rect 409022 315922 439314 315978
rect 439370 315922 439438 315978
rect 439494 315922 439562 315978
rect 439618 315922 439686 315978
rect 439742 315922 470034 315978
rect 470090 315922 470158 315978
rect 470214 315922 470282 315978
rect 470338 315922 470406 315978
rect 470462 315922 500754 315978
rect 500810 315922 500878 315978
rect 500934 315922 501002 315978
rect 501058 315922 501126 315978
rect 501182 315922 531474 315978
rect 531530 315922 531598 315978
rect 531654 315922 531722 315978
rect 531778 315922 531846 315978
rect 531902 315922 562194 315978
rect 562250 315922 562318 315978
rect 562374 315922 562442 315978
rect 562498 315922 562566 315978
rect 562622 315922 592914 315978
rect 592970 315922 593038 315978
rect 593094 315922 593162 315978
rect 593218 315922 593286 315978
rect 593342 315922 597456 315978
rect 597512 315922 597580 315978
rect 597636 315922 597704 315978
rect 597760 315922 597828 315978
rect 597884 315922 597980 315978
rect -1916 315826 597980 315922
rect -1916 310350 597980 310446
rect -1916 310294 -860 310350
rect -804 310294 -736 310350
rect -680 310294 -612 310350
rect -556 310294 -488 310350
rect -432 310294 5514 310350
rect 5570 310294 5638 310350
rect 5694 310294 5762 310350
rect 5818 310294 5886 310350
rect 5942 310294 36234 310350
rect 36290 310294 36358 310350
rect 36414 310294 36482 310350
rect 36538 310294 36606 310350
rect 36662 310294 66954 310350
rect 67010 310294 67078 310350
rect 67134 310294 67202 310350
rect 67258 310294 67326 310350
rect 67382 310294 97674 310350
rect 97730 310294 97798 310350
rect 97854 310294 97922 310350
rect 97978 310294 98046 310350
rect 98102 310294 128394 310350
rect 128450 310294 128518 310350
rect 128574 310294 128642 310350
rect 128698 310294 128766 310350
rect 128822 310294 159114 310350
rect 159170 310294 159238 310350
rect 159294 310294 159362 310350
rect 159418 310294 159486 310350
rect 159542 310294 189834 310350
rect 189890 310294 189958 310350
rect 190014 310294 190082 310350
rect 190138 310294 190206 310350
rect 190262 310294 220554 310350
rect 220610 310294 220678 310350
rect 220734 310294 220802 310350
rect 220858 310294 220926 310350
rect 220982 310294 251274 310350
rect 251330 310294 251398 310350
rect 251454 310294 251522 310350
rect 251578 310294 251646 310350
rect 251702 310294 281994 310350
rect 282050 310294 282118 310350
rect 282174 310294 282242 310350
rect 282298 310294 282366 310350
rect 282422 310294 312714 310350
rect 312770 310294 312838 310350
rect 312894 310294 312962 310350
rect 313018 310294 313086 310350
rect 313142 310294 343434 310350
rect 343490 310294 343558 310350
rect 343614 310294 343682 310350
rect 343738 310294 343806 310350
rect 343862 310294 374154 310350
rect 374210 310294 374278 310350
rect 374334 310294 374402 310350
rect 374458 310294 374526 310350
rect 374582 310294 404874 310350
rect 404930 310294 404998 310350
rect 405054 310294 405122 310350
rect 405178 310294 405246 310350
rect 405302 310294 435594 310350
rect 435650 310294 435718 310350
rect 435774 310294 435842 310350
rect 435898 310294 435966 310350
rect 436022 310294 466314 310350
rect 466370 310294 466438 310350
rect 466494 310294 466562 310350
rect 466618 310294 466686 310350
rect 466742 310294 497034 310350
rect 497090 310294 497158 310350
rect 497214 310294 497282 310350
rect 497338 310294 497406 310350
rect 497462 310294 527754 310350
rect 527810 310294 527878 310350
rect 527934 310294 528002 310350
rect 528058 310294 528126 310350
rect 528182 310294 558474 310350
rect 558530 310294 558598 310350
rect 558654 310294 558722 310350
rect 558778 310294 558846 310350
rect 558902 310294 589194 310350
rect 589250 310294 589318 310350
rect 589374 310294 589442 310350
rect 589498 310294 589566 310350
rect 589622 310294 596496 310350
rect 596552 310294 596620 310350
rect 596676 310294 596744 310350
rect 596800 310294 596868 310350
rect 596924 310294 597980 310350
rect -1916 310226 597980 310294
rect -1916 310170 -860 310226
rect -804 310170 -736 310226
rect -680 310170 -612 310226
rect -556 310170 -488 310226
rect -432 310170 5514 310226
rect 5570 310170 5638 310226
rect 5694 310170 5762 310226
rect 5818 310170 5886 310226
rect 5942 310170 36234 310226
rect 36290 310170 36358 310226
rect 36414 310170 36482 310226
rect 36538 310170 36606 310226
rect 36662 310170 66954 310226
rect 67010 310170 67078 310226
rect 67134 310170 67202 310226
rect 67258 310170 67326 310226
rect 67382 310170 97674 310226
rect 97730 310170 97798 310226
rect 97854 310170 97922 310226
rect 97978 310170 98046 310226
rect 98102 310170 128394 310226
rect 128450 310170 128518 310226
rect 128574 310170 128642 310226
rect 128698 310170 128766 310226
rect 128822 310170 159114 310226
rect 159170 310170 159238 310226
rect 159294 310170 159362 310226
rect 159418 310170 159486 310226
rect 159542 310170 189834 310226
rect 189890 310170 189958 310226
rect 190014 310170 190082 310226
rect 190138 310170 190206 310226
rect 190262 310170 220554 310226
rect 220610 310170 220678 310226
rect 220734 310170 220802 310226
rect 220858 310170 220926 310226
rect 220982 310170 251274 310226
rect 251330 310170 251398 310226
rect 251454 310170 251522 310226
rect 251578 310170 251646 310226
rect 251702 310170 281994 310226
rect 282050 310170 282118 310226
rect 282174 310170 282242 310226
rect 282298 310170 282366 310226
rect 282422 310170 312714 310226
rect 312770 310170 312838 310226
rect 312894 310170 312962 310226
rect 313018 310170 313086 310226
rect 313142 310170 343434 310226
rect 343490 310170 343558 310226
rect 343614 310170 343682 310226
rect 343738 310170 343806 310226
rect 343862 310170 374154 310226
rect 374210 310170 374278 310226
rect 374334 310170 374402 310226
rect 374458 310170 374526 310226
rect 374582 310170 404874 310226
rect 404930 310170 404998 310226
rect 405054 310170 405122 310226
rect 405178 310170 405246 310226
rect 405302 310170 435594 310226
rect 435650 310170 435718 310226
rect 435774 310170 435842 310226
rect 435898 310170 435966 310226
rect 436022 310170 466314 310226
rect 466370 310170 466438 310226
rect 466494 310170 466562 310226
rect 466618 310170 466686 310226
rect 466742 310170 497034 310226
rect 497090 310170 497158 310226
rect 497214 310170 497282 310226
rect 497338 310170 497406 310226
rect 497462 310170 527754 310226
rect 527810 310170 527878 310226
rect 527934 310170 528002 310226
rect 528058 310170 528126 310226
rect 528182 310170 558474 310226
rect 558530 310170 558598 310226
rect 558654 310170 558722 310226
rect 558778 310170 558846 310226
rect 558902 310170 589194 310226
rect 589250 310170 589318 310226
rect 589374 310170 589442 310226
rect 589498 310170 589566 310226
rect 589622 310170 596496 310226
rect 596552 310170 596620 310226
rect 596676 310170 596744 310226
rect 596800 310170 596868 310226
rect 596924 310170 597980 310226
rect -1916 310102 597980 310170
rect -1916 310046 -860 310102
rect -804 310046 -736 310102
rect -680 310046 -612 310102
rect -556 310046 -488 310102
rect -432 310046 5514 310102
rect 5570 310046 5638 310102
rect 5694 310046 5762 310102
rect 5818 310046 5886 310102
rect 5942 310046 36234 310102
rect 36290 310046 36358 310102
rect 36414 310046 36482 310102
rect 36538 310046 36606 310102
rect 36662 310046 66954 310102
rect 67010 310046 67078 310102
rect 67134 310046 67202 310102
rect 67258 310046 67326 310102
rect 67382 310046 97674 310102
rect 97730 310046 97798 310102
rect 97854 310046 97922 310102
rect 97978 310046 98046 310102
rect 98102 310046 128394 310102
rect 128450 310046 128518 310102
rect 128574 310046 128642 310102
rect 128698 310046 128766 310102
rect 128822 310046 159114 310102
rect 159170 310046 159238 310102
rect 159294 310046 159362 310102
rect 159418 310046 159486 310102
rect 159542 310046 189834 310102
rect 189890 310046 189958 310102
rect 190014 310046 190082 310102
rect 190138 310046 190206 310102
rect 190262 310046 220554 310102
rect 220610 310046 220678 310102
rect 220734 310046 220802 310102
rect 220858 310046 220926 310102
rect 220982 310046 251274 310102
rect 251330 310046 251398 310102
rect 251454 310046 251522 310102
rect 251578 310046 251646 310102
rect 251702 310046 281994 310102
rect 282050 310046 282118 310102
rect 282174 310046 282242 310102
rect 282298 310046 282366 310102
rect 282422 310046 312714 310102
rect 312770 310046 312838 310102
rect 312894 310046 312962 310102
rect 313018 310046 313086 310102
rect 313142 310046 343434 310102
rect 343490 310046 343558 310102
rect 343614 310046 343682 310102
rect 343738 310046 343806 310102
rect 343862 310046 374154 310102
rect 374210 310046 374278 310102
rect 374334 310046 374402 310102
rect 374458 310046 374526 310102
rect 374582 310046 404874 310102
rect 404930 310046 404998 310102
rect 405054 310046 405122 310102
rect 405178 310046 405246 310102
rect 405302 310046 435594 310102
rect 435650 310046 435718 310102
rect 435774 310046 435842 310102
rect 435898 310046 435966 310102
rect 436022 310046 466314 310102
rect 466370 310046 466438 310102
rect 466494 310046 466562 310102
rect 466618 310046 466686 310102
rect 466742 310046 497034 310102
rect 497090 310046 497158 310102
rect 497214 310046 497282 310102
rect 497338 310046 497406 310102
rect 497462 310046 527754 310102
rect 527810 310046 527878 310102
rect 527934 310046 528002 310102
rect 528058 310046 528126 310102
rect 528182 310046 558474 310102
rect 558530 310046 558598 310102
rect 558654 310046 558722 310102
rect 558778 310046 558846 310102
rect 558902 310046 589194 310102
rect 589250 310046 589318 310102
rect 589374 310046 589442 310102
rect 589498 310046 589566 310102
rect 589622 310046 596496 310102
rect 596552 310046 596620 310102
rect 596676 310046 596744 310102
rect 596800 310046 596868 310102
rect 596924 310046 597980 310102
rect -1916 309978 597980 310046
rect -1916 309922 -860 309978
rect -804 309922 -736 309978
rect -680 309922 -612 309978
rect -556 309922 -488 309978
rect -432 309922 5514 309978
rect 5570 309922 5638 309978
rect 5694 309922 5762 309978
rect 5818 309922 5886 309978
rect 5942 309922 36234 309978
rect 36290 309922 36358 309978
rect 36414 309922 36482 309978
rect 36538 309922 36606 309978
rect 36662 309922 66954 309978
rect 67010 309922 67078 309978
rect 67134 309922 67202 309978
rect 67258 309922 67326 309978
rect 67382 309922 97674 309978
rect 97730 309922 97798 309978
rect 97854 309922 97922 309978
rect 97978 309922 98046 309978
rect 98102 309922 128394 309978
rect 128450 309922 128518 309978
rect 128574 309922 128642 309978
rect 128698 309922 128766 309978
rect 128822 309922 159114 309978
rect 159170 309922 159238 309978
rect 159294 309922 159362 309978
rect 159418 309922 159486 309978
rect 159542 309922 189834 309978
rect 189890 309922 189958 309978
rect 190014 309922 190082 309978
rect 190138 309922 190206 309978
rect 190262 309922 220554 309978
rect 220610 309922 220678 309978
rect 220734 309922 220802 309978
rect 220858 309922 220926 309978
rect 220982 309922 251274 309978
rect 251330 309922 251398 309978
rect 251454 309922 251522 309978
rect 251578 309922 251646 309978
rect 251702 309922 281994 309978
rect 282050 309922 282118 309978
rect 282174 309922 282242 309978
rect 282298 309922 282366 309978
rect 282422 309922 312714 309978
rect 312770 309922 312838 309978
rect 312894 309922 312962 309978
rect 313018 309922 313086 309978
rect 313142 309922 343434 309978
rect 343490 309922 343558 309978
rect 343614 309922 343682 309978
rect 343738 309922 343806 309978
rect 343862 309922 374154 309978
rect 374210 309922 374278 309978
rect 374334 309922 374402 309978
rect 374458 309922 374526 309978
rect 374582 309922 404874 309978
rect 404930 309922 404998 309978
rect 405054 309922 405122 309978
rect 405178 309922 405246 309978
rect 405302 309922 435594 309978
rect 435650 309922 435718 309978
rect 435774 309922 435842 309978
rect 435898 309922 435966 309978
rect 436022 309922 466314 309978
rect 466370 309922 466438 309978
rect 466494 309922 466562 309978
rect 466618 309922 466686 309978
rect 466742 309922 497034 309978
rect 497090 309922 497158 309978
rect 497214 309922 497282 309978
rect 497338 309922 497406 309978
rect 497462 309922 527754 309978
rect 527810 309922 527878 309978
rect 527934 309922 528002 309978
rect 528058 309922 528126 309978
rect 528182 309922 558474 309978
rect 558530 309922 558598 309978
rect 558654 309922 558722 309978
rect 558778 309922 558846 309978
rect 558902 309922 589194 309978
rect 589250 309922 589318 309978
rect 589374 309922 589442 309978
rect 589498 309922 589566 309978
rect 589622 309922 596496 309978
rect 596552 309922 596620 309978
rect 596676 309922 596744 309978
rect 596800 309922 596868 309978
rect 596924 309922 597980 309978
rect -1916 309826 597980 309922
rect -1916 298350 597980 298446
rect -1916 298294 -1820 298350
rect -1764 298294 -1696 298350
rect -1640 298294 -1572 298350
rect -1516 298294 -1448 298350
rect -1392 298294 9234 298350
rect 9290 298294 9358 298350
rect 9414 298294 9482 298350
rect 9538 298294 9606 298350
rect 9662 298294 39954 298350
rect 40010 298294 40078 298350
rect 40134 298294 40202 298350
rect 40258 298294 40326 298350
rect 40382 298294 70674 298350
rect 70730 298294 70798 298350
rect 70854 298294 70922 298350
rect 70978 298294 71046 298350
rect 71102 298294 101394 298350
rect 101450 298294 101518 298350
rect 101574 298294 101642 298350
rect 101698 298294 101766 298350
rect 101822 298294 132114 298350
rect 132170 298294 132238 298350
rect 132294 298294 132362 298350
rect 132418 298294 132486 298350
rect 132542 298294 162834 298350
rect 162890 298294 162958 298350
rect 163014 298294 163082 298350
rect 163138 298294 163206 298350
rect 163262 298294 193554 298350
rect 193610 298294 193678 298350
rect 193734 298294 193802 298350
rect 193858 298294 193926 298350
rect 193982 298294 224274 298350
rect 224330 298294 224398 298350
rect 224454 298294 224522 298350
rect 224578 298294 224646 298350
rect 224702 298294 254994 298350
rect 255050 298294 255118 298350
rect 255174 298294 255242 298350
rect 255298 298294 255366 298350
rect 255422 298294 285714 298350
rect 285770 298294 285838 298350
rect 285894 298294 285962 298350
rect 286018 298294 286086 298350
rect 286142 298294 316434 298350
rect 316490 298294 316558 298350
rect 316614 298294 316682 298350
rect 316738 298294 316806 298350
rect 316862 298294 347154 298350
rect 347210 298294 347278 298350
rect 347334 298294 347402 298350
rect 347458 298294 347526 298350
rect 347582 298294 377874 298350
rect 377930 298294 377998 298350
rect 378054 298294 378122 298350
rect 378178 298294 378246 298350
rect 378302 298294 408594 298350
rect 408650 298294 408718 298350
rect 408774 298294 408842 298350
rect 408898 298294 408966 298350
rect 409022 298294 439314 298350
rect 439370 298294 439438 298350
rect 439494 298294 439562 298350
rect 439618 298294 439686 298350
rect 439742 298294 470034 298350
rect 470090 298294 470158 298350
rect 470214 298294 470282 298350
rect 470338 298294 470406 298350
rect 470462 298294 500754 298350
rect 500810 298294 500878 298350
rect 500934 298294 501002 298350
rect 501058 298294 501126 298350
rect 501182 298294 531474 298350
rect 531530 298294 531598 298350
rect 531654 298294 531722 298350
rect 531778 298294 531846 298350
rect 531902 298294 562194 298350
rect 562250 298294 562318 298350
rect 562374 298294 562442 298350
rect 562498 298294 562566 298350
rect 562622 298294 592914 298350
rect 592970 298294 593038 298350
rect 593094 298294 593162 298350
rect 593218 298294 593286 298350
rect 593342 298294 597456 298350
rect 597512 298294 597580 298350
rect 597636 298294 597704 298350
rect 597760 298294 597828 298350
rect 597884 298294 597980 298350
rect -1916 298226 597980 298294
rect -1916 298170 -1820 298226
rect -1764 298170 -1696 298226
rect -1640 298170 -1572 298226
rect -1516 298170 -1448 298226
rect -1392 298170 9234 298226
rect 9290 298170 9358 298226
rect 9414 298170 9482 298226
rect 9538 298170 9606 298226
rect 9662 298170 39954 298226
rect 40010 298170 40078 298226
rect 40134 298170 40202 298226
rect 40258 298170 40326 298226
rect 40382 298170 70674 298226
rect 70730 298170 70798 298226
rect 70854 298170 70922 298226
rect 70978 298170 71046 298226
rect 71102 298170 101394 298226
rect 101450 298170 101518 298226
rect 101574 298170 101642 298226
rect 101698 298170 101766 298226
rect 101822 298170 132114 298226
rect 132170 298170 132238 298226
rect 132294 298170 132362 298226
rect 132418 298170 132486 298226
rect 132542 298170 162834 298226
rect 162890 298170 162958 298226
rect 163014 298170 163082 298226
rect 163138 298170 163206 298226
rect 163262 298170 193554 298226
rect 193610 298170 193678 298226
rect 193734 298170 193802 298226
rect 193858 298170 193926 298226
rect 193982 298170 224274 298226
rect 224330 298170 224398 298226
rect 224454 298170 224522 298226
rect 224578 298170 224646 298226
rect 224702 298170 254994 298226
rect 255050 298170 255118 298226
rect 255174 298170 255242 298226
rect 255298 298170 255366 298226
rect 255422 298170 285714 298226
rect 285770 298170 285838 298226
rect 285894 298170 285962 298226
rect 286018 298170 286086 298226
rect 286142 298170 316434 298226
rect 316490 298170 316558 298226
rect 316614 298170 316682 298226
rect 316738 298170 316806 298226
rect 316862 298170 347154 298226
rect 347210 298170 347278 298226
rect 347334 298170 347402 298226
rect 347458 298170 347526 298226
rect 347582 298170 377874 298226
rect 377930 298170 377998 298226
rect 378054 298170 378122 298226
rect 378178 298170 378246 298226
rect 378302 298170 408594 298226
rect 408650 298170 408718 298226
rect 408774 298170 408842 298226
rect 408898 298170 408966 298226
rect 409022 298170 439314 298226
rect 439370 298170 439438 298226
rect 439494 298170 439562 298226
rect 439618 298170 439686 298226
rect 439742 298170 470034 298226
rect 470090 298170 470158 298226
rect 470214 298170 470282 298226
rect 470338 298170 470406 298226
rect 470462 298170 500754 298226
rect 500810 298170 500878 298226
rect 500934 298170 501002 298226
rect 501058 298170 501126 298226
rect 501182 298170 531474 298226
rect 531530 298170 531598 298226
rect 531654 298170 531722 298226
rect 531778 298170 531846 298226
rect 531902 298170 562194 298226
rect 562250 298170 562318 298226
rect 562374 298170 562442 298226
rect 562498 298170 562566 298226
rect 562622 298170 592914 298226
rect 592970 298170 593038 298226
rect 593094 298170 593162 298226
rect 593218 298170 593286 298226
rect 593342 298170 597456 298226
rect 597512 298170 597580 298226
rect 597636 298170 597704 298226
rect 597760 298170 597828 298226
rect 597884 298170 597980 298226
rect -1916 298102 597980 298170
rect -1916 298046 -1820 298102
rect -1764 298046 -1696 298102
rect -1640 298046 -1572 298102
rect -1516 298046 -1448 298102
rect -1392 298046 9234 298102
rect 9290 298046 9358 298102
rect 9414 298046 9482 298102
rect 9538 298046 9606 298102
rect 9662 298046 39954 298102
rect 40010 298046 40078 298102
rect 40134 298046 40202 298102
rect 40258 298046 40326 298102
rect 40382 298046 70674 298102
rect 70730 298046 70798 298102
rect 70854 298046 70922 298102
rect 70978 298046 71046 298102
rect 71102 298046 101394 298102
rect 101450 298046 101518 298102
rect 101574 298046 101642 298102
rect 101698 298046 101766 298102
rect 101822 298046 132114 298102
rect 132170 298046 132238 298102
rect 132294 298046 132362 298102
rect 132418 298046 132486 298102
rect 132542 298046 162834 298102
rect 162890 298046 162958 298102
rect 163014 298046 163082 298102
rect 163138 298046 163206 298102
rect 163262 298046 193554 298102
rect 193610 298046 193678 298102
rect 193734 298046 193802 298102
rect 193858 298046 193926 298102
rect 193982 298046 224274 298102
rect 224330 298046 224398 298102
rect 224454 298046 224522 298102
rect 224578 298046 224646 298102
rect 224702 298046 254994 298102
rect 255050 298046 255118 298102
rect 255174 298046 255242 298102
rect 255298 298046 255366 298102
rect 255422 298046 285714 298102
rect 285770 298046 285838 298102
rect 285894 298046 285962 298102
rect 286018 298046 286086 298102
rect 286142 298046 316434 298102
rect 316490 298046 316558 298102
rect 316614 298046 316682 298102
rect 316738 298046 316806 298102
rect 316862 298046 347154 298102
rect 347210 298046 347278 298102
rect 347334 298046 347402 298102
rect 347458 298046 347526 298102
rect 347582 298046 377874 298102
rect 377930 298046 377998 298102
rect 378054 298046 378122 298102
rect 378178 298046 378246 298102
rect 378302 298046 408594 298102
rect 408650 298046 408718 298102
rect 408774 298046 408842 298102
rect 408898 298046 408966 298102
rect 409022 298046 439314 298102
rect 439370 298046 439438 298102
rect 439494 298046 439562 298102
rect 439618 298046 439686 298102
rect 439742 298046 470034 298102
rect 470090 298046 470158 298102
rect 470214 298046 470282 298102
rect 470338 298046 470406 298102
rect 470462 298046 500754 298102
rect 500810 298046 500878 298102
rect 500934 298046 501002 298102
rect 501058 298046 501126 298102
rect 501182 298046 531474 298102
rect 531530 298046 531598 298102
rect 531654 298046 531722 298102
rect 531778 298046 531846 298102
rect 531902 298046 562194 298102
rect 562250 298046 562318 298102
rect 562374 298046 562442 298102
rect 562498 298046 562566 298102
rect 562622 298046 592914 298102
rect 592970 298046 593038 298102
rect 593094 298046 593162 298102
rect 593218 298046 593286 298102
rect 593342 298046 597456 298102
rect 597512 298046 597580 298102
rect 597636 298046 597704 298102
rect 597760 298046 597828 298102
rect 597884 298046 597980 298102
rect -1916 297978 597980 298046
rect -1916 297922 -1820 297978
rect -1764 297922 -1696 297978
rect -1640 297922 -1572 297978
rect -1516 297922 -1448 297978
rect -1392 297922 9234 297978
rect 9290 297922 9358 297978
rect 9414 297922 9482 297978
rect 9538 297922 9606 297978
rect 9662 297922 39954 297978
rect 40010 297922 40078 297978
rect 40134 297922 40202 297978
rect 40258 297922 40326 297978
rect 40382 297922 70674 297978
rect 70730 297922 70798 297978
rect 70854 297922 70922 297978
rect 70978 297922 71046 297978
rect 71102 297922 101394 297978
rect 101450 297922 101518 297978
rect 101574 297922 101642 297978
rect 101698 297922 101766 297978
rect 101822 297922 132114 297978
rect 132170 297922 132238 297978
rect 132294 297922 132362 297978
rect 132418 297922 132486 297978
rect 132542 297922 162834 297978
rect 162890 297922 162958 297978
rect 163014 297922 163082 297978
rect 163138 297922 163206 297978
rect 163262 297922 193554 297978
rect 193610 297922 193678 297978
rect 193734 297922 193802 297978
rect 193858 297922 193926 297978
rect 193982 297922 224274 297978
rect 224330 297922 224398 297978
rect 224454 297922 224522 297978
rect 224578 297922 224646 297978
rect 224702 297922 254994 297978
rect 255050 297922 255118 297978
rect 255174 297922 255242 297978
rect 255298 297922 255366 297978
rect 255422 297922 285714 297978
rect 285770 297922 285838 297978
rect 285894 297922 285962 297978
rect 286018 297922 286086 297978
rect 286142 297922 316434 297978
rect 316490 297922 316558 297978
rect 316614 297922 316682 297978
rect 316738 297922 316806 297978
rect 316862 297922 347154 297978
rect 347210 297922 347278 297978
rect 347334 297922 347402 297978
rect 347458 297922 347526 297978
rect 347582 297922 377874 297978
rect 377930 297922 377998 297978
rect 378054 297922 378122 297978
rect 378178 297922 378246 297978
rect 378302 297922 408594 297978
rect 408650 297922 408718 297978
rect 408774 297922 408842 297978
rect 408898 297922 408966 297978
rect 409022 297922 439314 297978
rect 439370 297922 439438 297978
rect 439494 297922 439562 297978
rect 439618 297922 439686 297978
rect 439742 297922 470034 297978
rect 470090 297922 470158 297978
rect 470214 297922 470282 297978
rect 470338 297922 470406 297978
rect 470462 297922 500754 297978
rect 500810 297922 500878 297978
rect 500934 297922 501002 297978
rect 501058 297922 501126 297978
rect 501182 297922 531474 297978
rect 531530 297922 531598 297978
rect 531654 297922 531722 297978
rect 531778 297922 531846 297978
rect 531902 297922 562194 297978
rect 562250 297922 562318 297978
rect 562374 297922 562442 297978
rect 562498 297922 562566 297978
rect 562622 297922 592914 297978
rect 592970 297922 593038 297978
rect 593094 297922 593162 297978
rect 593218 297922 593286 297978
rect 593342 297922 597456 297978
rect 597512 297922 597580 297978
rect 597636 297922 597704 297978
rect 597760 297922 597828 297978
rect 597884 297922 597980 297978
rect -1916 297826 597980 297922
rect -1916 292350 597980 292446
rect -1916 292294 -860 292350
rect -804 292294 -736 292350
rect -680 292294 -612 292350
rect -556 292294 -488 292350
rect -432 292294 5514 292350
rect 5570 292294 5638 292350
rect 5694 292294 5762 292350
rect 5818 292294 5886 292350
rect 5942 292294 36234 292350
rect 36290 292294 36358 292350
rect 36414 292294 36482 292350
rect 36538 292294 36606 292350
rect 36662 292294 66954 292350
rect 67010 292294 67078 292350
rect 67134 292294 67202 292350
rect 67258 292294 67326 292350
rect 67382 292294 97674 292350
rect 97730 292294 97798 292350
rect 97854 292294 97922 292350
rect 97978 292294 98046 292350
rect 98102 292294 128394 292350
rect 128450 292294 128518 292350
rect 128574 292294 128642 292350
rect 128698 292294 128766 292350
rect 128822 292294 159114 292350
rect 159170 292294 159238 292350
rect 159294 292294 159362 292350
rect 159418 292294 159486 292350
rect 159542 292294 189834 292350
rect 189890 292294 189958 292350
rect 190014 292294 190082 292350
rect 190138 292294 190206 292350
rect 190262 292294 220554 292350
rect 220610 292294 220678 292350
rect 220734 292294 220802 292350
rect 220858 292294 220926 292350
rect 220982 292294 251274 292350
rect 251330 292294 251398 292350
rect 251454 292294 251522 292350
rect 251578 292294 251646 292350
rect 251702 292294 281994 292350
rect 282050 292294 282118 292350
rect 282174 292294 282242 292350
rect 282298 292294 282366 292350
rect 282422 292294 312714 292350
rect 312770 292294 312838 292350
rect 312894 292294 312962 292350
rect 313018 292294 313086 292350
rect 313142 292294 343434 292350
rect 343490 292294 343558 292350
rect 343614 292294 343682 292350
rect 343738 292294 343806 292350
rect 343862 292294 374154 292350
rect 374210 292294 374278 292350
rect 374334 292294 374402 292350
rect 374458 292294 374526 292350
rect 374582 292294 404874 292350
rect 404930 292294 404998 292350
rect 405054 292294 405122 292350
rect 405178 292294 405246 292350
rect 405302 292294 435594 292350
rect 435650 292294 435718 292350
rect 435774 292294 435842 292350
rect 435898 292294 435966 292350
rect 436022 292294 466314 292350
rect 466370 292294 466438 292350
rect 466494 292294 466562 292350
rect 466618 292294 466686 292350
rect 466742 292294 497034 292350
rect 497090 292294 497158 292350
rect 497214 292294 497282 292350
rect 497338 292294 497406 292350
rect 497462 292294 527754 292350
rect 527810 292294 527878 292350
rect 527934 292294 528002 292350
rect 528058 292294 528126 292350
rect 528182 292294 558474 292350
rect 558530 292294 558598 292350
rect 558654 292294 558722 292350
rect 558778 292294 558846 292350
rect 558902 292294 589194 292350
rect 589250 292294 589318 292350
rect 589374 292294 589442 292350
rect 589498 292294 589566 292350
rect 589622 292294 596496 292350
rect 596552 292294 596620 292350
rect 596676 292294 596744 292350
rect 596800 292294 596868 292350
rect 596924 292294 597980 292350
rect -1916 292226 597980 292294
rect -1916 292170 -860 292226
rect -804 292170 -736 292226
rect -680 292170 -612 292226
rect -556 292170 -488 292226
rect -432 292170 5514 292226
rect 5570 292170 5638 292226
rect 5694 292170 5762 292226
rect 5818 292170 5886 292226
rect 5942 292170 36234 292226
rect 36290 292170 36358 292226
rect 36414 292170 36482 292226
rect 36538 292170 36606 292226
rect 36662 292170 66954 292226
rect 67010 292170 67078 292226
rect 67134 292170 67202 292226
rect 67258 292170 67326 292226
rect 67382 292170 97674 292226
rect 97730 292170 97798 292226
rect 97854 292170 97922 292226
rect 97978 292170 98046 292226
rect 98102 292170 128394 292226
rect 128450 292170 128518 292226
rect 128574 292170 128642 292226
rect 128698 292170 128766 292226
rect 128822 292170 159114 292226
rect 159170 292170 159238 292226
rect 159294 292170 159362 292226
rect 159418 292170 159486 292226
rect 159542 292170 189834 292226
rect 189890 292170 189958 292226
rect 190014 292170 190082 292226
rect 190138 292170 190206 292226
rect 190262 292170 220554 292226
rect 220610 292170 220678 292226
rect 220734 292170 220802 292226
rect 220858 292170 220926 292226
rect 220982 292170 251274 292226
rect 251330 292170 251398 292226
rect 251454 292170 251522 292226
rect 251578 292170 251646 292226
rect 251702 292170 281994 292226
rect 282050 292170 282118 292226
rect 282174 292170 282242 292226
rect 282298 292170 282366 292226
rect 282422 292170 312714 292226
rect 312770 292170 312838 292226
rect 312894 292170 312962 292226
rect 313018 292170 313086 292226
rect 313142 292170 343434 292226
rect 343490 292170 343558 292226
rect 343614 292170 343682 292226
rect 343738 292170 343806 292226
rect 343862 292170 374154 292226
rect 374210 292170 374278 292226
rect 374334 292170 374402 292226
rect 374458 292170 374526 292226
rect 374582 292170 404874 292226
rect 404930 292170 404998 292226
rect 405054 292170 405122 292226
rect 405178 292170 405246 292226
rect 405302 292170 435594 292226
rect 435650 292170 435718 292226
rect 435774 292170 435842 292226
rect 435898 292170 435966 292226
rect 436022 292170 466314 292226
rect 466370 292170 466438 292226
rect 466494 292170 466562 292226
rect 466618 292170 466686 292226
rect 466742 292170 497034 292226
rect 497090 292170 497158 292226
rect 497214 292170 497282 292226
rect 497338 292170 497406 292226
rect 497462 292170 527754 292226
rect 527810 292170 527878 292226
rect 527934 292170 528002 292226
rect 528058 292170 528126 292226
rect 528182 292170 558474 292226
rect 558530 292170 558598 292226
rect 558654 292170 558722 292226
rect 558778 292170 558846 292226
rect 558902 292170 589194 292226
rect 589250 292170 589318 292226
rect 589374 292170 589442 292226
rect 589498 292170 589566 292226
rect 589622 292170 596496 292226
rect 596552 292170 596620 292226
rect 596676 292170 596744 292226
rect 596800 292170 596868 292226
rect 596924 292170 597980 292226
rect -1916 292102 597980 292170
rect -1916 292046 -860 292102
rect -804 292046 -736 292102
rect -680 292046 -612 292102
rect -556 292046 -488 292102
rect -432 292046 5514 292102
rect 5570 292046 5638 292102
rect 5694 292046 5762 292102
rect 5818 292046 5886 292102
rect 5942 292046 36234 292102
rect 36290 292046 36358 292102
rect 36414 292046 36482 292102
rect 36538 292046 36606 292102
rect 36662 292046 66954 292102
rect 67010 292046 67078 292102
rect 67134 292046 67202 292102
rect 67258 292046 67326 292102
rect 67382 292046 97674 292102
rect 97730 292046 97798 292102
rect 97854 292046 97922 292102
rect 97978 292046 98046 292102
rect 98102 292046 128394 292102
rect 128450 292046 128518 292102
rect 128574 292046 128642 292102
rect 128698 292046 128766 292102
rect 128822 292046 159114 292102
rect 159170 292046 159238 292102
rect 159294 292046 159362 292102
rect 159418 292046 159486 292102
rect 159542 292046 189834 292102
rect 189890 292046 189958 292102
rect 190014 292046 190082 292102
rect 190138 292046 190206 292102
rect 190262 292046 220554 292102
rect 220610 292046 220678 292102
rect 220734 292046 220802 292102
rect 220858 292046 220926 292102
rect 220982 292046 251274 292102
rect 251330 292046 251398 292102
rect 251454 292046 251522 292102
rect 251578 292046 251646 292102
rect 251702 292046 281994 292102
rect 282050 292046 282118 292102
rect 282174 292046 282242 292102
rect 282298 292046 282366 292102
rect 282422 292046 312714 292102
rect 312770 292046 312838 292102
rect 312894 292046 312962 292102
rect 313018 292046 313086 292102
rect 313142 292046 343434 292102
rect 343490 292046 343558 292102
rect 343614 292046 343682 292102
rect 343738 292046 343806 292102
rect 343862 292046 374154 292102
rect 374210 292046 374278 292102
rect 374334 292046 374402 292102
rect 374458 292046 374526 292102
rect 374582 292046 404874 292102
rect 404930 292046 404998 292102
rect 405054 292046 405122 292102
rect 405178 292046 405246 292102
rect 405302 292046 435594 292102
rect 435650 292046 435718 292102
rect 435774 292046 435842 292102
rect 435898 292046 435966 292102
rect 436022 292046 466314 292102
rect 466370 292046 466438 292102
rect 466494 292046 466562 292102
rect 466618 292046 466686 292102
rect 466742 292046 497034 292102
rect 497090 292046 497158 292102
rect 497214 292046 497282 292102
rect 497338 292046 497406 292102
rect 497462 292046 527754 292102
rect 527810 292046 527878 292102
rect 527934 292046 528002 292102
rect 528058 292046 528126 292102
rect 528182 292046 558474 292102
rect 558530 292046 558598 292102
rect 558654 292046 558722 292102
rect 558778 292046 558846 292102
rect 558902 292046 589194 292102
rect 589250 292046 589318 292102
rect 589374 292046 589442 292102
rect 589498 292046 589566 292102
rect 589622 292046 596496 292102
rect 596552 292046 596620 292102
rect 596676 292046 596744 292102
rect 596800 292046 596868 292102
rect 596924 292046 597980 292102
rect -1916 291978 597980 292046
rect -1916 291922 -860 291978
rect -804 291922 -736 291978
rect -680 291922 -612 291978
rect -556 291922 -488 291978
rect -432 291922 5514 291978
rect 5570 291922 5638 291978
rect 5694 291922 5762 291978
rect 5818 291922 5886 291978
rect 5942 291922 36234 291978
rect 36290 291922 36358 291978
rect 36414 291922 36482 291978
rect 36538 291922 36606 291978
rect 36662 291922 66954 291978
rect 67010 291922 67078 291978
rect 67134 291922 67202 291978
rect 67258 291922 67326 291978
rect 67382 291922 97674 291978
rect 97730 291922 97798 291978
rect 97854 291922 97922 291978
rect 97978 291922 98046 291978
rect 98102 291922 128394 291978
rect 128450 291922 128518 291978
rect 128574 291922 128642 291978
rect 128698 291922 128766 291978
rect 128822 291922 159114 291978
rect 159170 291922 159238 291978
rect 159294 291922 159362 291978
rect 159418 291922 159486 291978
rect 159542 291922 189834 291978
rect 189890 291922 189958 291978
rect 190014 291922 190082 291978
rect 190138 291922 190206 291978
rect 190262 291922 220554 291978
rect 220610 291922 220678 291978
rect 220734 291922 220802 291978
rect 220858 291922 220926 291978
rect 220982 291922 251274 291978
rect 251330 291922 251398 291978
rect 251454 291922 251522 291978
rect 251578 291922 251646 291978
rect 251702 291922 281994 291978
rect 282050 291922 282118 291978
rect 282174 291922 282242 291978
rect 282298 291922 282366 291978
rect 282422 291922 312714 291978
rect 312770 291922 312838 291978
rect 312894 291922 312962 291978
rect 313018 291922 313086 291978
rect 313142 291922 343434 291978
rect 343490 291922 343558 291978
rect 343614 291922 343682 291978
rect 343738 291922 343806 291978
rect 343862 291922 374154 291978
rect 374210 291922 374278 291978
rect 374334 291922 374402 291978
rect 374458 291922 374526 291978
rect 374582 291922 404874 291978
rect 404930 291922 404998 291978
rect 405054 291922 405122 291978
rect 405178 291922 405246 291978
rect 405302 291922 435594 291978
rect 435650 291922 435718 291978
rect 435774 291922 435842 291978
rect 435898 291922 435966 291978
rect 436022 291922 466314 291978
rect 466370 291922 466438 291978
rect 466494 291922 466562 291978
rect 466618 291922 466686 291978
rect 466742 291922 497034 291978
rect 497090 291922 497158 291978
rect 497214 291922 497282 291978
rect 497338 291922 497406 291978
rect 497462 291922 527754 291978
rect 527810 291922 527878 291978
rect 527934 291922 528002 291978
rect 528058 291922 528126 291978
rect 528182 291922 558474 291978
rect 558530 291922 558598 291978
rect 558654 291922 558722 291978
rect 558778 291922 558846 291978
rect 558902 291922 589194 291978
rect 589250 291922 589318 291978
rect 589374 291922 589442 291978
rect 589498 291922 589566 291978
rect 589622 291922 596496 291978
rect 596552 291922 596620 291978
rect 596676 291922 596744 291978
rect 596800 291922 596868 291978
rect 596924 291922 597980 291978
rect -1916 291826 597980 291922
rect -1916 280350 597980 280446
rect -1916 280294 -1820 280350
rect -1764 280294 -1696 280350
rect -1640 280294 -1572 280350
rect -1516 280294 -1448 280350
rect -1392 280294 9234 280350
rect 9290 280294 9358 280350
rect 9414 280294 9482 280350
rect 9538 280294 9606 280350
rect 9662 280294 39954 280350
rect 40010 280294 40078 280350
rect 40134 280294 40202 280350
rect 40258 280294 40326 280350
rect 40382 280294 70674 280350
rect 70730 280294 70798 280350
rect 70854 280294 70922 280350
rect 70978 280294 71046 280350
rect 71102 280294 101394 280350
rect 101450 280294 101518 280350
rect 101574 280294 101642 280350
rect 101698 280294 101766 280350
rect 101822 280294 132114 280350
rect 132170 280294 132238 280350
rect 132294 280294 132362 280350
rect 132418 280294 132486 280350
rect 132542 280294 162834 280350
rect 162890 280294 162958 280350
rect 163014 280294 163082 280350
rect 163138 280294 163206 280350
rect 163262 280294 193554 280350
rect 193610 280294 193678 280350
rect 193734 280294 193802 280350
rect 193858 280294 193926 280350
rect 193982 280294 224274 280350
rect 224330 280294 224398 280350
rect 224454 280294 224522 280350
rect 224578 280294 224646 280350
rect 224702 280294 254994 280350
rect 255050 280294 255118 280350
rect 255174 280294 255242 280350
rect 255298 280294 255366 280350
rect 255422 280294 285714 280350
rect 285770 280294 285838 280350
rect 285894 280294 285962 280350
rect 286018 280294 286086 280350
rect 286142 280294 316434 280350
rect 316490 280294 316558 280350
rect 316614 280294 316682 280350
rect 316738 280294 316806 280350
rect 316862 280294 347154 280350
rect 347210 280294 347278 280350
rect 347334 280294 347402 280350
rect 347458 280294 347526 280350
rect 347582 280294 377874 280350
rect 377930 280294 377998 280350
rect 378054 280294 378122 280350
rect 378178 280294 378246 280350
rect 378302 280294 408594 280350
rect 408650 280294 408718 280350
rect 408774 280294 408842 280350
rect 408898 280294 408966 280350
rect 409022 280294 439314 280350
rect 439370 280294 439438 280350
rect 439494 280294 439562 280350
rect 439618 280294 439686 280350
rect 439742 280294 470034 280350
rect 470090 280294 470158 280350
rect 470214 280294 470282 280350
rect 470338 280294 470406 280350
rect 470462 280294 500754 280350
rect 500810 280294 500878 280350
rect 500934 280294 501002 280350
rect 501058 280294 501126 280350
rect 501182 280294 531474 280350
rect 531530 280294 531598 280350
rect 531654 280294 531722 280350
rect 531778 280294 531846 280350
rect 531902 280294 562194 280350
rect 562250 280294 562318 280350
rect 562374 280294 562442 280350
rect 562498 280294 562566 280350
rect 562622 280294 592914 280350
rect 592970 280294 593038 280350
rect 593094 280294 593162 280350
rect 593218 280294 593286 280350
rect 593342 280294 597456 280350
rect 597512 280294 597580 280350
rect 597636 280294 597704 280350
rect 597760 280294 597828 280350
rect 597884 280294 597980 280350
rect -1916 280226 597980 280294
rect -1916 280170 -1820 280226
rect -1764 280170 -1696 280226
rect -1640 280170 -1572 280226
rect -1516 280170 -1448 280226
rect -1392 280170 9234 280226
rect 9290 280170 9358 280226
rect 9414 280170 9482 280226
rect 9538 280170 9606 280226
rect 9662 280170 39954 280226
rect 40010 280170 40078 280226
rect 40134 280170 40202 280226
rect 40258 280170 40326 280226
rect 40382 280170 70674 280226
rect 70730 280170 70798 280226
rect 70854 280170 70922 280226
rect 70978 280170 71046 280226
rect 71102 280170 101394 280226
rect 101450 280170 101518 280226
rect 101574 280170 101642 280226
rect 101698 280170 101766 280226
rect 101822 280170 132114 280226
rect 132170 280170 132238 280226
rect 132294 280170 132362 280226
rect 132418 280170 132486 280226
rect 132542 280170 162834 280226
rect 162890 280170 162958 280226
rect 163014 280170 163082 280226
rect 163138 280170 163206 280226
rect 163262 280170 193554 280226
rect 193610 280170 193678 280226
rect 193734 280170 193802 280226
rect 193858 280170 193926 280226
rect 193982 280170 224274 280226
rect 224330 280170 224398 280226
rect 224454 280170 224522 280226
rect 224578 280170 224646 280226
rect 224702 280170 254994 280226
rect 255050 280170 255118 280226
rect 255174 280170 255242 280226
rect 255298 280170 255366 280226
rect 255422 280170 285714 280226
rect 285770 280170 285838 280226
rect 285894 280170 285962 280226
rect 286018 280170 286086 280226
rect 286142 280170 316434 280226
rect 316490 280170 316558 280226
rect 316614 280170 316682 280226
rect 316738 280170 316806 280226
rect 316862 280170 347154 280226
rect 347210 280170 347278 280226
rect 347334 280170 347402 280226
rect 347458 280170 347526 280226
rect 347582 280170 377874 280226
rect 377930 280170 377998 280226
rect 378054 280170 378122 280226
rect 378178 280170 378246 280226
rect 378302 280170 408594 280226
rect 408650 280170 408718 280226
rect 408774 280170 408842 280226
rect 408898 280170 408966 280226
rect 409022 280170 439314 280226
rect 439370 280170 439438 280226
rect 439494 280170 439562 280226
rect 439618 280170 439686 280226
rect 439742 280170 470034 280226
rect 470090 280170 470158 280226
rect 470214 280170 470282 280226
rect 470338 280170 470406 280226
rect 470462 280170 500754 280226
rect 500810 280170 500878 280226
rect 500934 280170 501002 280226
rect 501058 280170 501126 280226
rect 501182 280170 531474 280226
rect 531530 280170 531598 280226
rect 531654 280170 531722 280226
rect 531778 280170 531846 280226
rect 531902 280170 562194 280226
rect 562250 280170 562318 280226
rect 562374 280170 562442 280226
rect 562498 280170 562566 280226
rect 562622 280170 592914 280226
rect 592970 280170 593038 280226
rect 593094 280170 593162 280226
rect 593218 280170 593286 280226
rect 593342 280170 597456 280226
rect 597512 280170 597580 280226
rect 597636 280170 597704 280226
rect 597760 280170 597828 280226
rect 597884 280170 597980 280226
rect -1916 280102 597980 280170
rect -1916 280046 -1820 280102
rect -1764 280046 -1696 280102
rect -1640 280046 -1572 280102
rect -1516 280046 -1448 280102
rect -1392 280046 9234 280102
rect 9290 280046 9358 280102
rect 9414 280046 9482 280102
rect 9538 280046 9606 280102
rect 9662 280046 39954 280102
rect 40010 280046 40078 280102
rect 40134 280046 40202 280102
rect 40258 280046 40326 280102
rect 40382 280046 70674 280102
rect 70730 280046 70798 280102
rect 70854 280046 70922 280102
rect 70978 280046 71046 280102
rect 71102 280046 101394 280102
rect 101450 280046 101518 280102
rect 101574 280046 101642 280102
rect 101698 280046 101766 280102
rect 101822 280046 132114 280102
rect 132170 280046 132238 280102
rect 132294 280046 132362 280102
rect 132418 280046 132486 280102
rect 132542 280046 162834 280102
rect 162890 280046 162958 280102
rect 163014 280046 163082 280102
rect 163138 280046 163206 280102
rect 163262 280046 193554 280102
rect 193610 280046 193678 280102
rect 193734 280046 193802 280102
rect 193858 280046 193926 280102
rect 193982 280046 224274 280102
rect 224330 280046 224398 280102
rect 224454 280046 224522 280102
rect 224578 280046 224646 280102
rect 224702 280046 254994 280102
rect 255050 280046 255118 280102
rect 255174 280046 255242 280102
rect 255298 280046 255366 280102
rect 255422 280046 285714 280102
rect 285770 280046 285838 280102
rect 285894 280046 285962 280102
rect 286018 280046 286086 280102
rect 286142 280046 316434 280102
rect 316490 280046 316558 280102
rect 316614 280046 316682 280102
rect 316738 280046 316806 280102
rect 316862 280046 347154 280102
rect 347210 280046 347278 280102
rect 347334 280046 347402 280102
rect 347458 280046 347526 280102
rect 347582 280046 377874 280102
rect 377930 280046 377998 280102
rect 378054 280046 378122 280102
rect 378178 280046 378246 280102
rect 378302 280046 408594 280102
rect 408650 280046 408718 280102
rect 408774 280046 408842 280102
rect 408898 280046 408966 280102
rect 409022 280046 439314 280102
rect 439370 280046 439438 280102
rect 439494 280046 439562 280102
rect 439618 280046 439686 280102
rect 439742 280046 470034 280102
rect 470090 280046 470158 280102
rect 470214 280046 470282 280102
rect 470338 280046 470406 280102
rect 470462 280046 500754 280102
rect 500810 280046 500878 280102
rect 500934 280046 501002 280102
rect 501058 280046 501126 280102
rect 501182 280046 531474 280102
rect 531530 280046 531598 280102
rect 531654 280046 531722 280102
rect 531778 280046 531846 280102
rect 531902 280046 562194 280102
rect 562250 280046 562318 280102
rect 562374 280046 562442 280102
rect 562498 280046 562566 280102
rect 562622 280046 592914 280102
rect 592970 280046 593038 280102
rect 593094 280046 593162 280102
rect 593218 280046 593286 280102
rect 593342 280046 597456 280102
rect 597512 280046 597580 280102
rect 597636 280046 597704 280102
rect 597760 280046 597828 280102
rect 597884 280046 597980 280102
rect -1916 279978 597980 280046
rect -1916 279922 -1820 279978
rect -1764 279922 -1696 279978
rect -1640 279922 -1572 279978
rect -1516 279922 -1448 279978
rect -1392 279922 9234 279978
rect 9290 279922 9358 279978
rect 9414 279922 9482 279978
rect 9538 279922 9606 279978
rect 9662 279922 39954 279978
rect 40010 279922 40078 279978
rect 40134 279922 40202 279978
rect 40258 279922 40326 279978
rect 40382 279922 70674 279978
rect 70730 279922 70798 279978
rect 70854 279922 70922 279978
rect 70978 279922 71046 279978
rect 71102 279922 101394 279978
rect 101450 279922 101518 279978
rect 101574 279922 101642 279978
rect 101698 279922 101766 279978
rect 101822 279922 132114 279978
rect 132170 279922 132238 279978
rect 132294 279922 132362 279978
rect 132418 279922 132486 279978
rect 132542 279922 162834 279978
rect 162890 279922 162958 279978
rect 163014 279922 163082 279978
rect 163138 279922 163206 279978
rect 163262 279922 193554 279978
rect 193610 279922 193678 279978
rect 193734 279922 193802 279978
rect 193858 279922 193926 279978
rect 193982 279922 224274 279978
rect 224330 279922 224398 279978
rect 224454 279922 224522 279978
rect 224578 279922 224646 279978
rect 224702 279922 254994 279978
rect 255050 279922 255118 279978
rect 255174 279922 255242 279978
rect 255298 279922 255366 279978
rect 255422 279922 285714 279978
rect 285770 279922 285838 279978
rect 285894 279922 285962 279978
rect 286018 279922 286086 279978
rect 286142 279922 316434 279978
rect 316490 279922 316558 279978
rect 316614 279922 316682 279978
rect 316738 279922 316806 279978
rect 316862 279922 347154 279978
rect 347210 279922 347278 279978
rect 347334 279922 347402 279978
rect 347458 279922 347526 279978
rect 347582 279922 377874 279978
rect 377930 279922 377998 279978
rect 378054 279922 378122 279978
rect 378178 279922 378246 279978
rect 378302 279922 408594 279978
rect 408650 279922 408718 279978
rect 408774 279922 408842 279978
rect 408898 279922 408966 279978
rect 409022 279922 439314 279978
rect 439370 279922 439438 279978
rect 439494 279922 439562 279978
rect 439618 279922 439686 279978
rect 439742 279922 470034 279978
rect 470090 279922 470158 279978
rect 470214 279922 470282 279978
rect 470338 279922 470406 279978
rect 470462 279922 500754 279978
rect 500810 279922 500878 279978
rect 500934 279922 501002 279978
rect 501058 279922 501126 279978
rect 501182 279922 531474 279978
rect 531530 279922 531598 279978
rect 531654 279922 531722 279978
rect 531778 279922 531846 279978
rect 531902 279922 562194 279978
rect 562250 279922 562318 279978
rect 562374 279922 562442 279978
rect 562498 279922 562566 279978
rect 562622 279922 592914 279978
rect 592970 279922 593038 279978
rect 593094 279922 593162 279978
rect 593218 279922 593286 279978
rect 593342 279922 597456 279978
rect 597512 279922 597580 279978
rect 597636 279922 597704 279978
rect 597760 279922 597828 279978
rect 597884 279922 597980 279978
rect -1916 279826 597980 279922
rect -1916 274350 597980 274446
rect -1916 274294 -860 274350
rect -804 274294 -736 274350
rect -680 274294 -612 274350
rect -556 274294 -488 274350
rect -432 274294 5514 274350
rect 5570 274294 5638 274350
rect 5694 274294 5762 274350
rect 5818 274294 5886 274350
rect 5942 274294 36234 274350
rect 36290 274294 36358 274350
rect 36414 274294 36482 274350
rect 36538 274294 36606 274350
rect 36662 274294 66954 274350
rect 67010 274294 67078 274350
rect 67134 274294 67202 274350
rect 67258 274294 67326 274350
rect 67382 274294 97674 274350
rect 97730 274294 97798 274350
rect 97854 274294 97922 274350
rect 97978 274294 98046 274350
rect 98102 274294 128394 274350
rect 128450 274294 128518 274350
rect 128574 274294 128642 274350
rect 128698 274294 128766 274350
rect 128822 274294 159114 274350
rect 159170 274294 159238 274350
rect 159294 274294 159362 274350
rect 159418 274294 159486 274350
rect 159542 274294 189834 274350
rect 189890 274294 189958 274350
rect 190014 274294 190082 274350
rect 190138 274294 190206 274350
rect 190262 274294 220554 274350
rect 220610 274294 220678 274350
rect 220734 274294 220802 274350
rect 220858 274294 220926 274350
rect 220982 274294 251274 274350
rect 251330 274294 251398 274350
rect 251454 274294 251522 274350
rect 251578 274294 251646 274350
rect 251702 274294 281994 274350
rect 282050 274294 282118 274350
rect 282174 274294 282242 274350
rect 282298 274294 282366 274350
rect 282422 274294 312714 274350
rect 312770 274294 312838 274350
rect 312894 274294 312962 274350
rect 313018 274294 313086 274350
rect 313142 274294 343434 274350
rect 343490 274294 343558 274350
rect 343614 274294 343682 274350
rect 343738 274294 343806 274350
rect 343862 274294 374154 274350
rect 374210 274294 374278 274350
rect 374334 274294 374402 274350
rect 374458 274294 374526 274350
rect 374582 274294 404874 274350
rect 404930 274294 404998 274350
rect 405054 274294 405122 274350
rect 405178 274294 405246 274350
rect 405302 274294 435594 274350
rect 435650 274294 435718 274350
rect 435774 274294 435842 274350
rect 435898 274294 435966 274350
rect 436022 274294 466314 274350
rect 466370 274294 466438 274350
rect 466494 274294 466562 274350
rect 466618 274294 466686 274350
rect 466742 274294 497034 274350
rect 497090 274294 497158 274350
rect 497214 274294 497282 274350
rect 497338 274294 497406 274350
rect 497462 274294 527754 274350
rect 527810 274294 527878 274350
rect 527934 274294 528002 274350
rect 528058 274294 528126 274350
rect 528182 274294 558474 274350
rect 558530 274294 558598 274350
rect 558654 274294 558722 274350
rect 558778 274294 558846 274350
rect 558902 274294 589194 274350
rect 589250 274294 589318 274350
rect 589374 274294 589442 274350
rect 589498 274294 589566 274350
rect 589622 274294 596496 274350
rect 596552 274294 596620 274350
rect 596676 274294 596744 274350
rect 596800 274294 596868 274350
rect 596924 274294 597980 274350
rect -1916 274226 597980 274294
rect -1916 274170 -860 274226
rect -804 274170 -736 274226
rect -680 274170 -612 274226
rect -556 274170 -488 274226
rect -432 274170 5514 274226
rect 5570 274170 5638 274226
rect 5694 274170 5762 274226
rect 5818 274170 5886 274226
rect 5942 274170 36234 274226
rect 36290 274170 36358 274226
rect 36414 274170 36482 274226
rect 36538 274170 36606 274226
rect 36662 274170 66954 274226
rect 67010 274170 67078 274226
rect 67134 274170 67202 274226
rect 67258 274170 67326 274226
rect 67382 274170 97674 274226
rect 97730 274170 97798 274226
rect 97854 274170 97922 274226
rect 97978 274170 98046 274226
rect 98102 274170 128394 274226
rect 128450 274170 128518 274226
rect 128574 274170 128642 274226
rect 128698 274170 128766 274226
rect 128822 274170 159114 274226
rect 159170 274170 159238 274226
rect 159294 274170 159362 274226
rect 159418 274170 159486 274226
rect 159542 274170 189834 274226
rect 189890 274170 189958 274226
rect 190014 274170 190082 274226
rect 190138 274170 190206 274226
rect 190262 274170 220554 274226
rect 220610 274170 220678 274226
rect 220734 274170 220802 274226
rect 220858 274170 220926 274226
rect 220982 274170 251274 274226
rect 251330 274170 251398 274226
rect 251454 274170 251522 274226
rect 251578 274170 251646 274226
rect 251702 274170 281994 274226
rect 282050 274170 282118 274226
rect 282174 274170 282242 274226
rect 282298 274170 282366 274226
rect 282422 274170 312714 274226
rect 312770 274170 312838 274226
rect 312894 274170 312962 274226
rect 313018 274170 313086 274226
rect 313142 274170 343434 274226
rect 343490 274170 343558 274226
rect 343614 274170 343682 274226
rect 343738 274170 343806 274226
rect 343862 274170 374154 274226
rect 374210 274170 374278 274226
rect 374334 274170 374402 274226
rect 374458 274170 374526 274226
rect 374582 274170 404874 274226
rect 404930 274170 404998 274226
rect 405054 274170 405122 274226
rect 405178 274170 405246 274226
rect 405302 274170 435594 274226
rect 435650 274170 435718 274226
rect 435774 274170 435842 274226
rect 435898 274170 435966 274226
rect 436022 274170 466314 274226
rect 466370 274170 466438 274226
rect 466494 274170 466562 274226
rect 466618 274170 466686 274226
rect 466742 274170 497034 274226
rect 497090 274170 497158 274226
rect 497214 274170 497282 274226
rect 497338 274170 497406 274226
rect 497462 274170 527754 274226
rect 527810 274170 527878 274226
rect 527934 274170 528002 274226
rect 528058 274170 528126 274226
rect 528182 274170 558474 274226
rect 558530 274170 558598 274226
rect 558654 274170 558722 274226
rect 558778 274170 558846 274226
rect 558902 274170 589194 274226
rect 589250 274170 589318 274226
rect 589374 274170 589442 274226
rect 589498 274170 589566 274226
rect 589622 274170 596496 274226
rect 596552 274170 596620 274226
rect 596676 274170 596744 274226
rect 596800 274170 596868 274226
rect 596924 274170 597980 274226
rect -1916 274102 597980 274170
rect -1916 274046 -860 274102
rect -804 274046 -736 274102
rect -680 274046 -612 274102
rect -556 274046 -488 274102
rect -432 274046 5514 274102
rect 5570 274046 5638 274102
rect 5694 274046 5762 274102
rect 5818 274046 5886 274102
rect 5942 274046 36234 274102
rect 36290 274046 36358 274102
rect 36414 274046 36482 274102
rect 36538 274046 36606 274102
rect 36662 274046 66954 274102
rect 67010 274046 67078 274102
rect 67134 274046 67202 274102
rect 67258 274046 67326 274102
rect 67382 274046 97674 274102
rect 97730 274046 97798 274102
rect 97854 274046 97922 274102
rect 97978 274046 98046 274102
rect 98102 274046 128394 274102
rect 128450 274046 128518 274102
rect 128574 274046 128642 274102
rect 128698 274046 128766 274102
rect 128822 274046 159114 274102
rect 159170 274046 159238 274102
rect 159294 274046 159362 274102
rect 159418 274046 159486 274102
rect 159542 274046 189834 274102
rect 189890 274046 189958 274102
rect 190014 274046 190082 274102
rect 190138 274046 190206 274102
rect 190262 274046 220554 274102
rect 220610 274046 220678 274102
rect 220734 274046 220802 274102
rect 220858 274046 220926 274102
rect 220982 274046 251274 274102
rect 251330 274046 251398 274102
rect 251454 274046 251522 274102
rect 251578 274046 251646 274102
rect 251702 274046 281994 274102
rect 282050 274046 282118 274102
rect 282174 274046 282242 274102
rect 282298 274046 282366 274102
rect 282422 274046 312714 274102
rect 312770 274046 312838 274102
rect 312894 274046 312962 274102
rect 313018 274046 313086 274102
rect 313142 274046 343434 274102
rect 343490 274046 343558 274102
rect 343614 274046 343682 274102
rect 343738 274046 343806 274102
rect 343862 274046 374154 274102
rect 374210 274046 374278 274102
rect 374334 274046 374402 274102
rect 374458 274046 374526 274102
rect 374582 274046 404874 274102
rect 404930 274046 404998 274102
rect 405054 274046 405122 274102
rect 405178 274046 405246 274102
rect 405302 274046 435594 274102
rect 435650 274046 435718 274102
rect 435774 274046 435842 274102
rect 435898 274046 435966 274102
rect 436022 274046 466314 274102
rect 466370 274046 466438 274102
rect 466494 274046 466562 274102
rect 466618 274046 466686 274102
rect 466742 274046 497034 274102
rect 497090 274046 497158 274102
rect 497214 274046 497282 274102
rect 497338 274046 497406 274102
rect 497462 274046 527754 274102
rect 527810 274046 527878 274102
rect 527934 274046 528002 274102
rect 528058 274046 528126 274102
rect 528182 274046 558474 274102
rect 558530 274046 558598 274102
rect 558654 274046 558722 274102
rect 558778 274046 558846 274102
rect 558902 274046 589194 274102
rect 589250 274046 589318 274102
rect 589374 274046 589442 274102
rect 589498 274046 589566 274102
rect 589622 274046 596496 274102
rect 596552 274046 596620 274102
rect 596676 274046 596744 274102
rect 596800 274046 596868 274102
rect 596924 274046 597980 274102
rect -1916 273978 597980 274046
rect -1916 273922 -860 273978
rect -804 273922 -736 273978
rect -680 273922 -612 273978
rect -556 273922 -488 273978
rect -432 273922 5514 273978
rect 5570 273922 5638 273978
rect 5694 273922 5762 273978
rect 5818 273922 5886 273978
rect 5942 273922 36234 273978
rect 36290 273922 36358 273978
rect 36414 273922 36482 273978
rect 36538 273922 36606 273978
rect 36662 273922 66954 273978
rect 67010 273922 67078 273978
rect 67134 273922 67202 273978
rect 67258 273922 67326 273978
rect 67382 273922 97674 273978
rect 97730 273922 97798 273978
rect 97854 273922 97922 273978
rect 97978 273922 98046 273978
rect 98102 273922 128394 273978
rect 128450 273922 128518 273978
rect 128574 273922 128642 273978
rect 128698 273922 128766 273978
rect 128822 273922 159114 273978
rect 159170 273922 159238 273978
rect 159294 273922 159362 273978
rect 159418 273922 159486 273978
rect 159542 273922 189834 273978
rect 189890 273922 189958 273978
rect 190014 273922 190082 273978
rect 190138 273922 190206 273978
rect 190262 273922 220554 273978
rect 220610 273922 220678 273978
rect 220734 273922 220802 273978
rect 220858 273922 220926 273978
rect 220982 273922 251274 273978
rect 251330 273922 251398 273978
rect 251454 273922 251522 273978
rect 251578 273922 251646 273978
rect 251702 273922 281994 273978
rect 282050 273922 282118 273978
rect 282174 273922 282242 273978
rect 282298 273922 282366 273978
rect 282422 273922 312714 273978
rect 312770 273922 312838 273978
rect 312894 273922 312962 273978
rect 313018 273922 313086 273978
rect 313142 273922 343434 273978
rect 343490 273922 343558 273978
rect 343614 273922 343682 273978
rect 343738 273922 343806 273978
rect 343862 273922 374154 273978
rect 374210 273922 374278 273978
rect 374334 273922 374402 273978
rect 374458 273922 374526 273978
rect 374582 273922 404874 273978
rect 404930 273922 404998 273978
rect 405054 273922 405122 273978
rect 405178 273922 405246 273978
rect 405302 273922 435594 273978
rect 435650 273922 435718 273978
rect 435774 273922 435842 273978
rect 435898 273922 435966 273978
rect 436022 273922 466314 273978
rect 466370 273922 466438 273978
rect 466494 273922 466562 273978
rect 466618 273922 466686 273978
rect 466742 273922 497034 273978
rect 497090 273922 497158 273978
rect 497214 273922 497282 273978
rect 497338 273922 497406 273978
rect 497462 273922 527754 273978
rect 527810 273922 527878 273978
rect 527934 273922 528002 273978
rect 528058 273922 528126 273978
rect 528182 273922 558474 273978
rect 558530 273922 558598 273978
rect 558654 273922 558722 273978
rect 558778 273922 558846 273978
rect 558902 273922 589194 273978
rect 589250 273922 589318 273978
rect 589374 273922 589442 273978
rect 589498 273922 589566 273978
rect 589622 273922 596496 273978
rect 596552 273922 596620 273978
rect 596676 273922 596744 273978
rect 596800 273922 596868 273978
rect 596924 273922 597980 273978
rect -1916 273826 597980 273922
rect -1916 262350 597980 262446
rect -1916 262294 -1820 262350
rect -1764 262294 -1696 262350
rect -1640 262294 -1572 262350
rect -1516 262294 -1448 262350
rect -1392 262294 9234 262350
rect 9290 262294 9358 262350
rect 9414 262294 9482 262350
rect 9538 262294 9606 262350
rect 9662 262294 39954 262350
rect 40010 262294 40078 262350
rect 40134 262294 40202 262350
rect 40258 262294 40326 262350
rect 40382 262294 70674 262350
rect 70730 262294 70798 262350
rect 70854 262294 70922 262350
rect 70978 262294 71046 262350
rect 71102 262294 101394 262350
rect 101450 262294 101518 262350
rect 101574 262294 101642 262350
rect 101698 262294 101766 262350
rect 101822 262294 132114 262350
rect 132170 262294 132238 262350
rect 132294 262294 132362 262350
rect 132418 262294 132486 262350
rect 132542 262294 162834 262350
rect 162890 262294 162958 262350
rect 163014 262294 163082 262350
rect 163138 262294 163206 262350
rect 163262 262294 193554 262350
rect 193610 262294 193678 262350
rect 193734 262294 193802 262350
rect 193858 262294 193926 262350
rect 193982 262294 224274 262350
rect 224330 262294 224398 262350
rect 224454 262294 224522 262350
rect 224578 262294 224646 262350
rect 224702 262294 254994 262350
rect 255050 262294 255118 262350
rect 255174 262294 255242 262350
rect 255298 262294 255366 262350
rect 255422 262294 285714 262350
rect 285770 262294 285838 262350
rect 285894 262294 285962 262350
rect 286018 262294 286086 262350
rect 286142 262294 316434 262350
rect 316490 262294 316558 262350
rect 316614 262294 316682 262350
rect 316738 262294 316806 262350
rect 316862 262294 347154 262350
rect 347210 262294 347278 262350
rect 347334 262294 347402 262350
rect 347458 262294 347526 262350
rect 347582 262294 377874 262350
rect 377930 262294 377998 262350
rect 378054 262294 378122 262350
rect 378178 262294 378246 262350
rect 378302 262294 408594 262350
rect 408650 262294 408718 262350
rect 408774 262294 408842 262350
rect 408898 262294 408966 262350
rect 409022 262294 439314 262350
rect 439370 262294 439438 262350
rect 439494 262294 439562 262350
rect 439618 262294 439686 262350
rect 439742 262294 470034 262350
rect 470090 262294 470158 262350
rect 470214 262294 470282 262350
rect 470338 262294 470406 262350
rect 470462 262294 500754 262350
rect 500810 262294 500878 262350
rect 500934 262294 501002 262350
rect 501058 262294 501126 262350
rect 501182 262294 531474 262350
rect 531530 262294 531598 262350
rect 531654 262294 531722 262350
rect 531778 262294 531846 262350
rect 531902 262294 562194 262350
rect 562250 262294 562318 262350
rect 562374 262294 562442 262350
rect 562498 262294 562566 262350
rect 562622 262294 592914 262350
rect 592970 262294 593038 262350
rect 593094 262294 593162 262350
rect 593218 262294 593286 262350
rect 593342 262294 597456 262350
rect 597512 262294 597580 262350
rect 597636 262294 597704 262350
rect 597760 262294 597828 262350
rect 597884 262294 597980 262350
rect -1916 262226 597980 262294
rect -1916 262170 -1820 262226
rect -1764 262170 -1696 262226
rect -1640 262170 -1572 262226
rect -1516 262170 -1448 262226
rect -1392 262170 9234 262226
rect 9290 262170 9358 262226
rect 9414 262170 9482 262226
rect 9538 262170 9606 262226
rect 9662 262170 39954 262226
rect 40010 262170 40078 262226
rect 40134 262170 40202 262226
rect 40258 262170 40326 262226
rect 40382 262170 70674 262226
rect 70730 262170 70798 262226
rect 70854 262170 70922 262226
rect 70978 262170 71046 262226
rect 71102 262170 101394 262226
rect 101450 262170 101518 262226
rect 101574 262170 101642 262226
rect 101698 262170 101766 262226
rect 101822 262170 132114 262226
rect 132170 262170 132238 262226
rect 132294 262170 132362 262226
rect 132418 262170 132486 262226
rect 132542 262170 162834 262226
rect 162890 262170 162958 262226
rect 163014 262170 163082 262226
rect 163138 262170 163206 262226
rect 163262 262170 193554 262226
rect 193610 262170 193678 262226
rect 193734 262170 193802 262226
rect 193858 262170 193926 262226
rect 193982 262170 224274 262226
rect 224330 262170 224398 262226
rect 224454 262170 224522 262226
rect 224578 262170 224646 262226
rect 224702 262170 254994 262226
rect 255050 262170 255118 262226
rect 255174 262170 255242 262226
rect 255298 262170 255366 262226
rect 255422 262170 285714 262226
rect 285770 262170 285838 262226
rect 285894 262170 285962 262226
rect 286018 262170 286086 262226
rect 286142 262170 316434 262226
rect 316490 262170 316558 262226
rect 316614 262170 316682 262226
rect 316738 262170 316806 262226
rect 316862 262170 347154 262226
rect 347210 262170 347278 262226
rect 347334 262170 347402 262226
rect 347458 262170 347526 262226
rect 347582 262170 377874 262226
rect 377930 262170 377998 262226
rect 378054 262170 378122 262226
rect 378178 262170 378246 262226
rect 378302 262170 408594 262226
rect 408650 262170 408718 262226
rect 408774 262170 408842 262226
rect 408898 262170 408966 262226
rect 409022 262170 439314 262226
rect 439370 262170 439438 262226
rect 439494 262170 439562 262226
rect 439618 262170 439686 262226
rect 439742 262170 470034 262226
rect 470090 262170 470158 262226
rect 470214 262170 470282 262226
rect 470338 262170 470406 262226
rect 470462 262170 500754 262226
rect 500810 262170 500878 262226
rect 500934 262170 501002 262226
rect 501058 262170 501126 262226
rect 501182 262170 531474 262226
rect 531530 262170 531598 262226
rect 531654 262170 531722 262226
rect 531778 262170 531846 262226
rect 531902 262170 562194 262226
rect 562250 262170 562318 262226
rect 562374 262170 562442 262226
rect 562498 262170 562566 262226
rect 562622 262170 592914 262226
rect 592970 262170 593038 262226
rect 593094 262170 593162 262226
rect 593218 262170 593286 262226
rect 593342 262170 597456 262226
rect 597512 262170 597580 262226
rect 597636 262170 597704 262226
rect 597760 262170 597828 262226
rect 597884 262170 597980 262226
rect -1916 262102 597980 262170
rect -1916 262046 -1820 262102
rect -1764 262046 -1696 262102
rect -1640 262046 -1572 262102
rect -1516 262046 -1448 262102
rect -1392 262046 9234 262102
rect 9290 262046 9358 262102
rect 9414 262046 9482 262102
rect 9538 262046 9606 262102
rect 9662 262046 39954 262102
rect 40010 262046 40078 262102
rect 40134 262046 40202 262102
rect 40258 262046 40326 262102
rect 40382 262046 70674 262102
rect 70730 262046 70798 262102
rect 70854 262046 70922 262102
rect 70978 262046 71046 262102
rect 71102 262046 101394 262102
rect 101450 262046 101518 262102
rect 101574 262046 101642 262102
rect 101698 262046 101766 262102
rect 101822 262046 132114 262102
rect 132170 262046 132238 262102
rect 132294 262046 132362 262102
rect 132418 262046 132486 262102
rect 132542 262046 162834 262102
rect 162890 262046 162958 262102
rect 163014 262046 163082 262102
rect 163138 262046 163206 262102
rect 163262 262046 193554 262102
rect 193610 262046 193678 262102
rect 193734 262046 193802 262102
rect 193858 262046 193926 262102
rect 193982 262046 224274 262102
rect 224330 262046 224398 262102
rect 224454 262046 224522 262102
rect 224578 262046 224646 262102
rect 224702 262046 254994 262102
rect 255050 262046 255118 262102
rect 255174 262046 255242 262102
rect 255298 262046 255366 262102
rect 255422 262046 285714 262102
rect 285770 262046 285838 262102
rect 285894 262046 285962 262102
rect 286018 262046 286086 262102
rect 286142 262046 316434 262102
rect 316490 262046 316558 262102
rect 316614 262046 316682 262102
rect 316738 262046 316806 262102
rect 316862 262046 347154 262102
rect 347210 262046 347278 262102
rect 347334 262046 347402 262102
rect 347458 262046 347526 262102
rect 347582 262046 377874 262102
rect 377930 262046 377998 262102
rect 378054 262046 378122 262102
rect 378178 262046 378246 262102
rect 378302 262046 408594 262102
rect 408650 262046 408718 262102
rect 408774 262046 408842 262102
rect 408898 262046 408966 262102
rect 409022 262046 439314 262102
rect 439370 262046 439438 262102
rect 439494 262046 439562 262102
rect 439618 262046 439686 262102
rect 439742 262046 470034 262102
rect 470090 262046 470158 262102
rect 470214 262046 470282 262102
rect 470338 262046 470406 262102
rect 470462 262046 500754 262102
rect 500810 262046 500878 262102
rect 500934 262046 501002 262102
rect 501058 262046 501126 262102
rect 501182 262046 531474 262102
rect 531530 262046 531598 262102
rect 531654 262046 531722 262102
rect 531778 262046 531846 262102
rect 531902 262046 562194 262102
rect 562250 262046 562318 262102
rect 562374 262046 562442 262102
rect 562498 262046 562566 262102
rect 562622 262046 592914 262102
rect 592970 262046 593038 262102
rect 593094 262046 593162 262102
rect 593218 262046 593286 262102
rect 593342 262046 597456 262102
rect 597512 262046 597580 262102
rect 597636 262046 597704 262102
rect 597760 262046 597828 262102
rect 597884 262046 597980 262102
rect -1916 261978 597980 262046
rect -1916 261922 -1820 261978
rect -1764 261922 -1696 261978
rect -1640 261922 -1572 261978
rect -1516 261922 -1448 261978
rect -1392 261922 9234 261978
rect 9290 261922 9358 261978
rect 9414 261922 9482 261978
rect 9538 261922 9606 261978
rect 9662 261922 39954 261978
rect 40010 261922 40078 261978
rect 40134 261922 40202 261978
rect 40258 261922 40326 261978
rect 40382 261922 70674 261978
rect 70730 261922 70798 261978
rect 70854 261922 70922 261978
rect 70978 261922 71046 261978
rect 71102 261922 101394 261978
rect 101450 261922 101518 261978
rect 101574 261922 101642 261978
rect 101698 261922 101766 261978
rect 101822 261922 132114 261978
rect 132170 261922 132238 261978
rect 132294 261922 132362 261978
rect 132418 261922 132486 261978
rect 132542 261922 162834 261978
rect 162890 261922 162958 261978
rect 163014 261922 163082 261978
rect 163138 261922 163206 261978
rect 163262 261922 193554 261978
rect 193610 261922 193678 261978
rect 193734 261922 193802 261978
rect 193858 261922 193926 261978
rect 193982 261922 224274 261978
rect 224330 261922 224398 261978
rect 224454 261922 224522 261978
rect 224578 261922 224646 261978
rect 224702 261922 254994 261978
rect 255050 261922 255118 261978
rect 255174 261922 255242 261978
rect 255298 261922 255366 261978
rect 255422 261922 285714 261978
rect 285770 261922 285838 261978
rect 285894 261922 285962 261978
rect 286018 261922 286086 261978
rect 286142 261922 316434 261978
rect 316490 261922 316558 261978
rect 316614 261922 316682 261978
rect 316738 261922 316806 261978
rect 316862 261922 347154 261978
rect 347210 261922 347278 261978
rect 347334 261922 347402 261978
rect 347458 261922 347526 261978
rect 347582 261922 377874 261978
rect 377930 261922 377998 261978
rect 378054 261922 378122 261978
rect 378178 261922 378246 261978
rect 378302 261922 408594 261978
rect 408650 261922 408718 261978
rect 408774 261922 408842 261978
rect 408898 261922 408966 261978
rect 409022 261922 439314 261978
rect 439370 261922 439438 261978
rect 439494 261922 439562 261978
rect 439618 261922 439686 261978
rect 439742 261922 470034 261978
rect 470090 261922 470158 261978
rect 470214 261922 470282 261978
rect 470338 261922 470406 261978
rect 470462 261922 500754 261978
rect 500810 261922 500878 261978
rect 500934 261922 501002 261978
rect 501058 261922 501126 261978
rect 501182 261922 531474 261978
rect 531530 261922 531598 261978
rect 531654 261922 531722 261978
rect 531778 261922 531846 261978
rect 531902 261922 562194 261978
rect 562250 261922 562318 261978
rect 562374 261922 562442 261978
rect 562498 261922 562566 261978
rect 562622 261922 592914 261978
rect 592970 261922 593038 261978
rect 593094 261922 593162 261978
rect 593218 261922 593286 261978
rect 593342 261922 597456 261978
rect 597512 261922 597580 261978
rect 597636 261922 597704 261978
rect 597760 261922 597828 261978
rect 597884 261922 597980 261978
rect -1916 261826 597980 261922
rect -1916 256350 597980 256446
rect -1916 256294 -860 256350
rect -804 256294 -736 256350
rect -680 256294 -612 256350
rect -556 256294 -488 256350
rect -432 256294 5514 256350
rect 5570 256294 5638 256350
rect 5694 256294 5762 256350
rect 5818 256294 5886 256350
rect 5942 256294 36234 256350
rect 36290 256294 36358 256350
rect 36414 256294 36482 256350
rect 36538 256294 36606 256350
rect 36662 256294 66954 256350
rect 67010 256294 67078 256350
rect 67134 256294 67202 256350
rect 67258 256294 67326 256350
rect 67382 256294 97674 256350
rect 97730 256294 97798 256350
rect 97854 256294 97922 256350
rect 97978 256294 98046 256350
rect 98102 256294 128394 256350
rect 128450 256294 128518 256350
rect 128574 256294 128642 256350
rect 128698 256294 128766 256350
rect 128822 256294 159114 256350
rect 159170 256294 159238 256350
rect 159294 256294 159362 256350
rect 159418 256294 159486 256350
rect 159542 256294 189834 256350
rect 189890 256294 189958 256350
rect 190014 256294 190082 256350
rect 190138 256294 190206 256350
rect 190262 256294 220554 256350
rect 220610 256294 220678 256350
rect 220734 256294 220802 256350
rect 220858 256294 220926 256350
rect 220982 256294 251274 256350
rect 251330 256294 251398 256350
rect 251454 256294 251522 256350
rect 251578 256294 251646 256350
rect 251702 256294 281994 256350
rect 282050 256294 282118 256350
rect 282174 256294 282242 256350
rect 282298 256294 282366 256350
rect 282422 256294 312714 256350
rect 312770 256294 312838 256350
rect 312894 256294 312962 256350
rect 313018 256294 313086 256350
rect 313142 256294 343434 256350
rect 343490 256294 343558 256350
rect 343614 256294 343682 256350
rect 343738 256294 343806 256350
rect 343862 256294 374154 256350
rect 374210 256294 374278 256350
rect 374334 256294 374402 256350
rect 374458 256294 374526 256350
rect 374582 256294 404874 256350
rect 404930 256294 404998 256350
rect 405054 256294 405122 256350
rect 405178 256294 405246 256350
rect 405302 256294 435594 256350
rect 435650 256294 435718 256350
rect 435774 256294 435842 256350
rect 435898 256294 435966 256350
rect 436022 256294 466314 256350
rect 466370 256294 466438 256350
rect 466494 256294 466562 256350
rect 466618 256294 466686 256350
rect 466742 256294 497034 256350
rect 497090 256294 497158 256350
rect 497214 256294 497282 256350
rect 497338 256294 497406 256350
rect 497462 256294 527754 256350
rect 527810 256294 527878 256350
rect 527934 256294 528002 256350
rect 528058 256294 528126 256350
rect 528182 256294 558474 256350
rect 558530 256294 558598 256350
rect 558654 256294 558722 256350
rect 558778 256294 558846 256350
rect 558902 256294 589194 256350
rect 589250 256294 589318 256350
rect 589374 256294 589442 256350
rect 589498 256294 589566 256350
rect 589622 256294 596496 256350
rect 596552 256294 596620 256350
rect 596676 256294 596744 256350
rect 596800 256294 596868 256350
rect 596924 256294 597980 256350
rect -1916 256226 597980 256294
rect -1916 256170 -860 256226
rect -804 256170 -736 256226
rect -680 256170 -612 256226
rect -556 256170 -488 256226
rect -432 256170 5514 256226
rect 5570 256170 5638 256226
rect 5694 256170 5762 256226
rect 5818 256170 5886 256226
rect 5942 256170 36234 256226
rect 36290 256170 36358 256226
rect 36414 256170 36482 256226
rect 36538 256170 36606 256226
rect 36662 256170 66954 256226
rect 67010 256170 67078 256226
rect 67134 256170 67202 256226
rect 67258 256170 67326 256226
rect 67382 256170 97674 256226
rect 97730 256170 97798 256226
rect 97854 256170 97922 256226
rect 97978 256170 98046 256226
rect 98102 256170 128394 256226
rect 128450 256170 128518 256226
rect 128574 256170 128642 256226
rect 128698 256170 128766 256226
rect 128822 256170 159114 256226
rect 159170 256170 159238 256226
rect 159294 256170 159362 256226
rect 159418 256170 159486 256226
rect 159542 256170 189834 256226
rect 189890 256170 189958 256226
rect 190014 256170 190082 256226
rect 190138 256170 190206 256226
rect 190262 256170 220554 256226
rect 220610 256170 220678 256226
rect 220734 256170 220802 256226
rect 220858 256170 220926 256226
rect 220982 256170 251274 256226
rect 251330 256170 251398 256226
rect 251454 256170 251522 256226
rect 251578 256170 251646 256226
rect 251702 256170 281994 256226
rect 282050 256170 282118 256226
rect 282174 256170 282242 256226
rect 282298 256170 282366 256226
rect 282422 256170 312714 256226
rect 312770 256170 312838 256226
rect 312894 256170 312962 256226
rect 313018 256170 313086 256226
rect 313142 256170 343434 256226
rect 343490 256170 343558 256226
rect 343614 256170 343682 256226
rect 343738 256170 343806 256226
rect 343862 256170 374154 256226
rect 374210 256170 374278 256226
rect 374334 256170 374402 256226
rect 374458 256170 374526 256226
rect 374582 256170 404874 256226
rect 404930 256170 404998 256226
rect 405054 256170 405122 256226
rect 405178 256170 405246 256226
rect 405302 256170 435594 256226
rect 435650 256170 435718 256226
rect 435774 256170 435842 256226
rect 435898 256170 435966 256226
rect 436022 256170 466314 256226
rect 466370 256170 466438 256226
rect 466494 256170 466562 256226
rect 466618 256170 466686 256226
rect 466742 256170 497034 256226
rect 497090 256170 497158 256226
rect 497214 256170 497282 256226
rect 497338 256170 497406 256226
rect 497462 256170 527754 256226
rect 527810 256170 527878 256226
rect 527934 256170 528002 256226
rect 528058 256170 528126 256226
rect 528182 256170 558474 256226
rect 558530 256170 558598 256226
rect 558654 256170 558722 256226
rect 558778 256170 558846 256226
rect 558902 256170 589194 256226
rect 589250 256170 589318 256226
rect 589374 256170 589442 256226
rect 589498 256170 589566 256226
rect 589622 256170 596496 256226
rect 596552 256170 596620 256226
rect 596676 256170 596744 256226
rect 596800 256170 596868 256226
rect 596924 256170 597980 256226
rect -1916 256102 597980 256170
rect -1916 256046 -860 256102
rect -804 256046 -736 256102
rect -680 256046 -612 256102
rect -556 256046 -488 256102
rect -432 256046 5514 256102
rect 5570 256046 5638 256102
rect 5694 256046 5762 256102
rect 5818 256046 5886 256102
rect 5942 256046 36234 256102
rect 36290 256046 36358 256102
rect 36414 256046 36482 256102
rect 36538 256046 36606 256102
rect 36662 256046 66954 256102
rect 67010 256046 67078 256102
rect 67134 256046 67202 256102
rect 67258 256046 67326 256102
rect 67382 256046 97674 256102
rect 97730 256046 97798 256102
rect 97854 256046 97922 256102
rect 97978 256046 98046 256102
rect 98102 256046 128394 256102
rect 128450 256046 128518 256102
rect 128574 256046 128642 256102
rect 128698 256046 128766 256102
rect 128822 256046 159114 256102
rect 159170 256046 159238 256102
rect 159294 256046 159362 256102
rect 159418 256046 159486 256102
rect 159542 256046 189834 256102
rect 189890 256046 189958 256102
rect 190014 256046 190082 256102
rect 190138 256046 190206 256102
rect 190262 256046 220554 256102
rect 220610 256046 220678 256102
rect 220734 256046 220802 256102
rect 220858 256046 220926 256102
rect 220982 256046 251274 256102
rect 251330 256046 251398 256102
rect 251454 256046 251522 256102
rect 251578 256046 251646 256102
rect 251702 256046 281994 256102
rect 282050 256046 282118 256102
rect 282174 256046 282242 256102
rect 282298 256046 282366 256102
rect 282422 256046 312714 256102
rect 312770 256046 312838 256102
rect 312894 256046 312962 256102
rect 313018 256046 313086 256102
rect 313142 256046 343434 256102
rect 343490 256046 343558 256102
rect 343614 256046 343682 256102
rect 343738 256046 343806 256102
rect 343862 256046 374154 256102
rect 374210 256046 374278 256102
rect 374334 256046 374402 256102
rect 374458 256046 374526 256102
rect 374582 256046 404874 256102
rect 404930 256046 404998 256102
rect 405054 256046 405122 256102
rect 405178 256046 405246 256102
rect 405302 256046 435594 256102
rect 435650 256046 435718 256102
rect 435774 256046 435842 256102
rect 435898 256046 435966 256102
rect 436022 256046 466314 256102
rect 466370 256046 466438 256102
rect 466494 256046 466562 256102
rect 466618 256046 466686 256102
rect 466742 256046 497034 256102
rect 497090 256046 497158 256102
rect 497214 256046 497282 256102
rect 497338 256046 497406 256102
rect 497462 256046 527754 256102
rect 527810 256046 527878 256102
rect 527934 256046 528002 256102
rect 528058 256046 528126 256102
rect 528182 256046 558474 256102
rect 558530 256046 558598 256102
rect 558654 256046 558722 256102
rect 558778 256046 558846 256102
rect 558902 256046 589194 256102
rect 589250 256046 589318 256102
rect 589374 256046 589442 256102
rect 589498 256046 589566 256102
rect 589622 256046 596496 256102
rect 596552 256046 596620 256102
rect 596676 256046 596744 256102
rect 596800 256046 596868 256102
rect 596924 256046 597980 256102
rect -1916 255978 597980 256046
rect -1916 255922 -860 255978
rect -804 255922 -736 255978
rect -680 255922 -612 255978
rect -556 255922 -488 255978
rect -432 255922 5514 255978
rect 5570 255922 5638 255978
rect 5694 255922 5762 255978
rect 5818 255922 5886 255978
rect 5942 255922 36234 255978
rect 36290 255922 36358 255978
rect 36414 255922 36482 255978
rect 36538 255922 36606 255978
rect 36662 255922 66954 255978
rect 67010 255922 67078 255978
rect 67134 255922 67202 255978
rect 67258 255922 67326 255978
rect 67382 255922 97674 255978
rect 97730 255922 97798 255978
rect 97854 255922 97922 255978
rect 97978 255922 98046 255978
rect 98102 255922 128394 255978
rect 128450 255922 128518 255978
rect 128574 255922 128642 255978
rect 128698 255922 128766 255978
rect 128822 255922 159114 255978
rect 159170 255922 159238 255978
rect 159294 255922 159362 255978
rect 159418 255922 159486 255978
rect 159542 255922 189834 255978
rect 189890 255922 189958 255978
rect 190014 255922 190082 255978
rect 190138 255922 190206 255978
rect 190262 255922 220554 255978
rect 220610 255922 220678 255978
rect 220734 255922 220802 255978
rect 220858 255922 220926 255978
rect 220982 255922 251274 255978
rect 251330 255922 251398 255978
rect 251454 255922 251522 255978
rect 251578 255922 251646 255978
rect 251702 255922 281994 255978
rect 282050 255922 282118 255978
rect 282174 255922 282242 255978
rect 282298 255922 282366 255978
rect 282422 255922 312714 255978
rect 312770 255922 312838 255978
rect 312894 255922 312962 255978
rect 313018 255922 313086 255978
rect 313142 255922 343434 255978
rect 343490 255922 343558 255978
rect 343614 255922 343682 255978
rect 343738 255922 343806 255978
rect 343862 255922 374154 255978
rect 374210 255922 374278 255978
rect 374334 255922 374402 255978
rect 374458 255922 374526 255978
rect 374582 255922 404874 255978
rect 404930 255922 404998 255978
rect 405054 255922 405122 255978
rect 405178 255922 405246 255978
rect 405302 255922 435594 255978
rect 435650 255922 435718 255978
rect 435774 255922 435842 255978
rect 435898 255922 435966 255978
rect 436022 255922 466314 255978
rect 466370 255922 466438 255978
rect 466494 255922 466562 255978
rect 466618 255922 466686 255978
rect 466742 255922 497034 255978
rect 497090 255922 497158 255978
rect 497214 255922 497282 255978
rect 497338 255922 497406 255978
rect 497462 255922 527754 255978
rect 527810 255922 527878 255978
rect 527934 255922 528002 255978
rect 528058 255922 528126 255978
rect 528182 255922 558474 255978
rect 558530 255922 558598 255978
rect 558654 255922 558722 255978
rect 558778 255922 558846 255978
rect 558902 255922 589194 255978
rect 589250 255922 589318 255978
rect 589374 255922 589442 255978
rect 589498 255922 589566 255978
rect 589622 255922 596496 255978
rect 596552 255922 596620 255978
rect 596676 255922 596744 255978
rect 596800 255922 596868 255978
rect 596924 255922 597980 255978
rect -1916 255826 597980 255922
rect -1916 244350 597980 244446
rect -1916 244294 -1820 244350
rect -1764 244294 -1696 244350
rect -1640 244294 -1572 244350
rect -1516 244294 -1448 244350
rect -1392 244294 9234 244350
rect 9290 244294 9358 244350
rect 9414 244294 9482 244350
rect 9538 244294 9606 244350
rect 9662 244294 39954 244350
rect 40010 244294 40078 244350
rect 40134 244294 40202 244350
rect 40258 244294 40326 244350
rect 40382 244294 70674 244350
rect 70730 244294 70798 244350
rect 70854 244294 70922 244350
rect 70978 244294 71046 244350
rect 71102 244294 101394 244350
rect 101450 244294 101518 244350
rect 101574 244294 101642 244350
rect 101698 244294 101766 244350
rect 101822 244294 132114 244350
rect 132170 244294 132238 244350
rect 132294 244294 132362 244350
rect 132418 244294 132486 244350
rect 132542 244294 162834 244350
rect 162890 244294 162958 244350
rect 163014 244294 163082 244350
rect 163138 244294 163206 244350
rect 163262 244294 193554 244350
rect 193610 244294 193678 244350
rect 193734 244294 193802 244350
rect 193858 244294 193926 244350
rect 193982 244294 224274 244350
rect 224330 244294 224398 244350
rect 224454 244294 224522 244350
rect 224578 244294 224646 244350
rect 224702 244294 254994 244350
rect 255050 244294 255118 244350
rect 255174 244294 255242 244350
rect 255298 244294 255366 244350
rect 255422 244294 285714 244350
rect 285770 244294 285838 244350
rect 285894 244294 285962 244350
rect 286018 244294 286086 244350
rect 286142 244294 316434 244350
rect 316490 244294 316558 244350
rect 316614 244294 316682 244350
rect 316738 244294 316806 244350
rect 316862 244294 347154 244350
rect 347210 244294 347278 244350
rect 347334 244294 347402 244350
rect 347458 244294 347526 244350
rect 347582 244294 377874 244350
rect 377930 244294 377998 244350
rect 378054 244294 378122 244350
rect 378178 244294 378246 244350
rect 378302 244294 408594 244350
rect 408650 244294 408718 244350
rect 408774 244294 408842 244350
rect 408898 244294 408966 244350
rect 409022 244294 439314 244350
rect 439370 244294 439438 244350
rect 439494 244294 439562 244350
rect 439618 244294 439686 244350
rect 439742 244294 470034 244350
rect 470090 244294 470158 244350
rect 470214 244294 470282 244350
rect 470338 244294 470406 244350
rect 470462 244294 500754 244350
rect 500810 244294 500878 244350
rect 500934 244294 501002 244350
rect 501058 244294 501126 244350
rect 501182 244294 531474 244350
rect 531530 244294 531598 244350
rect 531654 244294 531722 244350
rect 531778 244294 531846 244350
rect 531902 244294 562194 244350
rect 562250 244294 562318 244350
rect 562374 244294 562442 244350
rect 562498 244294 562566 244350
rect 562622 244294 592914 244350
rect 592970 244294 593038 244350
rect 593094 244294 593162 244350
rect 593218 244294 593286 244350
rect 593342 244294 597456 244350
rect 597512 244294 597580 244350
rect 597636 244294 597704 244350
rect 597760 244294 597828 244350
rect 597884 244294 597980 244350
rect -1916 244226 597980 244294
rect -1916 244170 -1820 244226
rect -1764 244170 -1696 244226
rect -1640 244170 -1572 244226
rect -1516 244170 -1448 244226
rect -1392 244170 9234 244226
rect 9290 244170 9358 244226
rect 9414 244170 9482 244226
rect 9538 244170 9606 244226
rect 9662 244170 39954 244226
rect 40010 244170 40078 244226
rect 40134 244170 40202 244226
rect 40258 244170 40326 244226
rect 40382 244170 70674 244226
rect 70730 244170 70798 244226
rect 70854 244170 70922 244226
rect 70978 244170 71046 244226
rect 71102 244170 101394 244226
rect 101450 244170 101518 244226
rect 101574 244170 101642 244226
rect 101698 244170 101766 244226
rect 101822 244170 132114 244226
rect 132170 244170 132238 244226
rect 132294 244170 132362 244226
rect 132418 244170 132486 244226
rect 132542 244170 162834 244226
rect 162890 244170 162958 244226
rect 163014 244170 163082 244226
rect 163138 244170 163206 244226
rect 163262 244170 193554 244226
rect 193610 244170 193678 244226
rect 193734 244170 193802 244226
rect 193858 244170 193926 244226
rect 193982 244170 224274 244226
rect 224330 244170 224398 244226
rect 224454 244170 224522 244226
rect 224578 244170 224646 244226
rect 224702 244170 254994 244226
rect 255050 244170 255118 244226
rect 255174 244170 255242 244226
rect 255298 244170 255366 244226
rect 255422 244170 285714 244226
rect 285770 244170 285838 244226
rect 285894 244170 285962 244226
rect 286018 244170 286086 244226
rect 286142 244170 316434 244226
rect 316490 244170 316558 244226
rect 316614 244170 316682 244226
rect 316738 244170 316806 244226
rect 316862 244170 347154 244226
rect 347210 244170 347278 244226
rect 347334 244170 347402 244226
rect 347458 244170 347526 244226
rect 347582 244170 377874 244226
rect 377930 244170 377998 244226
rect 378054 244170 378122 244226
rect 378178 244170 378246 244226
rect 378302 244170 408594 244226
rect 408650 244170 408718 244226
rect 408774 244170 408842 244226
rect 408898 244170 408966 244226
rect 409022 244170 439314 244226
rect 439370 244170 439438 244226
rect 439494 244170 439562 244226
rect 439618 244170 439686 244226
rect 439742 244170 470034 244226
rect 470090 244170 470158 244226
rect 470214 244170 470282 244226
rect 470338 244170 470406 244226
rect 470462 244170 500754 244226
rect 500810 244170 500878 244226
rect 500934 244170 501002 244226
rect 501058 244170 501126 244226
rect 501182 244170 531474 244226
rect 531530 244170 531598 244226
rect 531654 244170 531722 244226
rect 531778 244170 531846 244226
rect 531902 244170 562194 244226
rect 562250 244170 562318 244226
rect 562374 244170 562442 244226
rect 562498 244170 562566 244226
rect 562622 244170 592914 244226
rect 592970 244170 593038 244226
rect 593094 244170 593162 244226
rect 593218 244170 593286 244226
rect 593342 244170 597456 244226
rect 597512 244170 597580 244226
rect 597636 244170 597704 244226
rect 597760 244170 597828 244226
rect 597884 244170 597980 244226
rect -1916 244102 597980 244170
rect -1916 244046 -1820 244102
rect -1764 244046 -1696 244102
rect -1640 244046 -1572 244102
rect -1516 244046 -1448 244102
rect -1392 244046 9234 244102
rect 9290 244046 9358 244102
rect 9414 244046 9482 244102
rect 9538 244046 9606 244102
rect 9662 244046 39954 244102
rect 40010 244046 40078 244102
rect 40134 244046 40202 244102
rect 40258 244046 40326 244102
rect 40382 244046 70674 244102
rect 70730 244046 70798 244102
rect 70854 244046 70922 244102
rect 70978 244046 71046 244102
rect 71102 244046 101394 244102
rect 101450 244046 101518 244102
rect 101574 244046 101642 244102
rect 101698 244046 101766 244102
rect 101822 244046 132114 244102
rect 132170 244046 132238 244102
rect 132294 244046 132362 244102
rect 132418 244046 132486 244102
rect 132542 244046 162834 244102
rect 162890 244046 162958 244102
rect 163014 244046 163082 244102
rect 163138 244046 163206 244102
rect 163262 244046 193554 244102
rect 193610 244046 193678 244102
rect 193734 244046 193802 244102
rect 193858 244046 193926 244102
rect 193982 244046 224274 244102
rect 224330 244046 224398 244102
rect 224454 244046 224522 244102
rect 224578 244046 224646 244102
rect 224702 244046 254994 244102
rect 255050 244046 255118 244102
rect 255174 244046 255242 244102
rect 255298 244046 255366 244102
rect 255422 244046 285714 244102
rect 285770 244046 285838 244102
rect 285894 244046 285962 244102
rect 286018 244046 286086 244102
rect 286142 244046 316434 244102
rect 316490 244046 316558 244102
rect 316614 244046 316682 244102
rect 316738 244046 316806 244102
rect 316862 244046 347154 244102
rect 347210 244046 347278 244102
rect 347334 244046 347402 244102
rect 347458 244046 347526 244102
rect 347582 244046 377874 244102
rect 377930 244046 377998 244102
rect 378054 244046 378122 244102
rect 378178 244046 378246 244102
rect 378302 244046 408594 244102
rect 408650 244046 408718 244102
rect 408774 244046 408842 244102
rect 408898 244046 408966 244102
rect 409022 244046 439314 244102
rect 439370 244046 439438 244102
rect 439494 244046 439562 244102
rect 439618 244046 439686 244102
rect 439742 244046 470034 244102
rect 470090 244046 470158 244102
rect 470214 244046 470282 244102
rect 470338 244046 470406 244102
rect 470462 244046 500754 244102
rect 500810 244046 500878 244102
rect 500934 244046 501002 244102
rect 501058 244046 501126 244102
rect 501182 244046 531474 244102
rect 531530 244046 531598 244102
rect 531654 244046 531722 244102
rect 531778 244046 531846 244102
rect 531902 244046 562194 244102
rect 562250 244046 562318 244102
rect 562374 244046 562442 244102
rect 562498 244046 562566 244102
rect 562622 244046 592914 244102
rect 592970 244046 593038 244102
rect 593094 244046 593162 244102
rect 593218 244046 593286 244102
rect 593342 244046 597456 244102
rect 597512 244046 597580 244102
rect 597636 244046 597704 244102
rect 597760 244046 597828 244102
rect 597884 244046 597980 244102
rect -1916 243978 597980 244046
rect -1916 243922 -1820 243978
rect -1764 243922 -1696 243978
rect -1640 243922 -1572 243978
rect -1516 243922 -1448 243978
rect -1392 243922 9234 243978
rect 9290 243922 9358 243978
rect 9414 243922 9482 243978
rect 9538 243922 9606 243978
rect 9662 243922 39954 243978
rect 40010 243922 40078 243978
rect 40134 243922 40202 243978
rect 40258 243922 40326 243978
rect 40382 243922 70674 243978
rect 70730 243922 70798 243978
rect 70854 243922 70922 243978
rect 70978 243922 71046 243978
rect 71102 243922 101394 243978
rect 101450 243922 101518 243978
rect 101574 243922 101642 243978
rect 101698 243922 101766 243978
rect 101822 243922 132114 243978
rect 132170 243922 132238 243978
rect 132294 243922 132362 243978
rect 132418 243922 132486 243978
rect 132542 243922 162834 243978
rect 162890 243922 162958 243978
rect 163014 243922 163082 243978
rect 163138 243922 163206 243978
rect 163262 243922 193554 243978
rect 193610 243922 193678 243978
rect 193734 243922 193802 243978
rect 193858 243922 193926 243978
rect 193982 243922 224274 243978
rect 224330 243922 224398 243978
rect 224454 243922 224522 243978
rect 224578 243922 224646 243978
rect 224702 243922 254994 243978
rect 255050 243922 255118 243978
rect 255174 243922 255242 243978
rect 255298 243922 255366 243978
rect 255422 243922 285714 243978
rect 285770 243922 285838 243978
rect 285894 243922 285962 243978
rect 286018 243922 286086 243978
rect 286142 243922 316434 243978
rect 316490 243922 316558 243978
rect 316614 243922 316682 243978
rect 316738 243922 316806 243978
rect 316862 243922 347154 243978
rect 347210 243922 347278 243978
rect 347334 243922 347402 243978
rect 347458 243922 347526 243978
rect 347582 243922 377874 243978
rect 377930 243922 377998 243978
rect 378054 243922 378122 243978
rect 378178 243922 378246 243978
rect 378302 243922 408594 243978
rect 408650 243922 408718 243978
rect 408774 243922 408842 243978
rect 408898 243922 408966 243978
rect 409022 243922 439314 243978
rect 439370 243922 439438 243978
rect 439494 243922 439562 243978
rect 439618 243922 439686 243978
rect 439742 243922 470034 243978
rect 470090 243922 470158 243978
rect 470214 243922 470282 243978
rect 470338 243922 470406 243978
rect 470462 243922 500754 243978
rect 500810 243922 500878 243978
rect 500934 243922 501002 243978
rect 501058 243922 501126 243978
rect 501182 243922 531474 243978
rect 531530 243922 531598 243978
rect 531654 243922 531722 243978
rect 531778 243922 531846 243978
rect 531902 243922 562194 243978
rect 562250 243922 562318 243978
rect 562374 243922 562442 243978
rect 562498 243922 562566 243978
rect 562622 243922 592914 243978
rect 592970 243922 593038 243978
rect 593094 243922 593162 243978
rect 593218 243922 593286 243978
rect 593342 243922 597456 243978
rect 597512 243922 597580 243978
rect 597636 243922 597704 243978
rect 597760 243922 597828 243978
rect 597884 243922 597980 243978
rect -1916 243826 597980 243922
rect -1916 238350 597980 238446
rect -1916 238294 -860 238350
rect -804 238294 -736 238350
rect -680 238294 -612 238350
rect -556 238294 -488 238350
rect -432 238294 5514 238350
rect 5570 238294 5638 238350
rect 5694 238294 5762 238350
rect 5818 238294 5886 238350
rect 5942 238294 36234 238350
rect 36290 238294 36358 238350
rect 36414 238294 36482 238350
rect 36538 238294 36606 238350
rect 36662 238294 66954 238350
rect 67010 238294 67078 238350
rect 67134 238294 67202 238350
rect 67258 238294 67326 238350
rect 67382 238294 97674 238350
rect 97730 238294 97798 238350
rect 97854 238294 97922 238350
rect 97978 238294 98046 238350
rect 98102 238294 128394 238350
rect 128450 238294 128518 238350
rect 128574 238294 128642 238350
rect 128698 238294 128766 238350
rect 128822 238294 159114 238350
rect 159170 238294 159238 238350
rect 159294 238294 159362 238350
rect 159418 238294 159486 238350
rect 159542 238294 189834 238350
rect 189890 238294 189958 238350
rect 190014 238294 190082 238350
rect 190138 238294 190206 238350
rect 190262 238294 220554 238350
rect 220610 238294 220678 238350
rect 220734 238294 220802 238350
rect 220858 238294 220926 238350
rect 220982 238294 251274 238350
rect 251330 238294 251398 238350
rect 251454 238294 251522 238350
rect 251578 238294 251646 238350
rect 251702 238294 281994 238350
rect 282050 238294 282118 238350
rect 282174 238294 282242 238350
rect 282298 238294 282366 238350
rect 282422 238294 312714 238350
rect 312770 238294 312838 238350
rect 312894 238294 312962 238350
rect 313018 238294 313086 238350
rect 313142 238294 343434 238350
rect 343490 238294 343558 238350
rect 343614 238294 343682 238350
rect 343738 238294 343806 238350
rect 343862 238294 374154 238350
rect 374210 238294 374278 238350
rect 374334 238294 374402 238350
rect 374458 238294 374526 238350
rect 374582 238294 404874 238350
rect 404930 238294 404998 238350
rect 405054 238294 405122 238350
rect 405178 238294 405246 238350
rect 405302 238294 435594 238350
rect 435650 238294 435718 238350
rect 435774 238294 435842 238350
rect 435898 238294 435966 238350
rect 436022 238294 466314 238350
rect 466370 238294 466438 238350
rect 466494 238294 466562 238350
rect 466618 238294 466686 238350
rect 466742 238294 497034 238350
rect 497090 238294 497158 238350
rect 497214 238294 497282 238350
rect 497338 238294 497406 238350
rect 497462 238294 527754 238350
rect 527810 238294 527878 238350
rect 527934 238294 528002 238350
rect 528058 238294 528126 238350
rect 528182 238294 558474 238350
rect 558530 238294 558598 238350
rect 558654 238294 558722 238350
rect 558778 238294 558846 238350
rect 558902 238294 589194 238350
rect 589250 238294 589318 238350
rect 589374 238294 589442 238350
rect 589498 238294 589566 238350
rect 589622 238294 596496 238350
rect 596552 238294 596620 238350
rect 596676 238294 596744 238350
rect 596800 238294 596868 238350
rect 596924 238294 597980 238350
rect -1916 238226 597980 238294
rect -1916 238170 -860 238226
rect -804 238170 -736 238226
rect -680 238170 -612 238226
rect -556 238170 -488 238226
rect -432 238170 5514 238226
rect 5570 238170 5638 238226
rect 5694 238170 5762 238226
rect 5818 238170 5886 238226
rect 5942 238170 36234 238226
rect 36290 238170 36358 238226
rect 36414 238170 36482 238226
rect 36538 238170 36606 238226
rect 36662 238170 66954 238226
rect 67010 238170 67078 238226
rect 67134 238170 67202 238226
rect 67258 238170 67326 238226
rect 67382 238170 97674 238226
rect 97730 238170 97798 238226
rect 97854 238170 97922 238226
rect 97978 238170 98046 238226
rect 98102 238170 128394 238226
rect 128450 238170 128518 238226
rect 128574 238170 128642 238226
rect 128698 238170 128766 238226
rect 128822 238170 159114 238226
rect 159170 238170 159238 238226
rect 159294 238170 159362 238226
rect 159418 238170 159486 238226
rect 159542 238170 189834 238226
rect 189890 238170 189958 238226
rect 190014 238170 190082 238226
rect 190138 238170 190206 238226
rect 190262 238170 220554 238226
rect 220610 238170 220678 238226
rect 220734 238170 220802 238226
rect 220858 238170 220926 238226
rect 220982 238170 251274 238226
rect 251330 238170 251398 238226
rect 251454 238170 251522 238226
rect 251578 238170 251646 238226
rect 251702 238170 281994 238226
rect 282050 238170 282118 238226
rect 282174 238170 282242 238226
rect 282298 238170 282366 238226
rect 282422 238170 312714 238226
rect 312770 238170 312838 238226
rect 312894 238170 312962 238226
rect 313018 238170 313086 238226
rect 313142 238170 343434 238226
rect 343490 238170 343558 238226
rect 343614 238170 343682 238226
rect 343738 238170 343806 238226
rect 343862 238170 374154 238226
rect 374210 238170 374278 238226
rect 374334 238170 374402 238226
rect 374458 238170 374526 238226
rect 374582 238170 404874 238226
rect 404930 238170 404998 238226
rect 405054 238170 405122 238226
rect 405178 238170 405246 238226
rect 405302 238170 435594 238226
rect 435650 238170 435718 238226
rect 435774 238170 435842 238226
rect 435898 238170 435966 238226
rect 436022 238170 466314 238226
rect 466370 238170 466438 238226
rect 466494 238170 466562 238226
rect 466618 238170 466686 238226
rect 466742 238170 497034 238226
rect 497090 238170 497158 238226
rect 497214 238170 497282 238226
rect 497338 238170 497406 238226
rect 497462 238170 527754 238226
rect 527810 238170 527878 238226
rect 527934 238170 528002 238226
rect 528058 238170 528126 238226
rect 528182 238170 558474 238226
rect 558530 238170 558598 238226
rect 558654 238170 558722 238226
rect 558778 238170 558846 238226
rect 558902 238170 589194 238226
rect 589250 238170 589318 238226
rect 589374 238170 589442 238226
rect 589498 238170 589566 238226
rect 589622 238170 596496 238226
rect 596552 238170 596620 238226
rect 596676 238170 596744 238226
rect 596800 238170 596868 238226
rect 596924 238170 597980 238226
rect -1916 238102 597980 238170
rect -1916 238046 -860 238102
rect -804 238046 -736 238102
rect -680 238046 -612 238102
rect -556 238046 -488 238102
rect -432 238046 5514 238102
rect 5570 238046 5638 238102
rect 5694 238046 5762 238102
rect 5818 238046 5886 238102
rect 5942 238046 36234 238102
rect 36290 238046 36358 238102
rect 36414 238046 36482 238102
rect 36538 238046 36606 238102
rect 36662 238046 66954 238102
rect 67010 238046 67078 238102
rect 67134 238046 67202 238102
rect 67258 238046 67326 238102
rect 67382 238046 97674 238102
rect 97730 238046 97798 238102
rect 97854 238046 97922 238102
rect 97978 238046 98046 238102
rect 98102 238046 128394 238102
rect 128450 238046 128518 238102
rect 128574 238046 128642 238102
rect 128698 238046 128766 238102
rect 128822 238046 159114 238102
rect 159170 238046 159238 238102
rect 159294 238046 159362 238102
rect 159418 238046 159486 238102
rect 159542 238046 189834 238102
rect 189890 238046 189958 238102
rect 190014 238046 190082 238102
rect 190138 238046 190206 238102
rect 190262 238046 220554 238102
rect 220610 238046 220678 238102
rect 220734 238046 220802 238102
rect 220858 238046 220926 238102
rect 220982 238046 251274 238102
rect 251330 238046 251398 238102
rect 251454 238046 251522 238102
rect 251578 238046 251646 238102
rect 251702 238046 281994 238102
rect 282050 238046 282118 238102
rect 282174 238046 282242 238102
rect 282298 238046 282366 238102
rect 282422 238046 312714 238102
rect 312770 238046 312838 238102
rect 312894 238046 312962 238102
rect 313018 238046 313086 238102
rect 313142 238046 343434 238102
rect 343490 238046 343558 238102
rect 343614 238046 343682 238102
rect 343738 238046 343806 238102
rect 343862 238046 374154 238102
rect 374210 238046 374278 238102
rect 374334 238046 374402 238102
rect 374458 238046 374526 238102
rect 374582 238046 404874 238102
rect 404930 238046 404998 238102
rect 405054 238046 405122 238102
rect 405178 238046 405246 238102
rect 405302 238046 435594 238102
rect 435650 238046 435718 238102
rect 435774 238046 435842 238102
rect 435898 238046 435966 238102
rect 436022 238046 466314 238102
rect 466370 238046 466438 238102
rect 466494 238046 466562 238102
rect 466618 238046 466686 238102
rect 466742 238046 497034 238102
rect 497090 238046 497158 238102
rect 497214 238046 497282 238102
rect 497338 238046 497406 238102
rect 497462 238046 527754 238102
rect 527810 238046 527878 238102
rect 527934 238046 528002 238102
rect 528058 238046 528126 238102
rect 528182 238046 558474 238102
rect 558530 238046 558598 238102
rect 558654 238046 558722 238102
rect 558778 238046 558846 238102
rect 558902 238046 589194 238102
rect 589250 238046 589318 238102
rect 589374 238046 589442 238102
rect 589498 238046 589566 238102
rect 589622 238046 596496 238102
rect 596552 238046 596620 238102
rect 596676 238046 596744 238102
rect 596800 238046 596868 238102
rect 596924 238046 597980 238102
rect -1916 237978 597980 238046
rect -1916 237922 -860 237978
rect -804 237922 -736 237978
rect -680 237922 -612 237978
rect -556 237922 -488 237978
rect -432 237922 5514 237978
rect 5570 237922 5638 237978
rect 5694 237922 5762 237978
rect 5818 237922 5886 237978
rect 5942 237922 36234 237978
rect 36290 237922 36358 237978
rect 36414 237922 36482 237978
rect 36538 237922 36606 237978
rect 36662 237922 66954 237978
rect 67010 237922 67078 237978
rect 67134 237922 67202 237978
rect 67258 237922 67326 237978
rect 67382 237922 97674 237978
rect 97730 237922 97798 237978
rect 97854 237922 97922 237978
rect 97978 237922 98046 237978
rect 98102 237922 128394 237978
rect 128450 237922 128518 237978
rect 128574 237922 128642 237978
rect 128698 237922 128766 237978
rect 128822 237922 159114 237978
rect 159170 237922 159238 237978
rect 159294 237922 159362 237978
rect 159418 237922 159486 237978
rect 159542 237922 189834 237978
rect 189890 237922 189958 237978
rect 190014 237922 190082 237978
rect 190138 237922 190206 237978
rect 190262 237922 220554 237978
rect 220610 237922 220678 237978
rect 220734 237922 220802 237978
rect 220858 237922 220926 237978
rect 220982 237922 251274 237978
rect 251330 237922 251398 237978
rect 251454 237922 251522 237978
rect 251578 237922 251646 237978
rect 251702 237922 281994 237978
rect 282050 237922 282118 237978
rect 282174 237922 282242 237978
rect 282298 237922 282366 237978
rect 282422 237922 312714 237978
rect 312770 237922 312838 237978
rect 312894 237922 312962 237978
rect 313018 237922 313086 237978
rect 313142 237922 343434 237978
rect 343490 237922 343558 237978
rect 343614 237922 343682 237978
rect 343738 237922 343806 237978
rect 343862 237922 374154 237978
rect 374210 237922 374278 237978
rect 374334 237922 374402 237978
rect 374458 237922 374526 237978
rect 374582 237922 404874 237978
rect 404930 237922 404998 237978
rect 405054 237922 405122 237978
rect 405178 237922 405246 237978
rect 405302 237922 435594 237978
rect 435650 237922 435718 237978
rect 435774 237922 435842 237978
rect 435898 237922 435966 237978
rect 436022 237922 466314 237978
rect 466370 237922 466438 237978
rect 466494 237922 466562 237978
rect 466618 237922 466686 237978
rect 466742 237922 497034 237978
rect 497090 237922 497158 237978
rect 497214 237922 497282 237978
rect 497338 237922 497406 237978
rect 497462 237922 527754 237978
rect 527810 237922 527878 237978
rect 527934 237922 528002 237978
rect 528058 237922 528126 237978
rect 528182 237922 558474 237978
rect 558530 237922 558598 237978
rect 558654 237922 558722 237978
rect 558778 237922 558846 237978
rect 558902 237922 589194 237978
rect 589250 237922 589318 237978
rect 589374 237922 589442 237978
rect 589498 237922 589566 237978
rect 589622 237922 596496 237978
rect 596552 237922 596620 237978
rect 596676 237922 596744 237978
rect 596800 237922 596868 237978
rect 596924 237922 597980 237978
rect -1916 237826 597980 237922
rect -1916 226350 597980 226446
rect -1916 226294 -1820 226350
rect -1764 226294 -1696 226350
rect -1640 226294 -1572 226350
rect -1516 226294 -1448 226350
rect -1392 226294 9234 226350
rect 9290 226294 9358 226350
rect 9414 226294 9482 226350
rect 9538 226294 9606 226350
rect 9662 226294 39954 226350
rect 40010 226294 40078 226350
rect 40134 226294 40202 226350
rect 40258 226294 40326 226350
rect 40382 226294 70674 226350
rect 70730 226294 70798 226350
rect 70854 226294 70922 226350
rect 70978 226294 71046 226350
rect 71102 226294 101394 226350
rect 101450 226294 101518 226350
rect 101574 226294 101642 226350
rect 101698 226294 101766 226350
rect 101822 226294 132114 226350
rect 132170 226294 132238 226350
rect 132294 226294 132362 226350
rect 132418 226294 132486 226350
rect 132542 226294 162834 226350
rect 162890 226294 162958 226350
rect 163014 226294 163082 226350
rect 163138 226294 163206 226350
rect 163262 226294 193554 226350
rect 193610 226294 193678 226350
rect 193734 226294 193802 226350
rect 193858 226294 193926 226350
rect 193982 226294 224274 226350
rect 224330 226294 224398 226350
rect 224454 226294 224522 226350
rect 224578 226294 224646 226350
rect 224702 226294 254994 226350
rect 255050 226294 255118 226350
rect 255174 226294 255242 226350
rect 255298 226294 255366 226350
rect 255422 226294 285714 226350
rect 285770 226294 285838 226350
rect 285894 226294 285962 226350
rect 286018 226294 286086 226350
rect 286142 226294 316434 226350
rect 316490 226294 316558 226350
rect 316614 226294 316682 226350
rect 316738 226294 316806 226350
rect 316862 226294 347154 226350
rect 347210 226294 347278 226350
rect 347334 226294 347402 226350
rect 347458 226294 347526 226350
rect 347582 226294 377874 226350
rect 377930 226294 377998 226350
rect 378054 226294 378122 226350
rect 378178 226294 378246 226350
rect 378302 226294 408594 226350
rect 408650 226294 408718 226350
rect 408774 226294 408842 226350
rect 408898 226294 408966 226350
rect 409022 226294 439314 226350
rect 439370 226294 439438 226350
rect 439494 226294 439562 226350
rect 439618 226294 439686 226350
rect 439742 226294 470034 226350
rect 470090 226294 470158 226350
rect 470214 226294 470282 226350
rect 470338 226294 470406 226350
rect 470462 226294 500754 226350
rect 500810 226294 500878 226350
rect 500934 226294 501002 226350
rect 501058 226294 501126 226350
rect 501182 226294 531474 226350
rect 531530 226294 531598 226350
rect 531654 226294 531722 226350
rect 531778 226294 531846 226350
rect 531902 226294 562194 226350
rect 562250 226294 562318 226350
rect 562374 226294 562442 226350
rect 562498 226294 562566 226350
rect 562622 226294 592914 226350
rect 592970 226294 593038 226350
rect 593094 226294 593162 226350
rect 593218 226294 593286 226350
rect 593342 226294 597456 226350
rect 597512 226294 597580 226350
rect 597636 226294 597704 226350
rect 597760 226294 597828 226350
rect 597884 226294 597980 226350
rect -1916 226226 597980 226294
rect -1916 226170 -1820 226226
rect -1764 226170 -1696 226226
rect -1640 226170 -1572 226226
rect -1516 226170 -1448 226226
rect -1392 226170 9234 226226
rect 9290 226170 9358 226226
rect 9414 226170 9482 226226
rect 9538 226170 9606 226226
rect 9662 226170 39954 226226
rect 40010 226170 40078 226226
rect 40134 226170 40202 226226
rect 40258 226170 40326 226226
rect 40382 226170 70674 226226
rect 70730 226170 70798 226226
rect 70854 226170 70922 226226
rect 70978 226170 71046 226226
rect 71102 226170 101394 226226
rect 101450 226170 101518 226226
rect 101574 226170 101642 226226
rect 101698 226170 101766 226226
rect 101822 226170 132114 226226
rect 132170 226170 132238 226226
rect 132294 226170 132362 226226
rect 132418 226170 132486 226226
rect 132542 226170 162834 226226
rect 162890 226170 162958 226226
rect 163014 226170 163082 226226
rect 163138 226170 163206 226226
rect 163262 226170 193554 226226
rect 193610 226170 193678 226226
rect 193734 226170 193802 226226
rect 193858 226170 193926 226226
rect 193982 226170 224274 226226
rect 224330 226170 224398 226226
rect 224454 226170 224522 226226
rect 224578 226170 224646 226226
rect 224702 226170 254994 226226
rect 255050 226170 255118 226226
rect 255174 226170 255242 226226
rect 255298 226170 255366 226226
rect 255422 226170 285714 226226
rect 285770 226170 285838 226226
rect 285894 226170 285962 226226
rect 286018 226170 286086 226226
rect 286142 226170 316434 226226
rect 316490 226170 316558 226226
rect 316614 226170 316682 226226
rect 316738 226170 316806 226226
rect 316862 226170 347154 226226
rect 347210 226170 347278 226226
rect 347334 226170 347402 226226
rect 347458 226170 347526 226226
rect 347582 226170 377874 226226
rect 377930 226170 377998 226226
rect 378054 226170 378122 226226
rect 378178 226170 378246 226226
rect 378302 226170 408594 226226
rect 408650 226170 408718 226226
rect 408774 226170 408842 226226
rect 408898 226170 408966 226226
rect 409022 226170 439314 226226
rect 439370 226170 439438 226226
rect 439494 226170 439562 226226
rect 439618 226170 439686 226226
rect 439742 226170 470034 226226
rect 470090 226170 470158 226226
rect 470214 226170 470282 226226
rect 470338 226170 470406 226226
rect 470462 226170 500754 226226
rect 500810 226170 500878 226226
rect 500934 226170 501002 226226
rect 501058 226170 501126 226226
rect 501182 226170 531474 226226
rect 531530 226170 531598 226226
rect 531654 226170 531722 226226
rect 531778 226170 531846 226226
rect 531902 226170 562194 226226
rect 562250 226170 562318 226226
rect 562374 226170 562442 226226
rect 562498 226170 562566 226226
rect 562622 226170 592914 226226
rect 592970 226170 593038 226226
rect 593094 226170 593162 226226
rect 593218 226170 593286 226226
rect 593342 226170 597456 226226
rect 597512 226170 597580 226226
rect 597636 226170 597704 226226
rect 597760 226170 597828 226226
rect 597884 226170 597980 226226
rect -1916 226102 597980 226170
rect -1916 226046 -1820 226102
rect -1764 226046 -1696 226102
rect -1640 226046 -1572 226102
rect -1516 226046 -1448 226102
rect -1392 226046 9234 226102
rect 9290 226046 9358 226102
rect 9414 226046 9482 226102
rect 9538 226046 9606 226102
rect 9662 226046 39954 226102
rect 40010 226046 40078 226102
rect 40134 226046 40202 226102
rect 40258 226046 40326 226102
rect 40382 226046 70674 226102
rect 70730 226046 70798 226102
rect 70854 226046 70922 226102
rect 70978 226046 71046 226102
rect 71102 226046 101394 226102
rect 101450 226046 101518 226102
rect 101574 226046 101642 226102
rect 101698 226046 101766 226102
rect 101822 226046 132114 226102
rect 132170 226046 132238 226102
rect 132294 226046 132362 226102
rect 132418 226046 132486 226102
rect 132542 226046 162834 226102
rect 162890 226046 162958 226102
rect 163014 226046 163082 226102
rect 163138 226046 163206 226102
rect 163262 226046 193554 226102
rect 193610 226046 193678 226102
rect 193734 226046 193802 226102
rect 193858 226046 193926 226102
rect 193982 226046 224274 226102
rect 224330 226046 224398 226102
rect 224454 226046 224522 226102
rect 224578 226046 224646 226102
rect 224702 226046 254994 226102
rect 255050 226046 255118 226102
rect 255174 226046 255242 226102
rect 255298 226046 255366 226102
rect 255422 226046 285714 226102
rect 285770 226046 285838 226102
rect 285894 226046 285962 226102
rect 286018 226046 286086 226102
rect 286142 226046 316434 226102
rect 316490 226046 316558 226102
rect 316614 226046 316682 226102
rect 316738 226046 316806 226102
rect 316862 226046 347154 226102
rect 347210 226046 347278 226102
rect 347334 226046 347402 226102
rect 347458 226046 347526 226102
rect 347582 226046 377874 226102
rect 377930 226046 377998 226102
rect 378054 226046 378122 226102
rect 378178 226046 378246 226102
rect 378302 226046 408594 226102
rect 408650 226046 408718 226102
rect 408774 226046 408842 226102
rect 408898 226046 408966 226102
rect 409022 226046 439314 226102
rect 439370 226046 439438 226102
rect 439494 226046 439562 226102
rect 439618 226046 439686 226102
rect 439742 226046 470034 226102
rect 470090 226046 470158 226102
rect 470214 226046 470282 226102
rect 470338 226046 470406 226102
rect 470462 226046 500754 226102
rect 500810 226046 500878 226102
rect 500934 226046 501002 226102
rect 501058 226046 501126 226102
rect 501182 226046 531474 226102
rect 531530 226046 531598 226102
rect 531654 226046 531722 226102
rect 531778 226046 531846 226102
rect 531902 226046 562194 226102
rect 562250 226046 562318 226102
rect 562374 226046 562442 226102
rect 562498 226046 562566 226102
rect 562622 226046 592914 226102
rect 592970 226046 593038 226102
rect 593094 226046 593162 226102
rect 593218 226046 593286 226102
rect 593342 226046 597456 226102
rect 597512 226046 597580 226102
rect 597636 226046 597704 226102
rect 597760 226046 597828 226102
rect 597884 226046 597980 226102
rect -1916 225978 597980 226046
rect -1916 225922 -1820 225978
rect -1764 225922 -1696 225978
rect -1640 225922 -1572 225978
rect -1516 225922 -1448 225978
rect -1392 225922 9234 225978
rect 9290 225922 9358 225978
rect 9414 225922 9482 225978
rect 9538 225922 9606 225978
rect 9662 225922 39954 225978
rect 40010 225922 40078 225978
rect 40134 225922 40202 225978
rect 40258 225922 40326 225978
rect 40382 225922 70674 225978
rect 70730 225922 70798 225978
rect 70854 225922 70922 225978
rect 70978 225922 71046 225978
rect 71102 225922 101394 225978
rect 101450 225922 101518 225978
rect 101574 225922 101642 225978
rect 101698 225922 101766 225978
rect 101822 225922 132114 225978
rect 132170 225922 132238 225978
rect 132294 225922 132362 225978
rect 132418 225922 132486 225978
rect 132542 225922 162834 225978
rect 162890 225922 162958 225978
rect 163014 225922 163082 225978
rect 163138 225922 163206 225978
rect 163262 225922 193554 225978
rect 193610 225922 193678 225978
rect 193734 225922 193802 225978
rect 193858 225922 193926 225978
rect 193982 225922 224274 225978
rect 224330 225922 224398 225978
rect 224454 225922 224522 225978
rect 224578 225922 224646 225978
rect 224702 225922 254994 225978
rect 255050 225922 255118 225978
rect 255174 225922 255242 225978
rect 255298 225922 255366 225978
rect 255422 225922 285714 225978
rect 285770 225922 285838 225978
rect 285894 225922 285962 225978
rect 286018 225922 286086 225978
rect 286142 225922 316434 225978
rect 316490 225922 316558 225978
rect 316614 225922 316682 225978
rect 316738 225922 316806 225978
rect 316862 225922 347154 225978
rect 347210 225922 347278 225978
rect 347334 225922 347402 225978
rect 347458 225922 347526 225978
rect 347582 225922 377874 225978
rect 377930 225922 377998 225978
rect 378054 225922 378122 225978
rect 378178 225922 378246 225978
rect 378302 225922 408594 225978
rect 408650 225922 408718 225978
rect 408774 225922 408842 225978
rect 408898 225922 408966 225978
rect 409022 225922 439314 225978
rect 439370 225922 439438 225978
rect 439494 225922 439562 225978
rect 439618 225922 439686 225978
rect 439742 225922 470034 225978
rect 470090 225922 470158 225978
rect 470214 225922 470282 225978
rect 470338 225922 470406 225978
rect 470462 225922 500754 225978
rect 500810 225922 500878 225978
rect 500934 225922 501002 225978
rect 501058 225922 501126 225978
rect 501182 225922 531474 225978
rect 531530 225922 531598 225978
rect 531654 225922 531722 225978
rect 531778 225922 531846 225978
rect 531902 225922 562194 225978
rect 562250 225922 562318 225978
rect 562374 225922 562442 225978
rect 562498 225922 562566 225978
rect 562622 225922 592914 225978
rect 592970 225922 593038 225978
rect 593094 225922 593162 225978
rect 593218 225922 593286 225978
rect 593342 225922 597456 225978
rect 597512 225922 597580 225978
rect 597636 225922 597704 225978
rect 597760 225922 597828 225978
rect 597884 225922 597980 225978
rect -1916 225826 597980 225922
rect -1916 220350 597980 220446
rect -1916 220294 -860 220350
rect -804 220294 -736 220350
rect -680 220294 -612 220350
rect -556 220294 -488 220350
rect -432 220294 5514 220350
rect 5570 220294 5638 220350
rect 5694 220294 5762 220350
rect 5818 220294 5886 220350
rect 5942 220294 36234 220350
rect 36290 220294 36358 220350
rect 36414 220294 36482 220350
rect 36538 220294 36606 220350
rect 36662 220294 66954 220350
rect 67010 220294 67078 220350
rect 67134 220294 67202 220350
rect 67258 220294 67326 220350
rect 67382 220294 97674 220350
rect 97730 220294 97798 220350
rect 97854 220294 97922 220350
rect 97978 220294 98046 220350
rect 98102 220294 128394 220350
rect 128450 220294 128518 220350
rect 128574 220294 128642 220350
rect 128698 220294 128766 220350
rect 128822 220294 159114 220350
rect 159170 220294 159238 220350
rect 159294 220294 159362 220350
rect 159418 220294 159486 220350
rect 159542 220294 189834 220350
rect 189890 220294 189958 220350
rect 190014 220294 190082 220350
rect 190138 220294 190206 220350
rect 190262 220294 220554 220350
rect 220610 220294 220678 220350
rect 220734 220294 220802 220350
rect 220858 220294 220926 220350
rect 220982 220294 251274 220350
rect 251330 220294 251398 220350
rect 251454 220294 251522 220350
rect 251578 220294 251646 220350
rect 251702 220294 281994 220350
rect 282050 220294 282118 220350
rect 282174 220294 282242 220350
rect 282298 220294 282366 220350
rect 282422 220294 312714 220350
rect 312770 220294 312838 220350
rect 312894 220294 312962 220350
rect 313018 220294 313086 220350
rect 313142 220294 343434 220350
rect 343490 220294 343558 220350
rect 343614 220294 343682 220350
rect 343738 220294 343806 220350
rect 343862 220294 374154 220350
rect 374210 220294 374278 220350
rect 374334 220294 374402 220350
rect 374458 220294 374526 220350
rect 374582 220294 404874 220350
rect 404930 220294 404998 220350
rect 405054 220294 405122 220350
rect 405178 220294 405246 220350
rect 405302 220294 435594 220350
rect 435650 220294 435718 220350
rect 435774 220294 435842 220350
rect 435898 220294 435966 220350
rect 436022 220294 466314 220350
rect 466370 220294 466438 220350
rect 466494 220294 466562 220350
rect 466618 220294 466686 220350
rect 466742 220294 497034 220350
rect 497090 220294 497158 220350
rect 497214 220294 497282 220350
rect 497338 220294 497406 220350
rect 497462 220294 527754 220350
rect 527810 220294 527878 220350
rect 527934 220294 528002 220350
rect 528058 220294 528126 220350
rect 528182 220294 558474 220350
rect 558530 220294 558598 220350
rect 558654 220294 558722 220350
rect 558778 220294 558846 220350
rect 558902 220294 589194 220350
rect 589250 220294 589318 220350
rect 589374 220294 589442 220350
rect 589498 220294 589566 220350
rect 589622 220294 596496 220350
rect 596552 220294 596620 220350
rect 596676 220294 596744 220350
rect 596800 220294 596868 220350
rect 596924 220294 597980 220350
rect -1916 220226 597980 220294
rect -1916 220170 -860 220226
rect -804 220170 -736 220226
rect -680 220170 -612 220226
rect -556 220170 -488 220226
rect -432 220170 5514 220226
rect 5570 220170 5638 220226
rect 5694 220170 5762 220226
rect 5818 220170 5886 220226
rect 5942 220170 36234 220226
rect 36290 220170 36358 220226
rect 36414 220170 36482 220226
rect 36538 220170 36606 220226
rect 36662 220170 66954 220226
rect 67010 220170 67078 220226
rect 67134 220170 67202 220226
rect 67258 220170 67326 220226
rect 67382 220170 97674 220226
rect 97730 220170 97798 220226
rect 97854 220170 97922 220226
rect 97978 220170 98046 220226
rect 98102 220170 128394 220226
rect 128450 220170 128518 220226
rect 128574 220170 128642 220226
rect 128698 220170 128766 220226
rect 128822 220170 159114 220226
rect 159170 220170 159238 220226
rect 159294 220170 159362 220226
rect 159418 220170 159486 220226
rect 159542 220170 189834 220226
rect 189890 220170 189958 220226
rect 190014 220170 190082 220226
rect 190138 220170 190206 220226
rect 190262 220170 220554 220226
rect 220610 220170 220678 220226
rect 220734 220170 220802 220226
rect 220858 220170 220926 220226
rect 220982 220170 251274 220226
rect 251330 220170 251398 220226
rect 251454 220170 251522 220226
rect 251578 220170 251646 220226
rect 251702 220170 281994 220226
rect 282050 220170 282118 220226
rect 282174 220170 282242 220226
rect 282298 220170 282366 220226
rect 282422 220170 312714 220226
rect 312770 220170 312838 220226
rect 312894 220170 312962 220226
rect 313018 220170 313086 220226
rect 313142 220170 343434 220226
rect 343490 220170 343558 220226
rect 343614 220170 343682 220226
rect 343738 220170 343806 220226
rect 343862 220170 374154 220226
rect 374210 220170 374278 220226
rect 374334 220170 374402 220226
rect 374458 220170 374526 220226
rect 374582 220170 404874 220226
rect 404930 220170 404998 220226
rect 405054 220170 405122 220226
rect 405178 220170 405246 220226
rect 405302 220170 435594 220226
rect 435650 220170 435718 220226
rect 435774 220170 435842 220226
rect 435898 220170 435966 220226
rect 436022 220170 466314 220226
rect 466370 220170 466438 220226
rect 466494 220170 466562 220226
rect 466618 220170 466686 220226
rect 466742 220170 497034 220226
rect 497090 220170 497158 220226
rect 497214 220170 497282 220226
rect 497338 220170 497406 220226
rect 497462 220170 527754 220226
rect 527810 220170 527878 220226
rect 527934 220170 528002 220226
rect 528058 220170 528126 220226
rect 528182 220170 558474 220226
rect 558530 220170 558598 220226
rect 558654 220170 558722 220226
rect 558778 220170 558846 220226
rect 558902 220170 589194 220226
rect 589250 220170 589318 220226
rect 589374 220170 589442 220226
rect 589498 220170 589566 220226
rect 589622 220170 596496 220226
rect 596552 220170 596620 220226
rect 596676 220170 596744 220226
rect 596800 220170 596868 220226
rect 596924 220170 597980 220226
rect -1916 220102 597980 220170
rect -1916 220046 -860 220102
rect -804 220046 -736 220102
rect -680 220046 -612 220102
rect -556 220046 -488 220102
rect -432 220046 5514 220102
rect 5570 220046 5638 220102
rect 5694 220046 5762 220102
rect 5818 220046 5886 220102
rect 5942 220046 36234 220102
rect 36290 220046 36358 220102
rect 36414 220046 36482 220102
rect 36538 220046 36606 220102
rect 36662 220046 66954 220102
rect 67010 220046 67078 220102
rect 67134 220046 67202 220102
rect 67258 220046 67326 220102
rect 67382 220046 97674 220102
rect 97730 220046 97798 220102
rect 97854 220046 97922 220102
rect 97978 220046 98046 220102
rect 98102 220046 128394 220102
rect 128450 220046 128518 220102
rect 128574 220046 128642 220102
rect 128698 220046 128766 220102
rect 128822 220046 159114 220102
rect 159170 220046 159238 220102
rect 159294 220046 159362 220102
rect 159418 220046 159486 220102
rect 159542 220046 189834 220102
rect 189890 220046 189958 220102
rect 190014 220046 190082 220102
rect 190138 220046 190206 220102
rect 190262 220046 220554 220102
rect 220610 220046 220678 220102
rect 220734 220046 220802 220102
rect 220858 220046 220926 220102
rect 220982 220046 251274 220102
rect 251330 220046 251398 220102
rect 251454 220046 251522 220102
rect 251578 220046 251646 220102
rect 251702 220046 281994 220102
rect 282050 220046 282118 220102
rect 282174 220046 282242 220102
rect 282298 220046 282366 220102
rect 282422 220046 312714 220102
rect 312770 220046 312838 220102
rect 312894 220046 312962 220102
rect 313018 220046 313086 220102
rect 313142 220046 343434 220102
rect 343490 220046 343558 220102
rect 343614 220046 343682 220102
rect 343738 220046 343806 220102
rect 343862 220046 374154 220102
rect 374210 220046 374278 220102
rect 374334 220046 374402 220102
rect 374458 220046 374526 220102
rect 374582 220046 404874 220102
rect 404930 220046 404998 220102
rect 405054 220046 405122 220102
rect 405178 220046 405246 220102
rect 405302 220046 435594 220102
rect 435650 220046 435718 220102
rect 435774 220046 435842 220102
rect 435898 220046 435966 220102
rect 436022 220046 466314 220102
rect 466370 220046 466438 220102
rect 466494 220046 466562 220102
rect 466618 220046 466686 220102
rect 466742 220046 497034 220102
rect 497090 220046 497158 220102
rect 497214 220046 497282 220102
rect 497338 220046 497406 220102
rect 497462 220046 527754 220102
rect 527810 220046 527878 220102
rect 527934 220046 528002 220102
rect 528058 220046 528126 220102
rect 528182 220046 558474 220102
rect 558530 220046 558598 220102
rect 558654 220046 558722 220102
rect 558778 220046 558846 220102
rect 558902 220046 589194 220102
rect 589250 220046 589318 220102
rect 589374 220046 589442 220102
rect 589498 220046 589566 220102
rect 589622 220046 596496 220102
rect 596552 220046 596620 220102
rect 596676 220046 596744 220102
rect 596800 220046 596868 220102
rect 596924 220046 597980 220102
rect -1916 219978 597980 220046
rect -1916 219922 -860 219978
rect -804 219922 -736 219978
rect -680 219922 -612 219978
rect -556 219922 -488 219978
rect -432 219922 5514 219978
rect 5570 219922 5638 219978
rect 5694 219922 5762 219978
rect 5818 219922 5886 219978
rect 5942 219922 36234 219978
rect 36290 219922 36358 219978
rect 36414 219922 36482 219978
rect 36538 219922 36606 219978
rect 36662 219922 66954 219978
rect 67010 219922 67078 219978
rect 67134 219922 67202 219978
rect 67258 219922 67326 219978
rect 67382 219922 97674 219978
rect 97730 219922 97798 219978
rect 97854 219922 97922 219978
rect 97978 219922 98046 219978
rect 98102 219922 128394 219978
rect 128450 219922 128518 219978
rect 128574 219922 128642 219978
rect 128698 219922 128766 219978
rect 128822 219922 159114 219978
rect 159170 219922 159238 219978
rect 159294 219922 159362 219978
rect 159418 219922 159486 219978
rect 159542 219922 189834 219978
rect 189890 219922 189958 219978
rect 190014 219922 190082 219978
rect 190138 219922 190206 219978
rect 190262 219922 220554 219978
rect 220610 219922 220678 219978
rect 220734 219922 220802 219978
rect 220858 219922 220926 219978
rect 220982 219922 251274 219978
rect 251330 219922 251398 219978
rect 251454 219922 251522 219978
rect 251578 219922 251646 219978
rect 251702 219922 281994 219978
rect 282050 219922 282118 219978
rect 282174 219922 282242 219978
rect 282298 219922 282366 219978
rect 282422 219922 312714 219978
rect 312770 219922 312838 219978
rect 312894 219922 312962 219978
rect 313018 219922 313086 219978
rect 313142 219922 343434 219978
rect 343490 219922 343558 219978
rect 343614 219922 343682 219978
rect 343738 219922 343806 219978
rect 343862 219922 374154 219978
rect 374210 219922 374278 219978
rect 374334 219922 374402 219978
rect 374458 219922 374526 219978
rect 374582 219922 404874 219978
rect 404930 219922 404998 219978
rect 405054 219922 405122 219978
rect 405178 219922 405246 219978
rect 405302 219922 435594 219978
rect 435650 219922 435718 219978
rect 435774 219922 435842 219978
rect 435898 219922 435966 219978
rect 436022 219922 466314 219978
rect 466370 219922 466438 219978
rect 466494 219922 466562 219978
rect 466618 219922 466686 219978
rect 466742 219922 497034 219978
rect 497090 219922 497158 219978
rect 497214 219922 497282 219978
rect 497338 219922 497406 219978
rect 497462 219922 527754 219978
rect 527810 219922 527878 219978
rect 527934 219922 528002 219978
rect 528058 219922 528126 219978
rect 528182 219922 558474 219978
rect 558530 219922 558598 219978
rect 558654 219922 558722 219978
rect 558778 219922 558846 219978
rect 558902 219922 589194 219978
rect 589250 219922 589318 219978
rect 589374 219922 589442 219978
rect 589498 219922 589566 219978
rect 589622 219922 596496 219978
rect 596552 219922 596620 219978
rect 596676 219922 596744 219978
rect 596800 219922 596868 219978
rect 596924 219922 597980 219978
rect -1916 219826 597980 219922
rect -1916 208350 597980 208446
rect -1916 208294 -1820 208350
rect -1764 208294 -1696 208350
rect -1640 208294 -1572 208350
rect -1516 208294 -1448 208350
rect -1392 208294 9234 208350
rect 9290 208294 9358 208350
rect 9414 208294 9482 208350
rect 9538 208294 9606 208350
rect 9662 208294 39954 208350
rect 40010 208294 40078 208350
rect 40134 208294 40202 208350
rect 40258 208294 40326 208350
rect 40382 208294 70674 208350
rect 70730 208294 70798 208350
rect 70854 208294 70922 208350
rect 70978 208294 71046 208350
rect 71102 208294 101394 208350
rect 101450 208294 101518 208350
rect 101574 208294 101642 208350
rect 101698 208294 101766 208350
rect 101822 208294 132114 208350
rect 132170 208294 132238 208350
rect 132294 208294 132362 208350
rect 132418 208294 132486 208350
rect 132542 208294 162834 208350
rect 162890 208294 162958 208350
rect 163014 208294 163082 208350
rect 163138 208294 163206 208350
rect 163262 208294 193554 208350
rect 193610 208294 193678 208350
rect 193734 208294 193802 208350
rect 193858 208294 193926 208350
rect 193982 208294 224274 208350
rect 224330 208294 224398 208350
rect 224454 208294 224522 208350
rect 224578 208294 224646 208350
rect 224702 208294 254994 208350
rect 255050 208294 255118 208350
rect 255174 208294 255242 208350
rect 255298 208294 255366 208350
rect 255422 208294 285714 208350
rect 285770 208294 285838 208350
rect 285894 208294 285962 208350
rect 286018 208294 286086 208350
rect 286142 208294 316434 208350
rect 316490 208294 316558 208350
rect 316614 208294 316682 208350
rect 316738 208294 316806 208350
rect 316862 208294 347154 208350
rect 347210 208294 347278 208350
rect 347334 208294 347402 208350
rect 347458 208294 347526 208350
rect 347582 208294 377874 208350
rect 377930 208294 377998 208350
rect 378054 208294 378122 208350
rect 378178 208294 378246 208350
rect 378302 208294 408594 208350
rect 408650 208294 408718 208350
rect 408774 208294 408842 208350
rect 408898 208294 408966 208350
rect 409022 208294 439314 208350
rect 439370 208294 439438 208350
rect 439494 208294 439562 208350
rect 439618 208294 439686 208350
rect 439742 208294 470034 208350
rect 470090 208294 470158 208350
rect 470214 208294 470282 208350
rect 470338 208294 470406 208350
rect 470462 208294 500754 208350
rect 500810 208294 500878 208350
rect 500934 208294 501002 208350
rect 501058 208294 501126 208350
rect 501182 208294 531474 208350
rect 531530 208294 531598 208350
rect 531654 208294 531722 208350
rect 531778 208294 531846 208350
rect 531902 208294 562194 208350
rect 562250 208294 562318 208350
rect 562374 208294 562442 208350
rect 562498 208294 562566 208350
rect 562622 208294 592914 208350
rect 592970 208294 593038 208350
rect 593094 208294 593162 208350
rect 593218 208294 593286 208350
rect 593342 208294 597456 208350
rect 597512 208294 597580 208350
rect 597636 208294 597704 208350
rect 597760 208294 597828 208350
rect 597884 208294 597980 208350
rect -1916 208226 597980 208294
rect -1916 208170 -1820 208226
rect -1764 208170 -1696 208226
rect -1640 208170 -1572 208226
rect -1516 208170 -1448 208226
rect -1392 208170 9234 208226
rect 9290 208170 9358 208226
rect 9414 208170 9482 208226
rect 9538 208170 9606 208226
rect 9662 208170 39954 208226
rect 40010 208170 40078 208226
rect 40134 208170 40202 208226
rect 40258 208170 40326 208226
rect 40382 208170 70674 208226
rect 70730 208170 70798 208226
rect 70854 208170 70922 208226
rect 70978 208170 71046 208226
rect 71102 208170 101394 208226
rect 101450 208170 101518 208226
rect 101574 208170 101642 208226
rect 101698 208170 101766 208226
rect 101822 208170 132114 208226
rect 132170 208170 132238 208226
rect 132294 208170 132362 208226
rect 132418 208170 132486 208226
rect 132542 208170 162834 208226
rect 162890 208170 162958 208226
rect 163014 208170 163082 208226
rect 163138 208170 163206 208226
rect 163262 208170 193554 208226
rect 193610 208170 193678 208226
rect 193734 208170 193802 208226
rect 193858 208170 193926 208226
rect 193982 208170 224274 208226
rect 224330 208170 224398 208226
rect 224454 208170 224522 208226
rect 224578 208170 224646 208226
rect 224702 208170 254994 208226
rect 255050 208170 255118 208226
rect 255174 208170 255242 208226
rect 255298 208170 255366 208226
rect 255422 208170 285714 208226
rect 285770 208170 285838 208226
rect 285894 208170 285962 208226
rect 286018 208170 286086 208226
rect 286142 208170 316434 208226
rect 316490 208170 316558 208226
rect 316614 208170 316682 208226
rect 316738 208170 316806 208226
rect 316862 208170 347154 208226
rect 347210 208170 347278 208226
rect 347334 208170 347402 208226
rect 347458 208170 347526 208226
rect 347582 208170 377874 208226
rect 377930 208170 377998 208226
rect 378054 208170 378122 208226
rect 378178 208170 378246 208226
rect 378302 208170 408594 208226
rect 408650 208170 408718 208226
rect 408774 208170 408842 208226
rect 408898 208170 408966 208226
rect 409022 208170 439314 208226
rect 439370 208170 439438 208226
rect 439494 208170 439562 208226
rect 439618 208170 439686 208226
rect 439742 208170 470034 208226
rect 470090 208170 470158 208226
rect 470214 208170 470282 208226
rect 470338 208170 470406 208226
rect 470462 208170 500754 208226
rect 500810 208170 500878 208226
rect 500934 208170 501002 208226
rect 501058 208170 501126 208226
rect 501182 208170 531474 208226
rect 531530 208170 531598 208226
rect 531654 208170 531722 208226
rect 531778 208170 531846 208226
rect 531902 208170 562194 208226
rect 562250 208170 562318 208226
rect 562374 208170 562442 208226
rect 562498 208170 562566 208226
rect 562622 208170 592914 208226
rect 592970 208170 593038 208226
rect 593094 208170 593162 208226
rect 593218 208170 593286 208226
rect 593342 208170 597456 208226
rect 597512 208170 597580 208226
rect 597636 208170 597704 208226
rect 597760 208170 597828 208226
rect 597884 208170 597980 208226
rect -1916 208102 597980 208170
rect -1916 208046 -1820 208102
rect -1764 208046 -1696 208102
rect -1640 208046 -1572 208102
rect -1516 208046 -1448 208102
rect -1392 208046 9234 208102
rect 9290 208046 9358 208102
rect 9414 208046 9482 208102
rect 9538 208046 9606 208102
rect 9662 208046 39954 208102
rect 40010 208046 40078 208102
rect 40134 208046 40202 208102
rect 40258 208046 40326 208102
rect 40382 208046 70674 208102
rect 70730 208046 70798 208102
rect 70854 208046 70922 208102
rect 70978 208046 71046 208102
rect 71102 208046 101394 208102
rect 101450 208046 101518 208102
rect 101574 208046 101642 208102
rect 101698 208046 101766 208102
rect 101822 208046 132114 208102
rect 132170 208046 132238 208102
rect 132294 208046 132362 208102
rect 132418 208046 132486 208102
rect 132542 208046 162834 208102
rect 162890 208046 162958 208102
rect 163014 208046 163082 208102
rect 163138 208046 163206 208102
rect 163262 208046 193554 208102
rect 193610 208046 193678 208102
rect 193734 208046 193802 208102
rect 193858 208046 193926 208102
rect 193982 208046 224274 208102
rect 224330 208046 224398 208102
rect 224454 208046 224522 208102
rect 224578 208046 224646 208102
rect 224702 208046 254994 208102
rect 255050 208046 255118 208102
rect 255174 208046 255242 208102
rect 255298 208046 255366 208102
rect 255422 208046 285714 208102
rect 285770 208046 285838 208102
rect 285894 208046 285962 208102
rect 286018 208046 286086 208102
rect 286142 208046 316434 208102
rect 316490 208046 316558 208102
rect 316614 208046 316682 208102
rect 316738 208046 316806 208102
rect 316862 208046 347154 208102
rect 347210 208046 347278 208102
rect 347334 208046 347402 208102
rect 347458 208046 347526 208102
rect 347582 208046 377874 208102
rect 377930 208046 377998 208102
rect 378054 208046 378122 208102
rect 378178 208046 378246 208102
rect 378302 208046 408594 208102
rect 408650 208046 408718 208102
rect 408774 208046 408842 208102
rect 408898 208046 408966 208102
rect 409022 208046 439314 208102
rect 439370 208046 439438 208102
rect 439494 208046 439562 208102
rect 439618 208046 439686 208102
rect 439742 208046 470034 208102
rect 470090 208046 470158 208102
rect 470214 208046 470282 208102
rect 470338 208046 470406 208102
rect 470462 208046 500754 208102
rect 500810 208046 500878 208102
rect 500934 208046 501002 208102
rect 501058 208046 501126 208102
rect 501182 208046 531474 208102
rect 531530 208046 531598 208102
rect 531654 208046 531722 208102
rect 531778 208046 531846 208102
rect 531902 208046 562194 208102
rect 562250 208046 562318 208102
rect 562374 208046 562442 208102
rect 562498 208046 562566 208102
rect 562622 208046 592914 208102
rect 592970 208046 593038 208102
rect 593094 208046 593162 208102
rect 593218 208046 593286 208102
rect 593342 208046 597456 208102
rect 597512 208046 597580 208102
rect 597636 208046 597704 208102
rect 597760 208046 597828 208102
rect 597884 208046 597980 208102
rect -1916 207978 597980 208046
rect -1916 207922 -1820 207978
rect -1764 207922 -1696 207978
rect -1640 207922 -1572 207978
rect -1516 207922 -1448 207978
rect -1392 207922 9234 207978
rect 9290 207922 9358 207978
rect 9414 207922 9482 207978
rect 9538 207922 9606 207978
rect 9662 207922 39954 207978
rect 40010 207922 40078 207978
rect 40134 207922 40202 207978
rect 40258 207922 40326 207978
rect 40382 207922 70674 207978
rect 70730 207922 70798 207978
rect 70854 207922 70922 207978
rect 70978 207922 71046 207978
rect 71102 207922 101394 207978
rect 101450 207922 101518 207978
rect 101574 207922 101642 207978
rect 101698 207922 101766 207978
rect 101822 207922 132114 207978
rect 132170 207922 132238 207978
rect 132294 207922 132362 207978
rect 132418 207922 132486 207978
rect 132542 207922 162834 207978
rect 162890 207922 162958 207978
rect 163014 207922 163082 207978
rect 163138 207922 163206 207978
rect 163262 207922 193554 207978
rect 193610 207922 193678 207978
rect 193734 207922 193802 207978
rect 193858 207922 193926 207978
rect 193982 207922 224274 207978
rect 224330 207922 224398 207978
rect 224454 207922 224522 207978
rect 224578 207922 224646 207978
rect 224702 207922 254994 207978
rect 255050 207922 255118 207978
rect 255174 207922 255242 207978
rect 255298 207922 255366 207978
rect 255422 207922 285714 207978
rect 285770 207922 285838 207978
rect 285894 207922 285962 207978
rect 286018 207922 286086 207978
rect 286142 207922 316434 207978
rect 316490 207922 316558 207978
rect 316614 207922 316682 207978
rect 316738 207922 316806 207978
rect 316862 207922 347154 207978
rect 347210 207922 347278 207978
rect 347334 207922 347402 207978
rect 347458 207922 347526 207978
rect 347582 207922 377874 207978
rect 377930 207922 377998 207978
rect 378054 207922 378122 207978
rect 378178 207922 378246 207978
rect 378302 207922 408594 207978
rect 408650 207922 408718 207978
rect 408774 207922 408842 207978
rect 408898 207922 408966 207978
rect 409022 207922 439314 207978
rect 439370 207922 439438 207978
rect 439494 207922 439562 207978
rect 439618 207922 439686 207978
rect 439742 207922 470034 207978
rect 470090 207922 470158 207978
rect 470214 207922 470282 207978
rect 470338 207922 470406 207978
rect 470462 207922 500754 207978
rect 500810 207922 500878 207978
rect 500934 207922 501002 207978
rect 501058 207922 501126 207978
rect 501182 207922 531474 207978
rect 531530 207922 531598 207978
rect 531654 207922 531722 207978
rect 531778 207922 531846 207978
rect 531902 207922 562194 207978
rect 562250 207922 562318 207978
rect 562374 207922 562442 207978
rect 562498 207922 562566 207978
rect 562622 207922 592914 207978
rect 592970 207922 593038 207978
rect 593094 207922 593162 207978
rect 593218 207922 593286 207978
rect 593342 207922 597456 207978
rect 597512 207922 597580 207978
rect 597636 207922 597704 207978
rect 597760 207922 597828 207978
rect 597884 207922 597980 207978
rect -1916 207826 597980 207922
rect -1916 202350 597980 202446
rect -1916 202294 -860 202350
rect -804 202294 -736 202350
rect -680 202294 -612 202350
rect -556 202294 -488 202350
rect -432 202294 5514 202350
rect 5570 202294 5638 202350
rect 5694 202294 5762 202350
rect 5818 202294 5886 202350
rect 5942 202294 36234 202350
rect 36290 202294 36358 202350
rect 36414 202294 36482 202350
rect 36538 202294 36606 202350
rect 36662 202294 66954 202350
rect 67010 202294 67078 202350
rect 67134 202294 67202 202350
rect 67258 202294 67326 202350
rect 67382 202294 97674 202350
rect 97730 202294 97798 202350
rect 97854 202294 97922 202350
rect 97978 202294 98046 202350
rect 98102 202294 128394 202350
rect 128450 202294 128518 202350
rect 128574 202294 128642 202350
rect 128698 202294 128766 202350
rect 128822 202294 159114 202350
rect 159170 202294 159238 202350
rect 159294 202294 159362 202350
rect 159418 202294 159486 202350
rect 159542 202294 189834 202350
rect 189890 202294 189958 202350
rect 190014 202294 190082 202350
rect 190138 202294 190206 202350
rect 190262 202294 220554 202350
rect 220610 202294 220678 202350
rect 220734 202294 220802 202350
rect 220858 202294 220926 202350
rect 220982 202294 251274 202350
rect 251330 202294 251398 202350
rect 251454 202294 251522 202350
rect 251578 202294 251646 202350
rect 251702 202294 281994 202350
rect 282050 202294 282118 202350
rect 282174 202294 282242 202350
rect 282298 202294 282366 202350
rect 282422 202294 312714 202350
rect 312770 202294 312838 202350
rect 312894 202294 312962 202350
rect 313018 202294 313086 202350
rect 313142 202294 343434 202350
rect 343490 202294 343558 202350
rect 343614 202294 343682 202350
rect 343738 202294 343806 202350
rect 343862 202294 374154 202350
rect 374210 202294 374278 202350
rect 374334 202294 374402 202350
rect 374458 202294 374526 202350
rect 374582 202294 404874 202350
rect 404930 202294 404998 202350
rect 405054 202294 405122 202350
rect 405178 202294 405246 202350
rect 405302 202294 435594 202350
rect 435650 202294 435718 202350
rect 435774 202294 435842 202350
rect 435898 202294 435966 202350
rect 436022 202294 466314 202350
rect 466370 202294 466438 202350
rect 466494 202294 466562 202350
rect 466618 202294 466686 202350
rect 466742 202294 497034 202350
rect 497090 202294 497158 202350
rect 497214 202294 497282 202350
rect 497338 202294 497406 202350
rect 497462 202294 527754 202350
rect 527810 202294 527878 202350
rect 527934 202294 528002 202350
rect 528058 202294 528126 202350
rect 528182 202294 558474 202350
rect 558530 202294 558598 202350
rect 558654 202294 558722 202350
rect 558778 202294 558846 202350
rect 558902 202294 589194 202350
rect 589250 202294 589318 202350
rect 589374 202294 589442 202350
rect 589498 202294 589566 202350
rect 589622 202294 596496 202350
rect 596552 202294 596620 202350
rect 596676 202294 596744 202350
rect 596800 202294 596868 202350
rect 596924 202294 597980 202350
rect -1916 202226 597980 202294
rect -1916 202170 -860 202226
rect -804 202170 -736 202226
rect -680 202170 -612 202226
rect -556 202170 -488 202226
rect -432 202170 5514 202226
rect 5570 202170 5638 202226
rect 5694 202170 5762 202226
rect 5818 202170 5886 202226
rect 5942 202170 36234 202226
rect 36290 202170 36358 202226
rect 36414 202170 36482 202226
rect 36538 202170 36606 202226
rect 36662 202170 66954 202226
rect 67010 202170 67078 202226
rect 67134 202170 67202 202226
rect 67258 202170 67326 202226
rect 67382 202170 97674 202226
rect 97730 202170 97798 202226
rect 97854 202170 97922 202226
rect 97978 202170 98046 202226
rect 98102 202170 128394 202226
rect 128450 202170 128518 202226
rect 128574 202170 128642 202226
rect 128698 202170 128766 202226
rect 128822 202170 159114 202226
rect 159170 202170 159238 202226
rect 159294 202170 159362 202226
rect 159418 202170 159486 202226
rect 159542 202170 189834 202226
rect 189890 202170 189958 202226
rect 190014 202170 190082 202226
rect 190138 202170 190206 202226
rect 190262 202170 220554 202226
rect 220610 202170 220678 202226
rect 220734 202170 220802 202226
rect 220858 202170 220926 202226
rect 220982 202170 251274 202226
rect 251330 202170 251398 202226
rect 251454 202170 251522 202226
rect 251578 202170 251646 202226
rect 251702 202170 281994 202226
rect 282050 202170 282118 202226
rect 282174 202170 282242 202226
rect 282298 202170 282366 202226
rect 282422 202170 312714 202226
rect 312770 202170 312838 202226
rect 312894 202170 312962 202226
rect 313018 202170 313086 202226
rect 313142 202170 343434 202226
rect 343490 202170 343558 202226
rect 343614 202170 343682 202226
rect 343738 202170 343806 202226
rect 343862 202170 374154 202226
rect 374210 202170 374278 202226
rect 374334 202170 374402 202226
rect 374458 202170 374526 202226
rect 374582 202170 404874 202226
rect 404930 202170 404998 202226
rect 405054 202170 405122 202226
rect 405178 202170 405246 202226
rect 405302 202170 435594 202226
rect 435650 202170 435718 202226
rect 435774 202170 435842 202226
rect 435898 202170 435966 202226
rect 436022 202170 466314 202226
rect 466370 202170 466438 202226
rect 466494 202170 466562 202226
rect 466618 202170 466686 202226
rect 466742 202170 497034 202226
rect 497090 202170 497158 202226
rect 497214 202170 497282 202226
rect 497338 202170 497406 202226
rect 497462 202170 527754 202226
rect 527810 202170 527878 202226
rect 527934 202170 528002 202226
rect 528058 202170 528126 202226
rect 528182 202170 558474 202226
rect 558530 202170 558598 202226
rect 558654 202170 558722 202226
rect 558778 202170 558846 202226
rect 558902 202170 589194 202226
rect 589250 202170 589318 202226
rect 589374 202170 589442 202226
rect 589498 202170 589566 202226
rect 589622 202170 596496 202226
rect 596552 202170 596620 202226
rect 596676 202170 596744 202226
rect 596800 202170 596868 202226
rect 596924 202170 597980 202226
rect -1916 202102 597980 202170
rect -1916 202046 -860 202102
rect -804 202046 -736 202102
rect -680 202046 -612 202102
rect -556 202046 -488 202102
rect -432 202046 5514 202102
rect 5570 202046 5638 202102
rect 5694 202046 5762 202102
rect 5818 202046 5886 202102
rect 5942 202046 36234 202102
rect 36290 202046 36358 202102
rect 36414 202046 36482 202102
rect 36538 202046 36606 202102
rect 36662 202046 66954 202102
rect 67010 202046 67078 202102
rect 67134 202046 67202 202102
rect 67258 202046 67326 202102
rect 67382 202046 97674 202102
rect 97730 202046 97798 202102
rect 97854 202046 97922 202102
rect 97978 202046 98046 202102
rect 98102 202046 128394 202102
rect 128450 202046 128518 202102
rect 128574 202046 128642 202102
rect 128698 202046 128766 202102
rect 128822 202046 159114 202102
rect 159170 202046 159238 202102
rect 159294 202046 159362 202102
rect 159418 202046 159486 202102
rect 159542 202046 189834 202102
rect 189890 202046 189958 202102
rect 190014 202046 190082 202102
rect 190138 202046 190206 202102
rect 190262 202046 220554 202102
rect 220610 202046 220678 202102
rect 220734 202046 220802 202102
rect 220858 202046 220926 202102
rect 220982 202046 251274 202102
rect 251330 202046 251398 202102
rect 251454 202046 251522 202102
rect 251578 202046 251646 202102
rect 251702 202046 281994 202102
rect 282050 202046 282118 202102
rect 282174 202046 282242 202102
rect 282298 202046 282366 202102
rect 282422 202046 312714 202102
rect 312770 202046 312838 202102
rect 312894 202046 312962 202102
rect 313018 202046 313086 202102
rect 313142 202046 343434 202102
rect 343490 202046 343558 202102
rect 343614 202046 343682 202102
rect 343738 202046 343806 202102
rect 343862 202046 374154 202102
rect 374210 202046 374278 202102
rect 374334 202046 374402 202102
rect 374458 202046 374526 202102
rect 374582 202046 404874 202102
rect 404930 202046 404998 202102
rect 405054 202046 405122 202102
rect 405178 202046 405246 202102
rect 405302 202046 435594 202102
rect 435650 202046 435718 202102
rect 435774 202046 435842 202102
rect 435898 202046 435966 202102
rect 436022 202046 466314 202102
rect 466370 202046 466438 202102
rect 466494 202046 466562 202102
rect 466618 202046 466686 202102
rect 466742 202046 497034 202102
rect 497090 202046 497158 202102
rect 497214 202046 497282 202102
rect 497338 202046 497406 202102
rect 497462 202046 527754 202102
rect 527810 202046 527878 202102
rect 527934 202046 528002 202102
rect 528058 202046 528126 202102
rect 528182 202046 558474 202102
rect 558530 202046 558598 202102
rect 558654 202046 558722 202102
rect 558778 202046 558846 202102
rect 558902 202046 589194 202102
rect 589250 202046 589318 202102
rect 589374 202046 589442 202102
rect 589498 202046 589566 202102
rect 589622 202046 596496 202102
rect 596552 202046 596620 202102
rect 596676 202046 596744 202102
rect 596800 202046 596868 202102
rect 596924 202046 597980 202102
rect -1916 201978 597980 202046
rect -1916 201922 -860 201978
rect -804 201922 -736 201978
rect -680 201922 -612 201978
rect -556 201922 -488 201978
rect -432 201922 5514 201978
rect 5570 201922 5638 201978
rect 5694 201922 5762 201978
rect 5818 201922 5886 201978
rect 5942 201922 36234 201978
rect 36290 201922 36358 201978
rect 36414 201922 36482 201978
rect 36538 201922 36606 201978
rect 36662 201922 66954 201978
rect 67010 201922 67078 201978
rect 67134 201922 67202 201978
rect 67258 201922 67326 201978
rect 67382 201922 97674 201978
rect 97730 201922 97798 201978
rect 97854 201922 97922 201978
rect 97978 201922 98046 201978
rect 98102 201922 128394 201978
rect 128450 201922 128518 201978
rect 128574 201922 128642 201978
rect 128698 201922 128766 201978
rect 128822 201922 159114 201978
rect 159170 201922 159238 201978
rect 159294 201922 159362 201978
rect 159418 201922 159486 201978
rect 159542 201922 189834 201978
rect 189890 201922 189958 201978
rect 190014 201922 190082 201978
rect 190138 201922 190206 201978
rect 190262 201922 220554 201978
rect 220610 201922 220678 201978
rect 220734 201922 220802 201978
rect 220858 201922 220926 201978
rect 220982 201922 251274 201978
rect 251330 201922 251398 201978
rect 251454 201922 251522 201978
rect 251578 201922 251646 201978
rect 251702 201922 281994 201978
rect 282050 201922 282118 201978
rect 282174 201922 282242 201978
rect 282298 201922 282366 201978
rect 282422 201922 312714 201978
rect 312770 201922 312838 201978
rect 312894 201922 312962 201978
rect 313018 201922 313086 201978
rect 313142 201922 343434 201978
rect 343490 201922 343558 201978
rect 343614 201922 343682 201978
rect 343738 201922 343806 201978
rect 343862 201922 374154 201978
rect 374210 201922 374278 201978
rect 374334 201922 374402 201978
rect 374458 201922 374526 201978
rect 374582 201922 404874 201978
rect 404930 201922 404998 201978
rect 405054 201922 405122 201978
rect 405178 201922 405246 201978
rect 405302 201922 435594 201978
rect 435650 201922 435718 201978
rect 435774 201922 435842 201978
rect 435898 201922 435966 201978
rect 436022 201922 466314 201978
rect 466370 201922 466438 201978
rect 466494 201922 466562 201978
rect 466618 201922 466686 201978
rect 466742 201922 497034 201978
rect 497090 201922 497158 201978
rect 497214 201922 497282 201978
rect 497338 201922 497406 201978
rect 497462 201922 527754 201978
rect 527810 201922 527878 201978
rect 527934 201922 528002 201978
rect 528058 201922 528126 201978
rect 528182 201922 558474 201978
rect 558530 201922 558598 201978
rect 558654 201922 558722 201978
rect 558778 201922 558846 201978
rect 558902 201922 589194 201978
rect 589250 201922 589318 201978
rect 589374 201922 589442 201978
rect 589498 201922 589566 201978
rect 589622 201922 596496 201978
rect 596552 201922 596620 201978
rect 596676 201922 596744 201978
rect 596800 201922 596868 201978
rect 596924 201922 597980 201978
rect -1916 201826 597980 201922
rect -1916 190350 597980 190446
rect -1916 190294 -1820 190350
rect -1764 190294 -1696 190350
rect -1640 190294 -1572 190350
rect -1516 190294 -1448 190350
rect -1392 190294 9234 190350
rect 9290 190294 9358 190350
rect 9414 190294 9482 190350
rect 9538 190294 9606 190350
rect 9662 190294 39954 190350
rect 40010 190294 40078 190350
rect 40134 190294 40202 190350
rect 40258 190294 40326 190350
rect 40382 190294 70674 190350
rect 70730 190294 70798 190350
rect 70854 190294 70922 190350
rect 70978 190294 71046 190350
rect 71102 190294 101394 190350
rect 101450 190294 101518 190350
rect 101574 190294 101642 190350
rect 101698 190294 101766 190350
rect 101822 190294 132114 190350
rect 132170 190294 132238 190350
rect 132294 190294 132362 190350
rect 132418 190294 132486 190350
rect 132542 190294 162834 190350
rect 162890 190294 162958 190350
rect 163014 190294 163082 190350
rect 163138 190294 163206 190350
rect 163262 190294 193554 190350
rect 193610 190294 193678 190350
rect 193734 190294 193802 190350
rect 193858 190294 193926 190350
rect 193982 190294 224274 190350
rect 224330 190294 224398 190350
rect 224454 190294 224522 190350
rect 224578 190294 224646 190350
rect 224702 190294 254994 190350
rect 255050 190294 255118 190350
rect 255174 190294 255242 190350
rect 255298 190294 255366 190350
rect 255422 190294 285714 190350
rect 285770 190294 285838 190350
rect 285894 190294 285962 190350
rect 286018 190294 286086 190350
rect 286142 190294 316434 190350
rect 316490 190294 316558 190350
rect 316614 190294 316682 190350
rect 316738 190294 316806 190350
rect 316862 190294 347154 190350
rect 347210 190294 347278 190350
rect 347334 190294 347402 190350
rect 347458 190294 347526 190350
rect 347582 190294 377874 190350
rect 377930 190294 377998 190350
rect 378054 190294 378122 190350
rect 378178 190294 378246 190350
rect 378302 190294 408594 190350
rect 408650 190294 408718 190350
rect 408774 190294 408842 190350
rect 408898 190294 408966 190350
rect 409022 190294 439314 190350
rect 439370 190294 439438 190350
rect 439494 190294 439562 190350
rect 439618 190294 439686 190350
rect 439742 190294 470034 190350
rect 470090 190294 470158 190350
rect 470214 190294 470282 190350
rect 470338 190294 470406 190350
rect 470462 190294 500754 190350
rect 500810 190294 500878 190350
rect 500934 190294 501002 190350
rect 501058 190294 501126 190350
rect 501182 190294 531474 190350
rect 531530 190294 531598 190350
rect 531654 190294 531722 190350
rect 531778 190294 531846 190350
rect 531902 190294 562194 190350
rect 562250 190294 562318 190350
rect 562374 190294 562442 190350
rect 562498 190294 562566 190350
rect 562622 190294 592914 190350
rect 592970 190294 593038 190350
rect 593094 190294 593162 190350
rect 593218 190294 593286 190350
rect 593342 190294 597456 190350
rect 597512 190294 597580 190350
rect 597636 190294 597704 190350
rect 597760 190294 597828 190350
rect 597884 190294 597980 190350
rect -1916 190226 597980 190294
rect -1916 190170 -1820 190226
rect -1764 190170 -1696 190226
rect -1640 190170 -1572 190226
rect -1516 190170 -1448 190226
rect -1392 190170 9234 190226
rect 9290 190170 9358 190226
rect 9414 190170 9482 190226
rect 9538 190170 9606 190226
rect 9662 190170 39954 190226
rect 40010 190170 40078 190226
rect 40134 190170 40202 190226
rect 40258 190170 40326 190226
rect 40382 190170 70674 190226
rect 70730 190170 70798 190226
rect 70854 190170 70922 190226
rect 70978 190170 71046 190226
rect 71102 190170 101394 190226
rect 101450 190170 101518 190226
rect 101574 190170 101642 190226
rect 101698 190170 101766 190226
rect 101822 190170 132114 190226
rect 132170 190170 132238 190226
rect 132294 190170 132362 190226
rect 132418 190170 132486 190226
rect 132542 190170 162834 190226
rect 162890 190170 162958 190226
rect 163014 190170 163082 190226
rect 163138 190170 163206 190226
rect 163262 190170 193554 190226
rect 193610 190170 193678 190226
rect 193734 190170 193802 190226
rect 193858 190170 193926 190226
rect 193982 190170 224274 190226
rect 224330 190170 224398 190226
rect 224454 190170 224522 190226
rect 224578 190170 224646 190226
rect 224702 190170 254994 190226
rect 255050 190170 255118 190226
rect 255174 190170 255242 190226
rect 255298 190170 255366 190226
rect 255422 190170 285714 190226
rect 285770 190170 285838 190226
rect 285894 190170 285962 190226
rect 286018 190170 286086 190226
rect 286142 190170 316434 190226
rect 316490 190170 316558 190226
rect 316614 190170 316682 190226
rect 316738 190170 316806 190226
rect 316862 190170 347154 190226
rect 347210 190170 347278 190226
rect 347334 190170 347402 190226
rect 347458 190170 347526 190226
rect 347582 190170 377874 190226
rect 377930 190170 377998 190226
rect 378054 190170 378122 190226
rect 378178 190170 378246 190226
rect 378302 190170 408594 190226
rect 408650 190170 408718 190226
rect 408774 190170 408842 190226
rect 408898 190170 408966 190226
rect 409022 190170 439314 190226
rect 439370 190170 439438 190226
rect 439494 190170 439562 190226
rect 439618 190170 439686 190226
rect 439742 190170 470034 190226
rect 470090 190170 470158 190226
rect 470214 190170 470282 190226
rect 470338 190170 470406 190226
rect 470462 190170 500754 190226
rect 500810 190170 500878 190226
rect 500934 190170 501002 190226
rect 501058 190170 501126 190226
rect 501182 190170 531474 190226
rect 531530 190170 531598 190226
rect 531654 190170 531722 190226
rect 531778 190170 531846 190226
rect 531902 190170 562194 190226
rect 562250 190170 562318 190226
rect 562374 190170 562442 190226
rect 562498 190170 562566 190226
rect 562622 190170 592914 190226
rect 592970 190170 593038 190226
rect 593094 190170 593162 190226
rect 593218 190170 593286 190226
rect 593342 190170 597456 190226
rect 597512 190170 597580 190226
rect 597636 190170 597704 190226
rect 597760 190170 597828 190226
rect 597884 190170 597980 190226
rect -1916 190102 597980 190170
rect -1916 190046 -1820 190102
rect -1764 190046 -1696 190102
rect -1640 190046 -1572 190102
rect -1516 190046 -1448 190102
rect -1392 190046 9234 190102
rect 9290 190046 9358 190102
rect 9414 190046 9482 190102
rect 9538 190046 9606 190102
rect 9662 190046 39954 190102
rect 40010 190046 40078 190102
rect 40134 190046 40202 190102
rect 40258 190046 40326 190102
rect 40382 190046 70674 190102
rect 70730 190046 70798 190102
rect 70854 190046 70922 190102
rect 70978 190046 71046 190102
rect 71102 190046 101394 190102
rect 101450 190046 101518 190102
rect 101574 190046 101642 190102
rect 101698 190046 101766 190102
rect 101822 190046 132114 190102
rect 132170 190046 132238 190102
rect 132294 190046 132362 190102
rect 132418 190046 132486 190102
rect 132542 190046 162834 190102
rect 162890 190046 162958 190102
rect 163014 190046 163082 190102
rect 163138 190046 163206 190102
rect 163262 190046 193554 190102
rect 193610 190046 193678 190102
rect 193734 190046 193802 190102
rect 193858 190046 193926 190102
rect 193982 190046 224274 190102
rect 224330 190046 224398 190102
rect 224454 190046 224522 190102
rect 224578 190046 224646 190102
rect 224702 190046 254994 190102
rect 255050 190046 255118 190102
rect 255174 190046 255242 190102
rect 255298 190046 255366 190102
rect 255422 190046 285714 190102
rect 285770 190046 285838 190102
rect 285894 190046 285962 190102
rect 286018 190046 286086 190102
rect 286142 190046 316434 190102
rect 316490 190046 316558 190102
rect 316614 190046 316682 190102
rect 316738 190046 316806 190102
rect 316862 190046 347154 190102
rect 347210 190046 347278 190102
rect 347334 190046 347402 190102
rect 347458 190046 347526 190102
rect 347582 190046 377874 190102
rect 377930 190046 377998 190102
rect 378054 190046 378122 190102
rect 378178 190046 378246 190102
rect 378302 190046 408594 190102
rect 408650 190046 408718 190102
rect 408774 190046 408842 190102
rect 408898 190046 408966 190102
rect 409022 190046 439314 190102
rect 439370 190046 439438 190102
rect 439494 190046 439562 190102
rect 439618 190046 439686 190102
rect 439742 190046 470034 190102
rect 470090 190046 470158 190102
rect 470214 190046 470282 190102
rect 470338 190046 470406 190102
rect 470462 190046 500754 190102
rect 500810 190046 500878 190102
rect 500934 190046 501002 190102
rect 501058 190046 501126 190102
rect 501182 190046 531474 190102
rect 531530 190046 531598 190102
rect 531654 190046 531722 190102
rect 531778 190046 531846 190102
rect 531902 190046 562194 190102
rect 562250 190046 562318 190102
rect 562374 190046 562442 190102
rect 562498 190046 562566 190102
rect 562622 190046 592914 190102
rect 592970 190046 593038 190102
rect 593094 190046 593162 190102
rect 593218 190046 593286 190102
rect 593342 190046 597456 190102
rect 597512 190046 597580 190102
rect 597636 190046 597704 190102
rect 597760 190046 597828 190102
rect 597884 190046 597980 190102
rect -1916 189978 597980 190046
rect -1916 189922 -1820 189978
rect -1764 189922 -1696 189978
rect -1640 189922 -1572 189978
rect -1516 189922 -1448 189978
rect -1392 189922 9234 189978
rect 9290 189922 9358 189978
rect 9414 189922 9482 189978
rect 9538 189922 9606 189978
rect 9662 189922 39954 189978
rect 40010 189922 40078 189978
rect 40134 189922 40202 189978
rect 40258 189922 40326 189978
rect 40382 189922 70674 189978
rect 70730 189922 70798 189978
rect 70854 189922 70922 189978
rect 70978 189922 71046 189978
rect 71102 189922 101394 189978
rect 101450 189922 101518 189978
rect 101574 189922 101642 189978
rect 101698 189922 101766 189978
rect 101822 189922 132114 189978
rect 132170 189922 132238 189978
rect 132294 189922 132362 189978
rect 132418 189922 132486 189978
rect 132542 189922 162834 189978
rect 162890 189922 162958 189978
rect 163014 189922 163082 189978
rect 163138 189922 163206 189978
rect 163262 189922 193554 189978
rect 193610 189922 193678 189978
rect 193734 189922 193802 189978
rect 193858 189922 193926 189978
rect 193982 189922 224274 189978
rect 224330 189922 224398 189978
rect 224454 189922 224522 189978
rect 224578 189922 224646 189978
rect 224702 189922 254994 189978
rect 255050 189922 255118 189978
rect 255174 189922 255242 189978
rect 255298 189922 255366 189978
rect 255422 189922 285714 189978
rect 285770 189922 285838 189978
rect 285894 189922 285962 189978
rect 286018 189922 286086 189978
rect 286142 189922 316434 189978
rect 316490 189922 316558 189978
rect 316614 189922 316682 189978
rect 316738 189922 316806 189978
rect 316862 189922 347154 189978
rect 347210 189922 347278 189978
rect 347334 189922 347402 189978
rect 347458 189922 347526 189978
rect 347582 189922 377874 189978
rect 377930 189922 377998 189978
rect 378054 189922 378122 189978
rect 378178 189922 378246 189978
rect 378302 189922 408594 189978
rect 408650 189922 408718 189978
rect 408774 189922 408842 189978
rect 408898 189922 408966 189978
rect 409022 189922 439314 189978
rect 439370 189922 439438 189978
rect 439494 189922 439562 189978
rect 439618 189922 439686 189978
rect 439742 189922 470034 189978
rect 470090 189922 470158 189978
rect 470214 189922 470282 189978
rect 470338 189922 470406 189978
rect 470462 189922 500754 189978
rect 500810 189922 500878 189978
rect 500934 189922 501002 189978
rect 501058 189922 501126 189978
rect 501182 189922 531474 189978
rect 531530 189922 531598 189978
rect 531654 189922 531722 189978
rect 531778 189922 531846 189978
rect 531902 189922 562194 189978
rect 562250 189922 562318 189978
rect 562374 189922 562442 189978
rect 562498 189922 562566 189978
rect 562622 189922 592914 189978
rect 592970 189922 593038 189978
rect 593094 189922 593162 189978
rect 593218 189922 593286 189978
rect 593342 189922 597456 189978
rect 597512 189922 597580 189978
rect 597636 189922 597704 189978
rect 597760 189922 597828 189978
rect 597884 189922 597980 189978
rect -1916 189826 597980 189922
rect -1916 184350 597980 184446
rect -1916 184294 -860 184350
rect -804 184294 -736 184350
rect -680 184294 -612 184350
rect -556 184294 -488 184350
rect -432 184294 5514 184350
rect 5570 184294 5638 184350
rect 5694 184294 5762 184350
rect 5818 184294 5886 184350
rect 5942 184294 36234 184350
rect 36290 184294 36358 184350
rect 36414 184294 36482 184350
rect 36538 184294 36606 184350
rect 36662 184294 66954 184350
rect 67010 184294 67078 184350
rect 67134 184294 67202 184350
rect 67258 184294 67326 184350
rect 67382 184294 97674 184350
rect 97730 184294 97798 184350
rect 97854 184294 97922 184350
rect 97978 184294 98046 184350
rect 98102 184294 128394 184350
rect 128450 184294 128518 184350
rect 128574 184294 128642 184350
rect 128698 184294 128766 184350
rect 128822 184294 159114 184350
rect 159170 184294 159238 184350
rect 159294 184294 159362 184350
rect 159418 184294 159486 184350
rect 159542 184294 189834 184350
rect 189890 184294 189958 184350
rect 190014 184294 190082 184350
rect 190138 184294 190206 184350
rect 190262 184294 220554 184350
rect 220610 184294 220678 184350
rect 220734 184294 220802 184350
rect 220858 184294 220926 184350
rect 220982 184294 251274 184350
rect 251330 184294 251398 184350
rect 251454 184294 251522 184350
rect 251578 184294 251646 184350
rect 251702 184294 281994 184350
rect 282050 184294 282118 184350
rect 282174 184294 282242 184350
rect 282298 184294 282366 184350
rect 282422 184294 312714 184350
rect 312770 184294 312838 184350
rect 312894 184294 312962 184350
rect 313018 184294 313086 184350
rect 313142 184294 343434 184350
rect 343490 184294 343558 184350
rect 343614 184294 343682 184350
rect 343738 184294 343806 184350
rect 343862 184294 374154 184350
rect 374210 184294 374278 184350
rect 374334 184294 374402 184350
rect 374458 184294 374526 184350
rect 374582 184294 404874 184350
rect 404930 184294 404998 184350
rect 405054 184294 405122 184350
rect 405178 184294 405246 184350
rect 405302 184294 435594 184350
rect 435650 184294 435718 184350
rect 435774 184294 435842 184350
rect 435898 184294 435966 184350
rect 436022 184294 466314 184350
rect 466370 184294 466438 184350
rect 466494 184294 466562 184350
rect 466618 184294 466686 184350
rect 466742 184294 497034 184350
rect 497090 184294 497158 184350
rect 497214 184294 497282 184350
rect 497338 184294 497406 184350
rect 497462 184294 527754 184350
rect 527810 184294 527878 184350
rect 527934 184294 528002 184350
rect 528058 184294 528126 184350
rect 528182 184294 558474 184350
rect 558530 184294 558598 184350
rect 558654 184294 558722 184350
rect 558778 184294 558846 184350
rect 558902 184294 589194 184350
rect 589250 184294 589318 184350
rect 589374 184294 589442 184350
rect 589498 184294 589566 184350
rect 589622 184294 596496 184350
rect 596552 184294 596620 184350
rect 596676 184294 596744 184350
rect 596800 184294 596868 184350
rect 596924 184294 597980 184350
rect -1916 184226 597980 184294
rect -1916 184170 -860 184226
rect -804 184170 -736 184226
rect -680 184170 -612 184226
rect -556 184170 -488 184226
rect -432 184170 5514 184226
rect 5570 184170 5638 184226
rect 5694 184170 5762 184226
rect 5818 184170 5886 184226
rect 5942 184170 36234 184226
rect 36290 184170 36358 184226
rect 36414 184170 36482 184226
rect 36538 184170 36606 184226
rect 36662 184170 66954 184226
rect 67010 184170 67078 184226
rect 67134 184170 67202 184226
rect 67258 184170 67326 184226
rect 67382 184170 97674 184226
rect 97730 184170 97798 184226
rect 97854 184170 97922 184226
rect 97978 184170 98046 184226
rect 98102 184170 128394 184226
rect 128450 184170 128518 184226
rect 128574 184170 128642 184226
rect 128698 184170 128766 184226
rect 128822 184170 159114 184226
rect 159170 184170 159238 184226
rect 159294 184170 159362 184226
rect 159418 184170 159486 184226
rect 159542 184170 189834 184226
rect 189890 184170 189958 184226
rect 190014 184170 190082 184226
rect 190138 184170 190206 184226
rect 190262 184170 220554 184226
rect 220610 184170 220678 184226
rect 220734 184170 220802 184226
rect 220858 184170 220926 184226
rect 220982 184170 251274 184226
rect 251330 184170 251398 184226
rect 251454 184170 251522 184226
rect 251578 184170 251646 184226
rect 251702 184170 281994 184226
rect 282050 184170 282118 184226
rect 282174 184170 282242 184226
rect 282298 184170 282366 184226
rect 282422 184170 312714 184226
rect 312770 184170 312838 184226
rect 312894 184170 312962 184226
rect 313018 184170 313086 184226
rect 313142 184170 343434 184226
rect 343490 184170 343558 184226
rect 343614 184170 343682 184226
rect 343738 184170 343806 184226
rect 343862 184170 374154 184226
rect 374210 184170 374278 184226
rect 374334 184170 374402 184226
rect 374458 184170 374526 184226
rect 374582 184170 404874 184226
rect 404930 184170 404998 184226
rect 405054 184170 405122 184226
rect 405178 184170 405246 184226
rect 405302 184170 435594 184226
rect 435650 184170 435718 184226
rect 435774 184170 435842 184226
rect 435898 184170 435966 184226
rect 436022 184170 466314 184226
rect 466370 184170 466438 184226
rect 466494 184170 466562 184226
rect 466618 184170 466686 184226
rect 466742 184170 497034 184226
rect 497090 184170 497158 184226
rect 497214 184170 497282 184226
rect 497338 184170 497406 184226
rect 497462 184170 527754 184226
rect 527810 184170 527878 184226
rect 527934 184170 528002 184226
rect 528058 184170 528126 184226
rect 528182 184170 558474 184226
rect 558530 184170 558598 184226
rect 558654 184170 558722 184226
rect 558778 184170 558846 184226
rect 558902 184170 589194 184226
rect 589250 184170 589318 184226
rect 589374 184170 589442 184226
rect 589498 184170 589566 184226
rect 589622 184170 596496 184226
rect 596552 184170 596620 184226
rect 596676 184170 596744 184226
rect 596800 184170 596868 184226
rect 596924 184170 597980 184226
rect -1916 184102 597980 184170
rect -1916 184046 -860 184102
rect -804 184046 -736 184102
rect -680 184046 -612 184102
rect -556 184046 -488 184102
rect -432 184046 5514 184102
rect 5570 184046 5638 184102
rect 5694 184046 5762 184102
rect 5818 184046 5886 184102
rect 5942 184046 36234 184102
rect 36290 184046 36358 184102
rect 36414 184046 36482 184102
rect 36538 184046 36606 184102
rect 36662 184046 66954 184102
rect 67010 184046 67078 184102
rect 67134 184046 67202 184102
rect 67258 184046 67326 184102
rect 67382 184046 97674 184102
rect 97730 184046 97798 184102
rect 97854 184046 97922 184102
rect 97978 184046 98046 184102
rect 98102 184046 128394 184102
rect 128450 184046 128518 184102
rect 128574 184046 128642 184102
rect 128698 184046 128766 184102
rect 128822 184046 159114 184102
rect 159170 184046 159238 184102
rect 159294 184046 159362 184102
rect 159418 184046 159486 184102
rect 159542 184046 189834 184102
rect 189890 184046 189958 184102
rect 190014 184046 190082 184102
rect 190138 184046 190206 184102
rect 190262 184046 220554 184102
rect 220610 184046 220678 184102
rect 220734 184046 220802 184102
rect 220858 184046 220926 184102
rect 220982 184046 251274 184102
rect 251330 184046 251398 184102
rect 251454 184046 251522 184102
rect 251578 184046 251646 184102
rect 251702 184046 281994 184102
rect 282050 184046 282118 184102
rect 282174 184046 282242 184102
rect 282298 184046 282366 184102
rect 282422 184046 312714 184102
rect 312770 184046 312838 184102
rect 312894 184046 312962 184102
rect 313018 184046 313086 184102
rect 313142 184046 343434 184102
rect 343490 184046 343558 184102
rect 343614 184046 343682 184102
rect 343738 184046 343806 184102
rect 343862 184046 374154 184102
rect 374210 184046 374278 184102
rect 374334 184046 374402 184102
rect 374458 184046 374526 184102
rect 374582 184046 404874 184102
rect 404930 184046 404998 184102
rect 405054 184046 405122 184102
rect 405178 184046 405246 184102
rect 405302 184046 435594 184102
rect 435650 184046 435718 184102
rect 435774 184046 435842 184102
rect 435898 184046 435966 184102
rect 436022 184046 466314 184102
rect 466370 184046 466438 184102
rect 466494 184046 466562 184102
rect 466618 184046 466686 184102
rect 466742 184046 497034 184102
rect 497090 184046 497158 184102
rect 497214 184046 497282 184102
rect 497338 184046 497406 184102
rect 497462 184046 527754 184102
rect 527810 184046 527878 184102
rect 527934 184046 528002 184102
rect 528058 184046 528126 184102
rect 528182 184046 558474 184102
rect 558530 184046 558598 184102
rect 558654 184046 558722 184102
rect 558778 184046 558846 184102
rect 558902 184046 589194 184102
rect 589250 184046 589318 184102
rect 589374 184046 589442 184102
rect 589498 184046 589566 184102
rect 589622 184046 596496 184102
rect 596552 184046 596620 184102
rect 596676 184046 596744 184102
rect 596800 184046 596868 184102
rect 596924 184046 597980 184102
rect -1916 183978 597980 184046
rect -1916 183922 -860 183978
rect -804 183922 -736 183978
rect -680 183922 -612 183978
rect -556 183922 -488 183978
rect -432 183922 5514 183978
rect 5570 183922 5638 183978
rect 5694 183922 5762 183978
rect 5818 183922 5886 183978
rect 5942 183922 36234 183978
rect 36290 183922 36358 183978
rect 36414 183922 36482 183978
rect 36538 183922 36606 183978
rect 36662 183922 66954 183978
rect 67010 183922 67078 183978
rect 67134 183922 67202 183978
rect 67258 183922 67326 183978
rect 67382 183922 97674 183978
rect 97730 183922 97798 183978
rect 97854 183922 97922 183978
rect 97978 183922 98046 183978
rect 98102 183922 128394 183978
rect 128450 183922 128518 183978
rect 128574 183922 128642 183978
rect 128698 183922 128766 183978
rect 128822 183922 159114 183978
rect 159170 183922 159238 183978
rect 159294 183922 159362 183978
rect 159418 183922 159486 183978
rect 159542 183922 189834 183978
rect 189890 183922 189958 183978
rect 190014 183922 190082 183978
rect 190138 183922 190206 183978
rect 190262 183922 220554 183978
rect 220610 183922 220678 183978
rect 220734 183922 220802 183978
rect 220858 183922 220926 183978
rect 220982 183922 251274 183978
rect 251330 183922 251398 183978
rect 251454 183922 251522 183978
rect 251578 183922 251646 183978
rect 251702 183922 281994 183978
rect 282050 183922 282118 183978
rect 282174 183922 282242 183978
rect 282298 183922 282366 183978
rect 282422 183922 312714 183978
rect 312770 183922 312838 183978
rect 312894 183922 312962 183978
rect 313018 183922 313086 183978
rect 313142 183922 343434 183978
rect 343490 183922 343558 183978
rect 343614 183922 343682 183978
rect 343738 183922 343806 183978
rect 343862 183922 374154 183978
rect 374210 183922 374278 183978
rect 374334 183922 374402 183978
rect 374458 183922 374526 183978
rect 374582 183922 404874 183978
rect 404930 183922 404998 183978
rect 405054 183922 405122 183978
rect 405178 183922 405246 183978
rect 405302 183922 435594 183978
rect 435650 183922 435718 183978
rect 435774 183922 435842 183978
rect 435898 183922 435966 183978
rect 436022 183922 466314 183978
rect 466370 183922 466438 183978
rect 466494 183922 466562 183978
rect 466618 183922 466686 183978
rect 466742 183922 497034 183978
rect 497090 183922 497158 183978
rect 497214 183922 497282 183978
rect 497338 183922 497406 183978
rect 497462 183922 527754 183978
rect 527810 183922 527878 183978
rect 527934 183922 528002 183978
rect 528058 183922 528126 183978
rect 528182 183922 558474 183978
rect 558530 183922 558598 183978
rect 558654 183922 558722 183978
rect 558778 183922 558846 183978
rect 558902 183922 589194 183978
rect 589250 183922 589318 183978
rect 589374 183922 589442 183978
rect 589498 183922 589566 183978
rect 589622 183922 596496 183978
rect 596552 183922 596620 183978
rect 596676 183922 596744 183978
rect 596800 183922 596868 183978
rect 596924 183922 597980 183978
rect -1916 183826 597980 183922
rect -1916 172350 597980 172446
rect -1916 172294 -1820 172350
rect -1764 172294 -1696 172350
rect -1640 172294 -1572 172350
rect -1516 172294 -1448 172350
rect -1392 172294 9234 172350
rect 9290 172294 9358 172350
rect 9414 172294 9482 172350
rect 9538 172294 9606 172350
rect 9662 172294 39954 172350
rect 40010 172294 40078 172350
rect 40134 172294 40202 172350
rect 40258 172294 40326 172350
rect 40382 172294 70674 172350
rect 70730 172294 70798 172350
rect 70854 172294 70922 172350
rect 70978 172294 71046 172350
rect 71102 172294 101394 172350
rect 101450 172294 101518 172350
rect 101574 172294 101642 172350
rect 101698 172294 101766 172350
rect 101822 172294 132114 172350
rect 132170 172294 132238 172350
rect 132294 172294 132362 172350
rect 132418 172294 132486 172350
rect 132542 172294 162834 172350
rect 162890 172294 162958 172350
rect 163014 172294 163082 172350
rect 163138 172294 163206 172350
rect 163262 172294 193554 172350
rect 193610 172294 193678 172350
rect 193734 172294 193802 172350
rect 193858 172294 193926 172350
rect 193982 172294 224274 172350
rect 224330 172294 224398 172350
rect 224454 172294 224522 172350
rect 224578 172294 224646 172350
rect 224702 172294 254994 172350
rect 255050 172294 255118 172350
rect 255174 172294 255242 172350
rect 255298 172294 255366 172350
rect 255422 172294 285714 172350
rect 285770 172294 285838 172350
rect 285894 172294 285962 172350
rect 286018 172294 286086 172350
rect 286142 172294 316434 172350
rect 316490 172294 316558 172350
rect 316614 172294 316682 172350
rect 316738 172294 316806 172350
rect 316862 172294 347154 172350
rect 347210 172294 347278 172350
rect 347334 172294 347402 172350
rect 347458 172294 347526 172350
rect 347582 172294 377874 172350
rect 377930 172294 377998 172350
rect 378054 172294 378122 172350
rect 378178 172294 378246 172350
rect 378302 172294 408594 172350
rect 408650 172294 408718 172350
rect 408774 172294 408842 172350
rect 408898 172294 408966 172350
rect 409022 172294 439314 172350
rect 439370 172294 439438 172350
rect 439494 172294 439562 172350
rect 439618 172294 439686 172350
rect 439742 172294 470034 172350
rect 470090 172294 470158 172350
rect 470214 172294 470282 172350
rect 470338 172294 470406 172350
rect 470462 172294 500754 172350
rect 500810 172294 500878 172350
rect 500934 172294 501002 172350
rect 501058 172294 501126 172350
rect 501182 172294 531474 172350
rect 531530 172294 531598 172350
rect 531654 172294 531722 172350
rect 531778 172294 531846 172350
rect 531902 172294 562194 172350
rect 562250 172294 562318 172350
rect 562374 172294 562442 172350
rect 562498 172294 562566 172350
rect 562622 172294 592914 172350
rect 592970 172294 593038 172350
rect 593094 172294 593162 172350
rect 593218 172294 593286 172350
rect 593342 172294 597456 172350
rect 597512 172294 597580 172350
rect 597636 172294 597704 172350
rect 597760 172294 597828 172350
rect 597884 172294 597980 172350
rect -1916 172226 597980 172294
rect -1916 172170 -1820 172226
rect -1764 172170 -1696 172226
rect -1640 172170 -1572 172226
rect -1516 172170 -1448 172226
rect -1392 172170 9234 172226
rect 9290 172170 9358 172226
rect 9414 172170 9482 172226
rect 9538 172170 9606 172226
rect 9662 172170 39954 172226
rect 40010 172170 40078 172226
rect 40134 172170 40202 172226
rect 40258 172170 40326 172226
rect 40382 172170 70674 172226
rect 70730 172170 70798 172226
rect 70854 172170 70922 172226
rect 70978 172170 71046 172226
rect 71102 172170 101394 172226
rect 101450 172170 101518 172226
rect 101574 172170 101642 172226
rect 101698 172170 101766 172226
rect 101822 172170 132114 172226
rect 132170 172170 132238 172226
rect 132294 172170 132362 172226
rect 132418 172170 132486 172226
rect 132542 172170 162834 172226
rect 162890 172170 162958 172226
rect 163014 172170 163082 172226
rect 163138 172170 163206 172226
rect 163262 172170 193554 172226
rect 193610 172170 193678 172226
rect 193734 172170 193802 172226
rect 193858 172170 193926 172226
rect 193982 172170 224274 172226
rect 224330 172170 224398 172226
rect 224454 172170 224522 172226
rect 224578 172170 224646 172226
rect 224702 172170 254994 172226
rect 255050 172170 255118 172226
rect 255174 172170 255242 172226
rect 255298 172170 255366 172226
rect 255422 172170 285714 172226
rect 285770 172170 285838 172226
rect 285894 172170 285962 172226
rect 286018 172170 286086 172226
rect 286142 172170 316434 172226
rect 316490 172170 316558 172226
rect 316614 172170 316682 172226
rect 316738 172170 316806 172226
rect 316862 172170 347154 172226
rect 347210 172170 347278 172226
rect 347334 172170 347402 172226
rect 347458 172170 347526 172226
rect 347582 172170 377874 172226
rect 377930 172170 377998 172226
rect 378054 172170 378122 172226
rect 378178 172170 378246 172226
rect 378302 172170 408594 172226
rect 408650 172170 408718 172226
rect 408774 172170 408842 172226
rect 408898 172170 408966 172226
rect 409022 172170 439314 172226
rect 439370 172170 439438 172226
rect 439494 172170 439562 172226
rect 439618 172170 439686 172226
rect 439742 172170 470034 172226
rect 470090 172170 470158 172226
rect 470214 172170 470282 172226
rect 470338 172170 470406 172226
rect 470462 172170 500754 172226
rect 500810 172170 500878 172226
rect 500934 172170 501002 172226
rect 501058 172170 501126 172226
rect 501182 172170 531474 172226
rect 531530 172170 531598 172226
rect 531654 172170 531722 172226
rect 531778 172170 531846 172226
rect 531902 172170 562194 172226
rect 562250 172170 562318 172226
rect 562374 172170 562442 172226
rect 562498 172170 562566 172226
rect 562622 172170 592914 172226
rect 592970 172170 593038 172226
rect 593094 172170 593162 172226
rect 593218 172170 593286 172226
rect 593342 172170 597456 172226
rect 597512 172170 597580 172226
rect 597636 172170 597704 172226
rect 597760 172170 597828 172226
rect 597884 172170 597980 172226
rect -1916 172102 597980 172170
rect -1916 172046 -1820 172102
rect -1764 172046 -1696 172102
rect -1640 172046 -1572 172102
rect -1516 172046 -1448 172102
rect -1392 172046 9234 172102
rect 9290 172046 9358 172102
rect 9414 172046 9482 172102
rect 9538 172046 9606 172102
rect 9662 172046 39954 172102
rect 40010 172046 40078 172102
rect 40134 172046 40202 172102
rect 40258 172046 40326 172102
rect 40382 172046 70674 172102
rect 70730 172046 70798 172102
rect 70854 172046 70922 172102
rect 70978 172046 71046 172102
rect 71102 172046 101394 172102
rect 101450 172046 101518 172102
rect 101574 172046 101642 172102
rect 101698 172046 101766 172102
rect 101822 172046 132114 172102
rect 132170 172046 132238 172102
rect 132294 172046 132362 172102
rect 132418 172046 132486 172102
rect 132542 172046 162834 172102
rect 162890 172046 162958 172102
rect 163014 172046 163082 172102
rect 163138 172046 163206 172102
rect 163262 172046 193554 172102
rect 193610 172046 193678 172102
rect 193734 172046 193802 172102
rect 193858 172046 193926 172102
rect 193982 172046 224274 172102
rect 224330 172046 224398 172102
rect 224454 172046 224522 172102
rect 224578 172046 224646 172102
rect 224702 172046 254994 172102
rect 255050 172046 255118 172102
rect 255174 172046 255242 172102
rect 255298 172046 255366 172102
rect 255422 172046 285714 172102
rect 285770 172046 285838 172102
rect 285894 172046 285962 172102
rect 286018 172046 286086 172102
rect 286142 172046 316434 172102
rect 316490 172046 316558 172102
rect 316614 172046 316682 172102
rect 316738 172046 316806 172102
rect 316862 172046 347154 172102
rect 347210 172046 347278 172102
rect 347334 172046 347402 172102
rect 347458 172046 347526 172102
rect 347582 172046 377874 172102
rect 377930 172046 377998 172102
rect 378054 172046 378122 172102
rect 378178 172046 378246 172102
rect 378302 172046 408594 172102
rect 408650 172046 408718 172102
rect 408774 172046 408842 172102
rect 408898 172046 408966 172102
rect 409022 172046 439314 172102
rect 439370 172046 439438 172102
rect 439494 172046 439562 172102
rect 439618 172046 439686 172102
rect 439742 172046 470034 172102
rect 470090 172046 470158 172102
rect 470214 172046 470282 172102
rect 470338 172046 470406 172102
rect 470462 172046 500754 172102
rect 500810 172046 500878 172102
rect 500934 172046 501002 172102
rect 501058 172046 501126 172102
rect 501182 172046 531474 172102
rect 531530 172046 531598 172102
rect 531654 172046 531722 172102
rect 531778 172046 531846 172102
rect 531902 172046 562194 172102
rect 562250 172046 562318 172102
rect 562374 172046 562442 172102
rect 562498 172046 562566 172102
rect 562622 172046 592914 172102
rect 592970 172046 593038 172102
rect 593094 172046 593162 172102
rect 593218 172046 593286 172102
rect 593342 172046 597456 172102
rect 597512 172046 597580 172102
rect 597636 172046 597704 172102
rect 597760 172046 597828 172102
rect 597884 172046 597980 172102
rect -1916 171978 597980 172046
rect -1916 171922 -1820 171978
rect -1764 171922 -1696 171978
rect -1640 171922 -1572 171978
rect -1516 171922 -1448 171978
rect -1392 171922 9234 171978
rect 9290 171922 9358 171978
rect 9414 171922 9482 171978
rect 9538 171922 9606 171978
rect 9662 171922 39954 171978
rect 40010 171922 40078 171978
rect 40134 171922 40202 171978
rect 40258 171922 40326 171978
rect 40382 171922 70674 171978
rect 70730 171922 70798 171978
rect 70854 171922 70922 171978
rect 70978 171922 71046 171978
rect 71102 171922 101394 171978
rect 101450 171922 101518 171978
rect 101574 171922 101642 171978
rect 101698 171922 101766 171978
rect 101822 171922 132114 171978
rect 132170 171922 132238 171978
rect 132294 171922 132362 171978
rect 132418 171922 132486 171978
rect 132542 171922 162834 171978
rect 162890 171922 162958 171978
rect 163014 171922 163082 171978
rect 163138 171922 163206 171978
rect 163262 171922 193554 171978
rect 193610 171922 193678 171978
rect 193734 171922 193802 171978
rect 193858 171922 193926 171978
rect 193982 171922 224274 171978
rect 224330 171922 224398 171978
rect 224454 171922 224522 171978
rect 224578 171922 224646 171978
rect 224702 171922 254994 171978
rect 255050 171922 255118 171978
rect 255174 171922 255242 171978
rect 255298 171922 255366 171978
rect 255422 171922 285714 171978
rect 285770 171922 285838 171978
rect 285894 171922 285962 171978
rect 286018 171922 286086 171978
rect 286142 171922 316434 171978
rect 316490 171922 316558 171978
rect 316614 171922 316682 171978
rect 316738 171922 316806 171978
rect 316862 171922 347154 171978
rect 347210 171922 347278 171978
rect 347334 171922 347402 171978
rect 347458 171922 347526 171978
rect 347582 171922 377874 171978
rect 377930 171922 377998 171978
rect 378054 171922 378122 171978
rect 378178 171922 378246 171978
rect 378302 171922 408594 171978
rect 408650 171922 408718 171978
rect 408774 171922 408842 171978
rect 408898 171922 408966 171978
rect 409022 171922 439314 171978
rect 439370 171922 439438 171978
rect 439494 171922 439562 171978
rect 439618 171922 439686 171978
rect 439742 171922 470034 171978
rect 470090 171922 470158 171978
rect 470214 171922 470282 171978
rect 470338 171922 470406 171978
rect 470462 171922 500754 171978
rect 500810 171922 500878 171978
rect 500934 171922 501002 171978
rect 501058 171922 501126 171978
rect 501182 171922 531474 171978
rect 531530 171922 531598 171978
rect 531654 171922 531722 171978
rect 531778 171922 531846 171978
rect 531902 171922 562194 171978
rect 562250 171922 562318 171978
rect 562374 171922 562442 171978
rect 562498 171922 562566 171978
rect 562622 171922 592914 171978
rect 592970 171922 593038 171978
rect 593094 171922 593162 171978
rect 593218 171922 593286 171978
rect 593342 171922 597456 171978
rect 597512 171922 597580 171978
rect 597636 171922 597704 171978
rect 597760 171922 597828 171978
rect 597884 171922 597980 171978
rect -1916 171826 597980 171922
rect -1916 166350 597980 166446
rect -1916 166294 -860 166350
rect -804 166294 -736 166350
rect -680 166294 -612 166350
rect -556 166294 -488 166350
rect -432 166294 5514 166350
rect 5570 166294 5638 166350
rect 5694 166294 5762 166350
rect 5818 166294 5886 166350
rect 5942 166294 36234 166350
rect 36290 166294 36358 166350
rect 36414 166294 36482 166350
rect 36538 166294 36606 166350
rect 36662 166294 66954 166350
rect 67010 166294 67078 166350
rect 67134 166294 67202 166350
rect 67258 166294 67326 166350
rect 67382 166294 97674 166350
rect 97730 166294 97798 166350
rect 97854 166294 97922 166350
rect 97978 166294 98046 166350
rect 98102 166294 128394 166350
rect 128450 166294 128518 166350
rect 128574 166294 128642 166350
rect 128698 166294 128766 166350
rect 128822 166294 159114 166350
rect 159170 166294 159238 166350
rect 159294 166294 159362 166350
rect 159418 166294 159486 166350
rect 159542 166294 189834 166350
rect 189890 166294 189958 166350
rect 190014 166294 190082 166350
rect 190138 166294 190206 166350
rect 190262 166294 220554 166350
rect 220610 166294 220678 166350
rect 220734 166294 220802 166350
rect 220858 166294 220926 166350
rect 220982 166294 251274 166350
rect 251330 166294 251398 166350
rect 251454 166294 251522 166350
rect 251578 166294 251646 166350
rect 251702 166294 281994 166350
rect 282050 166294 282118 166350
rect 282174 166294 282242 166350
rect 282298 166294 282366 166350
rect 282422 166294 312714 166350
rect 312770 166294 312838 166350
rect 312894 166294 312962 166350
rect 313018 166294 313086 166350
rect 313142 166294 343434 166350
rect 343490 166294 343558 166350
rect 343614 166294 343682 166350
rect 343738 166294 343806 166350
rect 343862 166294 374154 166350
rect 374210 166294 374278 166350
rect 374334 166294 374402 166350
rect 374458 166294 374526 166350
rect 374582 166294 404874 166350
rect 404930 166294 404998 166350
rect 405054 166294 405122 166350
rect 405178 166294 405246 166350
rect 405302 166294 435594 166350
rect 435650 166294 435718 166350
rect 435774 166294 435842 166350
rect 435898 166294 435966 166350
rect 436022 166294 466314 166350
rect 466370 166294 466438 166350
rect 466494 166294 466562 166350
rect 466618 166294 466686 166350
rect 466742 166294 497034 166350
rect 497090 166294 497158 166350
rect 497214 166294 497282 166350
rect 497338 166294 497406 166350
rect 497462 166294 527754 166350
rect 527810 166294 527878 166350
rect 527934 166294 528002 166350
rect 528058 166294 528126 166350
rect 528182 166294 558474 166350
rect 558530 166294 558598 166350
rect 558654 166294 558722 166350
rect 558778 166294 558846 166350
rect 558902 166294 589194 166350
rect 589250 166294 589318 166350
rect 589374 166294 589442 166350
rect 589498 166294 589566 166350
rect 589622 166294 596496 166350
rect 596552 166294 596620 166350
rect 596676 166294 596744 166350
rect 596800 166294 596868 166350
rect 596924 166294 597980 166350
rect -1916 166226 597980 166294
rect -1916 166170 -860 166226
rect -804 166170 -736 166226
rect -680 166170 -612 166226
rect -556 166170 -488 166226
rect -432 166170 5514 166226
rect 5570 166170 5638 166226
rect 5694 166170 5762 166226
rect 5818 166170 5886 166226
rect 5942 166170 36234 166226
rect 36290 166170 36358 166226
rect 36414 166170 36482 166226
rect 36538 166170 36606 166226
rect 36662 166170 66954 166226
rect 67010 166170 67078 166226
rect 67134 166170 67202 166226
rect 67258 166170 67326 166226
rect 67382 166170 97674 166226
rect 97730 166170 97798 166226
rect 97854 166170 97922 166226
rect 97978 166170 98046 166226
rect 98102 166170 128394 166226
rect 128450 166170 128518 166226
rect 128574 166170 128642 166226
rect 128698 166170 128766 166226
rect 128822 166170 159114 166226
rect 159170 166170 159238 166226
rect 159294 166170 159362 166226
rect 159418 166170 159486 166226
rect 159542 166170 189834 166226
rect 189890 166170 189958 166226
rect 190014 166170 190082 166226
rect 190138 166170 190206 166226
rect 190262 166170 220554 166226
rect 220610 166170 220678 166226
rect 220734 166170 220802 166226
rect 220858 166170 220926 166226
rect 220982 166170 251274 166226
rect 251330 166170 251398 166226
rect 251454 166170 251522 166226
rect 251578 166170 251646 166226
rect 251702 166170 281994 166226
rect 282050 166170 282118 166226
rect 282174 166170 282242 166226
rect 282298 166170 282366 166226
rect 282422 166170 312714 166226
rect 312770 166170 312838 166226
rect 312894 166170 312962 166226
rect 313018 166170 313086 166226
rect 313142 166170 343434 166226
rect 343490 166170 343558 166226
rect 343614 166170 343682 166226
rect 343738 166170 343806 166226
rect 343862 166170 374154 166226
rect 374210 166170 374278 166226
rect 374334 166170 374402 166226
rect 374458 166170 374526 166226
rect 374582 166170 404874 166226
rect 404930 166170 404998 166226
rect 405054 166170 405122 166226
rect 405178 166170 405246 166226
rect 405302 166170 435594 166226
rect 435650 166170 435718 166226
rect 435774 166170 435842 166226
rect 435898 166170 435966 166226
rect 436022 166170 466314 166226
rect 466370 166170 466438 166226
rect 466494 166170 466562 166226
rect 466618 166170 466686 166226
rect 466742 166170 497034 166226
rect 497090 166170 497158 166226
rect 497214 166170 497282 166226
rect 497338 166170 497406 166226
rect 497462 166170 527754 166226
rect 527810 166170 527878 166226
rect 527934 166170 528002 166226
rect 528058 166170 528126 166226
rect 528182 166170 558474 166226
rect 558530 166170 558598 166226
rect 558654 166170 558722 166226
rect 558778 166170 558846 166226
rect 558902 166170 589194 166226
rect 589250 166170 589318 166226
rect 589374 166170 589442 166226
rect 589498 166170 589566 166226
rect 589622 166170 596496 166226
rect 596552 166170 596620 166226
rect 596676 166170 596744 166226
rect 596800 166170 596868 166226
rect 596924 166170 597980 166226
rect -1916 166102 597980 166170
rect -1916 166046 -860 166102
rect -804 166046 -736 166102
rect -680 166046 -612 166102
rect -556 166046 -488 166102
rect -432 166046 5514 166102
rect 5570 166046 5638 166102
rect 5694 166046 5762 166102
rect 5818 166046 5886 166102
rect 5942 166046 36234 166102
rect 36290 166046 36358 166102
rect 36414 166046 36482 166102
rect 36538 166046 36606 166102
rect 36662 166046 66954 166102
rect 67010 166046 67078 166102
rect 67134 166046 67202 166102
rect 67258 166046 67326 166102
rect 67382 166046 97674 166102
rect 97730 166046 97798 166102
rect 97854 166046 97922 166102
rect 97978 166046 98046 166102
rect 98102 166046 128394 166102
rect 128450 166046 128518 166102
rect 128574 166046 128642 166102
rect 128698 166046 128766 166102
rect 128822 166046 159114 166102
rect 159170 166046 159238 166102
rect 159294 166046 159362 166102
rect 159418 166046 159486 166102
rect 159542 166046 189834 166102
rect 189890 166046 189958 166102
rect 190014 166046 190082 166102
rect 190138 166046 190206 166102
rect 190262 166046 220554 166102
rect 220610 166046 220678 166102
rect 220734 166046 220802 166102
rect 220858 166046 220926 166102
rect 220982 166046 251274 166102
rect 251330 166046 251398 166102
rect 251454 166046 251522 166102
rect 251578 166046 251646 166102
rect 251702 166046 281994 166102
rect 282050 166046 282118 166102
rect 282174 166046 282242 166102
rect 282298 166046 282366 166102
rect 282422 166046 312714 166102
rect 312770 166046 312838 166102
rect 312894 166046 312962 166102
rect 313018 166046 313086 166102
rect 313142 166046 343434 166102
rect 343490 166046 343558 166102
rect 343614 166046 343682 166102
rect 343738 166046 343806 166102
rect 343862 166046 374154 166102
rect 374210 166046 374278 166102
rect 374334 166046 374402 166102
rect 374458 166046 374526 166102
rect 374582 166046 404874 166102
rect 404930 166046 404998 166102
rect 405054 166046 405122 166102
rect 405178 166046 405246 166102
rect 405302 166046 435594 166102
rect 435650 166046 435718 166102
rect 435774 166046 435842 166102
rect 435898 166046 435966 166102
rect 436022 166046 466314 166102
rect 466370 166046 466438 166102
rect 466494 166046 466562 166102
rect 466618 166046 466686 166102
rect 466742 166046 497034 166102
rect 497090 166046 497158 166102
rect 497214 166046 497282 166102
rect 497338 166046 497406 166102
rect 497462 166046 527754 166102
rect 527810 166046 527878 166102
rect 527934 166046 528002 166102
rect 528058 166046 528126 166102
rect 528182 166046 558474 166102
rect 558530 166046 558598 166102
rect 558654 166046 558722 166102
rect 558778 166046 558846 166102
rect 558902 166046 589194 166102
rect 589250 166046 589318 166102
rect 589374 166046 589442 166102
rect 589498 166046 589566 166102
rect 589622 166046 596496 166102
rect 596552 166046 596620 166102
rect 596676 166046 596744 166102
rect 596800 166046 596868 166102
rect 596924 166046 597980 166102
rect -1916 165978 597980 166046
rect -1916 165922 -860 165978
rect -804 165922 -736 165978
rect -680 165922 -612 165978
rect -556 165922 -488 165978
rect -432 165922 5514 165978
rect 5570 165922 5638 165978
rect 5694 165922 5762 165978
rect 5818 165922 5886 165978
rect 5942 165922 36234 165978
rect 36290 165922 36358 165978
rect 36414 165922 36482 165978
rect 36538 165922 36606 165978
rect 36662 165922 66954 165978
rect 67010 165922 67078 165978
rect 67134 165922 67202 165978
rect 67258 165922 67326 165978
rect 67382 165922 97674 165978
rect 97730 165922 97798 165978
rect 97854 165922 97922 165978
rect 97978 165922 98046 165978
rect 98102 165922 128394 165978
rect 128450 165922 128518 165978
rect 128574 165922 128642 165978
rect 128698 165922 128766 165978
rect 128822 165922 159114 165978
rect 159170 165922 159238 165978
rect 159294 165922 159362 165978
rect 159418 165922 159486 165978
rect 159542 165922 189834 165978
rect 189890 165922 189958 165978
rect 190014 165922 190082 165978
rect 190138 165922 190206 165978
rect 190262 165922 220554 165978
rect 220610 165922 220678 165978
rect 220734 165922 220802 165978
rect 220858 165922 220926 165978
rect 220982 165922 251274 165978
rect 251330 165922 251398 165978
rect 251454 165922 251522 165978
rect 251578 165922 251646 165978
rect 251702 165922 281994 165978
rect 282050 165922 282118 165978
rect 282174 165922 282242 165978
rect 282298 165922 282366 165978
rect 282422 165922 312714 165978
rect 312770 165922 312838 165978
rect 312894 165922 312962 165978
rect 313018 165922 313086 165978
rect 313142 165922 343434 165978
rect 343490 165922 343558 165978
rect 343614 165922 343682 165978
rect 343738 165922 343806 165978
rect 343862 165922 374154 165978
rect 374210 165922 374278 165978
rect 374334 165922 374402 165978
rect 374458 165922 374526 165978
rect 374582 165922 404874 165978
rect 404930 165922 404998 165978
rect 405054 165922 405122 165978
rect 405178 165922 405246 165978
rect 405302 165922 435594 165978
rect 435650 165922 435718 165978
rect 435774 165922 435842 165978
rect 435898 165922 435966 165978
rect 436022 165922 466314 165978
rect 466370 165922 466438 165978
rect 466494 165922 466562 165978
rect 466618 165922 466686 165978
rect 466742 165922 497034 165978
rect 497090 165922 497158 165978
rect 497214 165922 497282 165978
rect 497338 165922 497406 165978
rect 497462 165922 527754 165978
rect 527810 165922 527878 165978
rect 527934 165922 528002 165978
rect 528058 165922 528126 165978
rect 528182 165922 558474 165978
rect 558530 165922 558598 165978
rect 558654 165922 558722 165978
rect 558778 165922 558846 165978
rect 558902 165922 589194 165978
rect 589250 165922 589318 165978
rect 589374 165922 589442 165978
rect 589498 165922 589566 165978
rect 589622 165922 596496 165978
rect 596552 165922 596620 165978
rect 596676 165922 596744 165978
rect 596800 165922 596868 165978
rect 596924 165922 597980 165978
rect -1916 165826 597980 165922
rect -1916 154350 597980 154446
rect -1916 154294 -1820 154350
rect -1764 154294 -1696 154350
rect -1640 154294 -1572 154350
rect -1516 154294 -1448 154350
rect -1392 154294 9234 154350
rect 9290 154294 9358 154350
rect 9414 154294 9482 154350
rect 9538 154294 9606 154350
rect 9662 154294 39954 154350
rect 40010 154294 40078 154350
rect 40134 154294 40202 154350
rect 40258 154294 40326 154350
rect 40382 154294 70674 154350
rect 70730 154294 70798 154350
rect 70854 154294 70922 154350
rect 70978 154294 71046 154350
rect 71102 154294 101394 154350
rect 101450 154294 101518 154350
rect 101574 154294 101642 154350
rect 101698 154294 101766 154350
rect 101822 154294 132114 154350
rect 132170 154294 132238 154350
rect 132294 154294 132362 154350
rect 132418 154294 132486 154350
rect 132542 154294 162834 154350
rect 162890 154294 162958 154350
rect 163014 154294 163082 154350
rect 163138 154294 163206 154350
rect 163262 154294 193554 154350
rect 193610 154294 193678 154350
rect 193734 154294 193802 154350
rect 193858 154294 193926 154350
rect 193982 154294 224274 154350
rect 224330 154294 224398 154350
rect 224454 154294 224522 154350
rect 224578 154294 224646 154350
rect 224702 154294 254994 154350
rect 255050 154294 255118 154350
rect 255174 154294 255242 154350
rect 255298 154294 255366 154350
rect 255422 154294 285714 154350
rect 285770 154294 285838 154350
rect 285894 154294 285962 154350
rect 286018 154294 286086 154350
rect 286142 154294 316434 154350
rect 316490 154294 316558 154350
rect 316614 154294 316682 154350
rect 316738 154294 316806 154350
rect 316862 154294 347154 154350
rect 347210 154294 347278 154350
rect 347334 154294 347402 154350
rect 347458 154294 347526 154350
rect 347582 154294 377874 154350
rect 377930 154294 377998 154350
rect 378054 154294 378122 154350
rect 378178 154294 378246 154350
rect 378302 154294 408594 154350
rect 408650 154294 408718 154350
rect 408774 154294 408842 154350
rect 408898 154294 408966 154350
rect 409022 154294 439314 154350
rect 439370 154294 439438 154350
rect 439494 154294 439562 154350
rect 439618 154294 439686 154350
rect 439742 154294 470034 154350
rect 470090 154294 470158 154350
rect 470214 154294 470282 154350
rect 470338 154294 470406 154350
rect 470462 154294 500754 154350
rect 500810 154294 500878 154350
rect 500934 154294 501002 154350
rect 501058 154294 501126 154350
rect 501182 154294 531474 154350
rect 531530 154294 531598 154350
rect 531654 154294 531722 154350
rect 531778 154294 531846 154350
rect 531902 154294 562194 154350
rect 562250 154294 562318 154350
rect 562374 154294 562442 154350
rect 562498 154294 562566 154350
rect 562622 154294 592914 154350
rect 592970 154294 593038 154350
rect 593094 154294 593162 154350
rect 593218 154294 593286 154350
rect 593342 154294 597456 154350
rect 597512 154294 597580 154350
rect 597636 154294 597704 154350
rect 597760 154294 597828 154350
rect 597884 154294 597980 154350
rect -1916 154226 597980 154294
rect -1916 154170 -1820 154226
rect -1764 154170 -1696 154226
rect -1640 154170 -1572 154226
rect -1516 154170 -1448 154226
rect -1392 154170 9234 154226
rect 9290 154170 9358 154226
rect 9414 154170 9482 154226
rect 9538 154170 9606 154226
rect 9662 154170 39954 154226
rect 40010 154170 40078 154226
rect 40134 154170 40202 154226
rect 40258 154170 40326 154226
rect 40382 154170 70674 154226
rect 70730 154170 70798 154226
rect 70854 154170 70922 154226
rect 70978 154170 71046 154226
rect 71102 154170 101394 154226
rect 101450 154170 101518 154226
rect 101574 154170 101642 154226
rect 101698 154170 101766 154226
rect 101822 154170 132114 154226
rect 132170 154170 132238 154226
rect 132294 154170 132362 154226
rect 132418 154170 132486 154226
rect 132542 154170 162834 154226
rect 162890 154170 162958 154226
rect 163014 154170 163082 154226
rect 163138 154170 163206 154226
rect 163262 154170 193554 154226
rect 193610 154170 193678 154226
rect 193734 154170 193802 154226
rect 193858 154170 193926 154226
rect 193982 154170 224274 154226
rect 224330 154170 224398 154226
rect 224454 154170 224522 154226
rect 224578 154170 224646 154226
rect 224702 154170 254994 154226
rect 255050 154170 255118 154226
rect 255174 154170 255242 154226
rect 255298 154170 255366 154226
rect 255422 154170 285714 154226
rect 285770 154170 285838 154226
rect 285894 154170 285962 154226
rect 286018 154170 286086 154226
rect 286142 154170 316434 154226
rect 316490 154170 316558 154226
rect 316614 154170 316682 154226
rect 316738 154170 316806 154226
rect 316862 154170 347154 154226
rect 347210 154170 347278 154226
rect 347334 154170 347402 154226
rect 347458 154170 347526 154226
rect 347582 154170 377874 154226
rect 377930 154170 377998 154226
rect 378054 154170 378122 154226
rect 378178 154170 378246 154226
rect 378302 154170 408594 154226
rect 408650 154170 408718 154226
rect 408774 154170 408842 154226
rect 408898 154170 408966 154226
rect 409022 154170 439314 154226
rect 439370 154170 439438 154226
rect 439494 154170 439562 154226
rect 439618 154170 439686 154226
rect 439742 154170 470034 154226
rect 470090 154170 470158 154226
rect 470214 154170 470282 154226
rect 470338 154170 470406 154226
rect 470462 154170 500754 154226
rect 500810 154170 500878 154226
rect 500934 154170 501002 154226
rect 501058 154170 501126 154226
rect 501182 154170 531474 154226
rect 531530 154170 531598 154226
rect 531654 154170 531722 154226
rect 531778 154170 531846 154226
rect 531902 154170 562194 154226
rect 562250 154170 562318 154226
rect 562374 154170 562442 154226
rect 562498 154170 562566 154226
rect 562622 154170 592914 154226
rect 592970 154170 593038 154226
rect 593094 154170 593162 154226
rect 593218 154170 593286 154226
rect 593342 154170 597456 154226
rect 597512 154170 597580 154226
rect 597636 154170 597704 154226
rect 597760 154170 597828 154226
rect 597884 154170 597980 154226
rect -1916 154102 597980 154170
rect -1916 154046 -1820 154102
rect -1764 154046 -1696 154102
rect -1640 154046 -1572 154102
rect -1516 154046 -1448 154102
rect -1392 154046 9234 154102
rect 9290 154046 9358 154102
rect 9414 154046 9482 154102
rect 9538 154046 9606 154102
rect 9662 154046 39954 154102
rect 40010 154046 40078 154102
rect 40134 154046 40202 154102
rect 40258 154046 40326 154102
rect 40382 154046 70674 154102
rect 70730 154046 70798 154102
rect 70854 154046 70922 154102
rect 70978 154046 71046 154102
rect 71102 154046 101394 154102
rect 101450 154046 101518 154102
rect 101574 154046 101642 154102
rect 101698 154046 101766 154102
rect 101822 154046 132114 154102
rect 132170 154046 132238 154102
rect 132294 154046 132362 154102
rect 132418 154046 132486 154102
rect 132542 154046 162834 154102
rect 162890 154046 162958 154102
rect 163014 154046 163082 154102
rect 163138 154046 163206 154102
rect 163262 154046 193554 154102
rect 193610 154046 193678 154102
rect 193734 154046 193802 154102
rect 193858 154046 193926 154102
rect 193982 154046 224274 154102
rect 224330 154046 224398 154102
rect 224454 154046 224522 154102
rect 224578 154046 224646 154102
rect 224702 154046 254994 154102
rect 255050 154046 255118 154102
rect 255174 154046 255242 154102
rect 255298 154046 255366 154102
rect 255422 154046 285714 154102
rect 285770 154046 285838 154102
rect 285894 154046 285962 154102
rect 286018 154046 286086 154102
rect 286142 154046 316434 154102
rect 316490 154046 316558 154102
rect 316614 154046 316682 154102
rect 316738 154046 316806 154102
rect 316862 154046 347154 154102
rect 347210 154046 347278 154102
rect 347334 154046 347402 154102
rect 347458 154046 347526 154102
rect 347582 154046 377874 154102
rect 377930 154046 377998 154102
rect 378054 154046 378122 154102
rect 378178 154046 378246 154102
rect 378302 154046 408594 154102
rect 408650 154046 408718 154102
rect 408774 154046 408842 154102
rect 408898 154046 408966 154102
rect 409022 154046 439314 154102
rect 439370 154046 439438 154102
rect 439494 154046 439562 154102
rect 439618 154046 439686 154102
rect 439742 154046 470034 154102
rect 470090 154046 470158 154102
rect 470214 154046 470282 154102
rect 470338 154046 470406 154102
rect 470462 154046 500754 154102
rect 500810 154046 500878 154102
rect 500934 154046 501002 154102
rect 501058 154046 501126 154102
rect 501182 154046 531474 154102
rect 531530 154046 531598 154102
rect 531654 154046 531722 154102
rect 531778 154046 531846 154102
rect 531902 154046 562194 154102
rect 562250 154046 562318 154102
rect 562374 154046 562442 154102
rect 562498 154046 562566 154102
rect 562622 154046 592914 154102
rect 592970 154046 593038 154102
rect 593094 154046 593162 154102
rect 593218 154046 593286 154102
rect 593342 154046 597456 154102
rect 597512 154046 597580 154102
rect 597636 154046 597704 154102
rect 597760 154046 597828 154102
rect 597884 154046 597980 154102
rect -1916 153978 597980 154046
rect -1916 153922 -1820 153978
rect -1764 153922 -1696 153978
rect -1640 153922 -1572 153978
rect -1516 153922 -1448 153978
rect -1392 153922 9234 153978
rect 9290 153922 9358 153978
rect 9414 153922 9482 153978
rect 9538 153922 9606 153978
rect 9662 153922 39954 153978
rect 40010 153922 40078 153978
rect 40134 153922 40202 153978
rect 40258 153922 40326 153978
rect 40382 153922 70674 153978
rect 70730 153922 70798 153978
rect 70854 153922 70922 153978
rect 70978 153922 71046 153978
rect 71102 153922 101394 153978
rect 101450 153922 101518 153978
rect 101574 153922 101642 153978
rect 101698 153922 101766 153978
rect 101822 153922 132114 153978
rect 132170 153922 132238 153978
rect 132294 153922 132362 153978
rect 132418 153922 132486 153978
rect 132542 153922 162834 153978
rect 162890 153922 162958 153978
rect 163014 153922 163082 153978
rect 163138 153922 163206 153978
rect 163262 153922 193554 153978
rect 193610 153922 193678 153978
rect 193734 153922 193802 153978
rect 193858 153922 193926 153978
rect 193982 153922 224274 153978
rect 224330 153922 224398 153978
rect 224454 153922 224522 153978
rect 224578 153922 224646 153978
rect 224702 153922 254994 153978
rect 255050 153922 255118 153978
rect 255174 153922 255242 153978
rect 255298 153922 255366 153978
rect 255422 153922 285714 153978
rect 285770 153922 285838 153978
rect 285894 153922 285962 153978
rect 286018 153922 286086 153978
rect 286142 153922 316434 153978
rect 316490 153922 316558 153978
rect 316614 153922 316682 153978
rect 316738 153922 316806 153978
rect 316862 153922 347154 153978
rect 347210 153922 347278 153978
rect 347334 153922 347402 153978
rect 347458 153922 347526 153978
rect 347582 153922 377874 153978
rect 377930 153922 377998 153978
rect 378054 153922 378122 153978
rect 378178 153922 378246 153978
rect 378302 153922 408594 153978
rect 408650 153922 408718 153978
rect 408774 153922 408842 153978
rect 408898 153922 408966 153978
rect 409022 153922 439314 153978
rect 439370 153922 439438 153978
rect 439494 153922 439562 153978
rect 439618 153922 439686 153978
rect 439742 153922 470034 153978
rect 470090 153922 470158 153978
rect 470214 153922 470282 153978
rect 470338 153922 470406 153978
rect 470462 153922 500754 153978
rect 500810 153922 500878 153978
rect 500934 153922 501002 153978
rect 501058 153922 501126 153978
rect 501182 153922 531474 153978
rect 531530 153922 531598 153978
rect 531654 153922 531722 153978
rect 531778 153922 531846 153978
rect 531902 153922 562194 153978
rect 562250 153922 562318 153978
rect 562374 153922 562442 153978
rect 562498 153922 562566 153978
rect 562622 153922 592914 153978
rect 592970 153922 593038 153978
rect 593094 153922 593162 153978
rect 593218 153922 593286 153978
rect 593342 153922 597456 153978
rect 597512 153922 597580 153978
rect 597636 153922 597704 153978
rect 597760 153922 597828 153978
rect 597884 153922 597980 153978
rect -1916 153826 597980 153922
rect -1916 148350 597980 148446
rect -1916 148294 -860 148350
rect -804 148294 -736 148350
rect -680 148294 -612 148350
rect -556 148294 -488 148350
rect -432 148294 5514 148350
rect 5570 148294 5638 148350
rect 5694 148294 5762 148350
rect 5818 148294 5886 148350
rect 5942 148294 36234 148350
rect 36290 148294 36358 148350
rect 36414 148294 36482 148350
rect 36538 148294 36606 148350
rect 36662 148294 66954 148350
rect 67010 148294 67078 148350
rect 67134 148294 67202 148350
rect 67258 148294 67326 148350
rect 67382 148294 97674 148350
rect 97730 148294 97798 148350
rect 97854 148294 97922 148350
rect 97978 148294 98046 148350
rect 98102 148294 128394 148350
rect 128450 148294 128518 148350
rect 128574 148294 128642 148350
rect 128698 148294 128766 148350
rect 128822 148294 159114 148350
rect 159170 148294 159238 148350
rect 159294 148294 159362 148350
rect 159418 148294 159486 148350
rect 159542 148294 189834 148350
rect 189890 148294 189958 148350
rect 190014 148294 190082 148350
rect 190138 148294 190206 148350
rect 190262 148294 220554 148350
rect 220610 148294 220678 148350
rect 220734 148294 220802 148350
rect 220858 148294 220926 148350
rect 220982 148294 251274 148350
rect 251330 148294 251398 148350
rect 251454 148294 251522 148350
rect 251578 148294 251646 148350
rect 251702 148294 281994 148350
rect 282050 148294 282118 148350
rect 282174 148294 282242 148350
rect 282298 148294 282366 148350
rect 282422 148294 312714 148350
rect 312770 148294 312838 148350
rect 312894 148294 312962 148350
rect 313018 148294 313086 148350
rect 313142 148294 343434 148350
rect 343490 148294 343558 148350
rect 343614 148294 343682 148350
rect 343738 148294 343806 148350
rect 343862 148294 374154 148350
rect 374210 148294 374278 148350
rect 374334 148294 374402 148350
rect 374458 148294 374526 148350
rect 374582 148294 404874 148350
rect 404930 148294 404998 148350
rect 405054 148294 405122 148350
rect 405178 148294 405246 148350
rect 405302 148294 435594 148350
rect 435650 148294 435718 148350
rect 435774 148294 435842 148350
rect 435898 148294 435966 148350
rect 436022 148294 466314 148350
rect 466370 148294 466438 148350
rect 466494 148294 466562 148350
rect 466618 148294 466686 148350
rect 466742 148294 497034 148350
rect 497090 148294 497158 148350
rect 497214 148294 497282 148350
rect 497338 148294 497406 148350
rect 497462 148294 527754 148350
rect 527810 148294 527878 148350
rect 527934 148294 528002 148350
rect 528058 148294 528126 148350
rect 528182 148294 558474 148350
rect 558530 148294 558598 148350
rect 558654 148294 558722 148350
rect 558778 148294 558846 148350
rect 558902 148294 589194 148350
rect 589250 148294 589318 148350
rect 589374 148294 589442 148350
rect 589498 148294 589566 148350
rect 589622 148294 596496 148350
rect 596552 148294 596620 148350
rect 596676 148294 596744 148350
rect 596800 148294 596868 148350
rect 596924 148294 597980 148350
rect -1916 148226 597980 148294
rect -1916 148170 -860 148226
rect -804 148170 -736 148226
rect -680 148170 -612 148226
rect -556 148170 -488 148226
rect -432 148170 5514 148226
rect 5570 148170 5638 148226
rect 5694 148170 5762 148226
rect 5818 148170 5886 148226
rect 5942 148170 36234 148226
rect 36290 148170 36358 148226
rect 36414 148170 36482 148226
rect 36538 148170 36606 148226
rect 36662 148170 66954 148226
rect 67010 148170 67078 148226
rect 67134 148170 67202 148226
rect 67258 148170 67326 148226
rect 67382 148170 97674 148226
rect 97730 148170 97798 148226
rect 97854 148170 97922 148226
rect 97978 148170 98046 148226
rect 98102 148170 128394 148226
rect 128450 148170 128518 148226
rect 128574 148170 128642 148226
rect 128698 148170 128766 148226
rect 128822 148170 159114 148226
rect 159170 148170 159238 148226
rect 159294 148170 159362 148226
rect 159418 148170 159486 148226
rect 159542 148170 189834 148226
rect 189890 148170 189958 148226
rect 190014 148170 190082 148226
rect 190138 148170 190206 148226
rect 190262 148170 220554 148226
rect 220610 148170 220678 148226
rect 220734 148170 220802 148226
rect 220858 148170 220926 148226
rect 220982 148170 251274 148226
rect 251330 148170 251398 148226
rect 251454 148170 251522 148226
rect 251578 148170 251646 148226
rect 251702 148170 281994 148226
rect 282050 148170 282118 148226
rect 282174 148170 282242 148226
rect 282298 148170 282366 148226
rect 282422 148170 312714 148226
rect 312770 148170 312838 148226
rect 312894 148170 312962 148226
rect 313018 148170 313086 148226
rect 313142 148170 343434 148226
rect 343490 148170 343558 148226
rect 343614 148170 343682 148226
rect 343738 148170 343806 148226
rect 343862 148170 374154 148226
rect 374210 148170 374278 148226
rect 374334 148170 374402 148226
rect 374458 148170 374526 148226
rect 374582 148170 404874 148226
rect 404930 148170 404998 148226
rect 405054 148170 405122 148226
rect 405178 148170 405246 148226
rect 405302 148170 435594 148226
rect 435650 148170 435718 148226
rect 435774 148170 435842 148226
rect 435898 148170 435966 148226
rect 436022 148170 466314 148226
rect 466370 148170 466438 148226
rect 466494 148170 466562 148226
rect 466618 148170 466686 148226
rect 466742 148170 497034 148226
rect 497090 148170 497158 148226
rect 497214 148170 497282 148226
rect 497338 148170 497406 148226
rect 497462 148170 527754 148226
rect 527810 148170 527878 148226
rect 527934 148170 528002 148226
rect 528058 148170 528126 148226
rect 528182 148170 558474 148226
rect 558530 148170 558598 148226
rect 558654 148170 558722 148226
rect 558778 148170 558846 148226
rect 558902 148170 589194 148226
rect 589250 148170 589318 148226
rect 589374 148170 589442 148226
rect 589498 148170 589566 148226
rect 589622 148170 596496 148226
rect 596552 148170 596620 148226
rect 596676 148170 596744 148226
rect 596800 148170 596868 148226
rect 596924 148170 597980 148226
rect -1916 148102 597980 148170
rect -1916 148046 -860 148102
rect -804 148046 -736 148102
rect -680 148046 -612 148102
rect -556 148046 -488 148102
rect -432 148046 5514 148102
rect 5570 148046 5638 148102
rect 5694 148046 5762 148102
rect 5818 148046 5886 148102
rect 5942 148046 36234 148102
rect 36290 148046 36358 148102
rect 36414 148046 36482 148102
rect 36538 148046 36606 148102
rect 36662 148046 66954 148102
rect 67010 148046 67078 148102
rect 67134 148046 67202 148102
rect 67258 148046 67326 148102
rect 67382 148046 97674 148102
rect 97730 148046 97798 148102
rect 97854 148046 97922 148102
rect 97978 148046 98046 148102
rect 98102 148046 128394 148102
rect 128450 148046 128518 148102
rect 128574 148046 128642 148102
rect 128698 148046 128766 148102
rect 128822 148046 159114 148102
rect 159170 148046 159238 148102
rect 159294 148046 159362 148102
rect 159418 148046 159486 148102
rect 159542 148046 189834 148102
rect 189890 148046 189958 148102
rect 190014 148046 190082 148102
rect 190138 148046 190206 148102
rect 190262 148046 220554 148102
rect 220610 148046 220678 148102
rect 220734 148046 220802 148102
rect 220858 148046 220926 148102
rect 220982 148046 251274 148102
rect 251330 148046 251398 148102
rect 251454 148046 251522 148102
rect 251578 148046 251646 148102
rect 251702 148046 281994 148102
rect 282050 148046 282118 148102
rect 282174 148046 282242 148102
rect 282298 148046 282366 148102
rect 282422 148046 312714 148102
rect 312770 148046 312838 148102
rect 312894 148046 312962 148102
rect 313018 148046 313086 148102
rect 313142 148046 343434 148102
rect 343490 148046 343558 148102
rect 343614 148046 343682 148102
rect 343738 148046 343806 148102
rect 343862 148046 374154 148102
rect 374210 148046 374278 148102
rect 374334 148046 374402 148102
rect 374458 148046 374526 148102
rect 374582 148046 404874 148102
rect 404930 148046 404998 148102
rect 405054 148046 405122 148102
rect 405178 148046 405246 148102
rect 405302 148046 435594 148102
rect 435650 148046 435718 148102
rect 435774 148046 435842 148102
rect 435898 148046 435966 148102
rect 436022 148046 466314 148102
rect 466370 148046 466438 148102
rect 466494 148046 466562 148102
rect 466618 148046 466686 148102
rect 466742 148046 497034 148102
rect 497090 148046 497158 148102
rect 497214 148046 497282 148102
rect 497338 148046 497406 148102
rect 497462 148046 527754 148102
rect 527810 148046 527878 148102
rect 527934 148046 528002 148102
rect 528058 148046 528126 148102
rect 528182 148046 558474 148102
rect 558530 148046 558598 148102
rect 558654 148046 558722 148102
rect 558778 148046 558846 148102
rect 558902 148046 589194 148102
rect 589250 148046 589318 148102
rect 589374 148046 589442 148102
rect 589498 148046 589566 148102
rect 589622 148046 596496 148102
rect 596552 148046 596620 148102
rect 596676 148046 596744 148102
rect 596800 148046 596868 148102
rect 596924 148046 597980 148102
rect -1916 147978 597980 148046
rect -1916 147922 -860 147978
rect -804 147922 -736 147978
rect -680 147922 -612 147978
rect -556 147922 -488 147978
rect -432 147922 5514 147978
rect 5570 147922 5638 147978
rect 5694 147922 5762 147978
rect 5818 147922 5886 147978
rect 5942 147922 36234 147978
rect 36290 147922 36358 147978
rect 36414 147922 36482 147978
rect 36538 147922 36606 147978
rect 36662 147922 66954 147978
rect 67010 147922 67078 147978
rect 67134 147922 67202 147978
rect 67258 147922 67326 147978
rect 67382 147922 97674 147978
rect 97730 147922 97798 147978
rect 97854 147922 97922 147978
rect 97978 147922 98046 147978
rect 98102 147922 128394 147978
rect 128450 147922 128518 147978
rect 128574 147922 128642 147978
rect 128698 147922 128766 147978
rect 128822 147922 159114 147978
rect 159170 147922 159238 147978
rect 159294 147922 159362 147978
rect 159418 147922 159486 147978
rect 159542 147922 189834 147978
rect 189890 147922 189958 147978
rect 190014 147922 190082 147978
rect 190138 147922 190206 147978
rect 190262 147922 220554 147978
rect 220610 147922 220678 147978
rect 220734 147922 220802 147978
rect 220858 147922 220926 147978
rect 220982 147922 251274 147978
rect 251330 147922 251398 147978
rect 251454 147922 251522 147978
rect 251578 147922 251646 147978
rect 251702 147922 281994 147978
rect 282050 147922 282118 147978
rect 282174 147922 282242 147978
rect 282298 147922 282366 147978
rect 282422 147922 312714 147978
rect 312770 147922 312838 147978
rect 312894 147922 312962 147978
rect 313018 147922 313086 147978
rect 313142 147922 343434 147978
rect 343490 147922 343558 147978
rect 343614 147922 343682 147978
rect 343738 147922 343806 147978
rect 343862 147922 374154 147978
rect 374210 147922 374278 147978
rect 374334 147922 374402 147978
rect 374458 147922 374526 147978
rect 374582 147922 404874 147978
rect 404930 147922 404998 147978
rect 405054 147922 405122 147978
rect 405178 147922 405246 147978
rect 405302 147922 435594 147978
rect 435650 147922 435718 147978
rect 435774 147922 435842 147978
rect 435898 147922 435966 147978
rect 436022 147922 466314 147978
rect 466370 147922 466438 147978
rect 466494 147922 466562 147978
rect 466618 147922 466686 147978
rect 466742 147922 497034 147978
rect 497090 147922 497158 147978
rect 497214 147922 497282 147978
rect 497338 147922 497406 147978
rect 497462 147922 527754 147978
rect 527810 147922 527878 147978
rect 527934 147922 528002 147978
rect 528058 147922 528126 147978
rect 528182 147922 558474 147978
rect 558530 147922 558598 147978
rect 558654 147922 558722 147978
rect 558778 147922 558846 147978
rect 558902 147922 589194 147978
rect 589250 147922 589318 147978
rect 589374 147922 589442 147978
rect 589498 147922 589566 147978
rect 589622 147922 596496 147978
rect 596552 147922 596620 147978
rect 596676 147922 596744 147978
rect 596800 147922 596868 147978
rect 596924 147922 597980 147978
rect -1916 147826 597980 147922
rect -1916 136350 597980 136446
rect -1916 136294 -1820 136350
rect -1764 136294 -1696 136350
rect -1640 136294 -1572 136350
rect -1516 136294 -1448 136350
rect -1392 136294 9234 136350
rect 9290 136294 9358 136350
rect 9414 136294 9482 136350
rect 9538 136294 9606 136350
rect 9662 136294 39954 136350
rect 40010 136294 40078 136350
rect 40134 136294 40202 136350
rect 40258 136294 40326 136350
rect 40382 136294 70674 136350
rect 70730 136294 70798 136350
rect 70854 136294 70922 136350
rect 70978 136294 71046 136350
rect 71102 136294 101394 136350
rect 101450 136294 101518 136350
rect 101574 136294 101642 136350
rect 101698 136294 101766 136350
rect 101822 136294 132114 136350
rect 132170 136294 132238 136350
rect 132294 136294 132362 136350
rect 132418 136294 132486 136350
rect 132542 136294 162834 136350
rect 162890 136294 162958 136350
rect 163014 136294 163082 136350
rect 163138 136294 163206 136350
rect 163262 136294 193554 136350
rect 193610 136294 193678 136350
rect 193734 136294 193802 136350
rect 193858 136294 193926 136350
rect 193982 136294 224274 136350
rect 224330 136294 224398 136350
rect 224454 136294 224522 136350
rect 224578 136294 224646 136350
rect 224702 136294 254994 136350
rect 255050 136294 255118 136350
rect 255174 136294 255242 136350
rect 255298 136294 255366 136350
rect 255422 136294 285714 136350
rect 285770 136294 285838 136350
rect 285894 136294 285962 136350
rect 286018 136294 286086 136350
rect 286142 136294 316434 136350
rect 316490 136294 316558 136350
rect 316614 136294 316682 136350
rect 316738 136294 316806 136350
rect 316862 136294 347154 136350
rect 347210 136294 347278 136350
rect 347334 136294 347402 136350
rect 347458 136294 347526 136350
rect 347582 136294 377874 136350
rect 377930 136294 377998 136350
rect 378054 136294 378122 136350
rect 378178 136294 378246 136350
rect 378302 136294 408594 136350
rect 408650 136294 408718 136350
rect 408774 136294 408842 136350
rect 408898 136294 408966 136350
rect 409022 136294 439314 136350
rect 439370 136294 439438 136350
rect 439494 136294 439562 136350
rect 439618 136294 439686 136350
rect 439742 136294 470034 136350
rect 470090 136294 470158 136350
rect 470214 136294 470282 136350
rect 470338 136294 470406 136350
rect 470462 136294 500754 136350
rect 500810 136294 500878 136350
rect 500934 136294 501002 136350
rect 501058 136294 501126 136350
rect 501182 136294 531474 136350
rect 531530 136294 531598 136350
rect 531654 136294 531722 136350
rect 531778 136294 531846 136350
rect 531902 136294 562194 136350
rect 562250 136294 562318 136350
rect 562374 136294 562442 136350
rect 562498 136294 562566 136350
rect 562622 136294 592914 136350
rect 592970 136294 593038 136350
rect 593094 136294 593162 136350
rect 593218 136294 593286 136350
rect 593342 136294 597456 136350
rect 597512 136294 597580 136350
rect 597636 136294 597704 136350
rect 597760 136294 597828 136350
rect 597884 136294 597980 136350
rect -1916 136226 597980 136294
rect -1916 136170 -1820 136226
rect -1764 136170 -1696 136226
rect -1640 136170 -1572 136226
rect -1516 136170 -1448 136226
rect -1392 136170 9234 136226
rect 9290 136170 9358 136226
rect 9414 136170 9482 136226
rect 9538 136170 9606 136226
rect 9662 136170 39954 136226
rect 40010 136170 40078 136226
rect 40134 136170 40202 136226
rect 40258 136170 40326 136226
rect 40382 136170 70674 136226
rect 70730 136170 70798 136226
rect 70854 136170 70922 136226
rect 70978 136170 71046 136226
rect 71102 136170 101394 136226
rect 101450 136170 101518 136226
rect 101574 136170 101642 136226
rect 101698 136170 101766 136226
rect 101822 136170 132114 136226
rect 132170 136170 132238 136226
rect 132294 136170 132362 136226
rect 132418 136170 132486 136226
rect 132542 136170 162834 136226
rect 162890 136170 162958 136226
rect 163014 136170 163082 136226
rect 163138 136170 163206 136226
rect 163262 136170 193554 136226
rect 193610 136170 193678 136226
rect 193734 136170 193802 136226
rect 193858 136170 193926 136226
rect 193982 136170 224274 136226
rect 224330 136170 224398 136226
rect 224454 136170 224522 136226
rect 224578 136170 224646 136226
rect 224702 136170 254994 136226
rect 255050 136170 255118 136226
rect 255174 136170 255242 136226
rect 255298 136170 255366 136226
rect 255422 136170 285714 136226
rect 285770 136170 285838 136226
rect 285894 136170 285962 136226
rect 286018 136170 286086 136226
rect 286142 136170 316434 136226
rect 316490 136170 316558 136226
rect 316614 136170 316682 136226
rect 316738 136170 316806 136226
rect 316862 136170 347154 136226
rect 347210 136170 347278 136226
rect 347334 136170 347402 136226
rect 347458 136170 347526 136226
rect 347582 136170 377874 136226
rect 377930 136170 377998 136226
rect 378054 136170 378122 136226
rect 378178 136170 378246 136226
rect 378302 136170 408594 136226
rect 408650 136170 408718 136226
rect 408774 136170 408842 136226
rect 408898 136170 408966 136226
rect 409022 136170 439314 136226
rect 439370 136170 439438 136226
rect 439494 136170 439562 136226
rect 439618 136170 439686 136226
rect 439742 136170 470034 136226
rect 470090 136170 470158 136226
rect 470214 136170 470282 136226
rect 470338 136170 470406 136226
rect 470462 136170 500754 136226
rect 500810 136170 500878 136226
rect 500934 136170 501002 136226
rect 501058 136170 501126 136226
rect 501182 136170 531474 136226
rect 531530 136170 531598 136226
rect 531654 136170 531722 136226
rect 531778 136170 531846 136226
rect 531902 136170 562194 136226
rect 562250 136170 562318 136226
rect 562374 136170 562442 136226
rect 562498 136170 562566 136226
rect 562622 136170 592914 136226
rect 592970 136170 593038 136226
rect 593094 136170 593162 136226
rect 593218 136170 593286 136226
rect 593342 136170 597456 136226
rect 597512 136170 597580 136226
rect 597636 136170 597704 136226
rect 597760 136170 597828 136226
rect 597884 136170 597980 136226
rect -1916 136102 597980 136170
rect -1916 136046 -1820 136102
rect -1764 136046 -1696 136102
rect -1640 136046 -1572 136102
rect -1516 136046 -1448 136102
rect -1392 136046 9234 136102
rect 9290 136046 9358 136102
rect 9414 136046 9482 136102
rect 9538 136046 9606 136102
rect 9662 136046 39954 136102
rect 40010 136046 40078 136102
rect 40134 136046 40202 136102
rect 40258 136046 40326 136102
rect 40382 136046 70674 136102
rect 70730 136046 70798 136102
rect 70854 136046 70922 136102
rect 70978 136046 71046 136102
rect 71102 136046 101394 136102
rect 101450 136046 101518 136102
rect 101574 136046 101642 136102
rect 101698 136046 101766 136102
rect 101822 136046 132114 136102
rect 132170 136046 132238 136102
rect 132294 136046 132362 136102
rect 132418 136046 132486 136102
rect 132542 136046 162834 136102
rect 162890 136046 162958 136102
rect 163014 136046 163082 136102
rect 163138 136046 163206 136102
rect 163262 136046 193554 136102
rect 193610 136046 193678 136102
rect 193734 136046 193802 136102
rect 193858 136046 193926 136102
rect 193982 136046 224274 136102
rect 224330 136046 224398 136102
rect 224454 136046 224522 136102
rect 224578 136046 224646 136102
rect 224702 136046 254994 136102
rect 255050 136046 255118 136102
rect 255174 136046 255242 136102
rect 255298 136046 255366 136102
rect 255422 136046 285714 136102
rect 285770 136046 285838 136102
rect 285894 136046 285962 136102
rect 286018 136046 286086 136102
rect 286142 136046 316434 136102
rect 316490 136046 316558 136102
rect 316614 136046 316682 136102
rect 316738 136046 316806 136102
rect 316862 136046 347154 136102
rect 347210 136046 347278 136102
rect 347334 136046 347402 136102
rect 347458 136046 347526 136102
rect 347582 136046 377874 136102
rect 377930 136046 377998 136102
rect 378054 136046 378122 136102
rect 378178 136046 378246 136102
rect 378302 136046 408594 136102
rect 408650 136046 408718 136102
rect 408774 136046 408842 136102
rect 408898 136046 408966 136102
rect 409022 136046 439314 136102
rect 439370 136046 439438 136102
rect 439494 136046 439562 136102
rect 439618 136046 439686 136102
rect 439742 136046 470034 136102
rect 470090 136046 470158 136102
rect 470214 136046 470282 136102
rect 470338 136046 470406 136102
rect 470462 136046 500754 136102
rect 500810 136046 500878 136102
rect 500934 136046 501002 136102
rect 501058 136046 501126 136102
rect 501182 136046 531474 136102
rect 531530 136046 531598 136102
rect 531654 136046 531722 136102
rect 531778 136046 531846 136102
rect 531902 136046 562194 136102
rect 562250 136046 562318 136102
rect 562374 136046 562442 136102
rect 562498 136046 562566 136102
rect 562622 136046 592914 136102
rect 592970 136046 593038 136102
rect 593094 136046 593162 136102
rect 593218 136046 593286 136102
rect 593342 136046 597456 136102
rect 597512 136046 597580 136102
rect 597636 136046 597704 136102
rect 597760 136046 597828 136102
rect 597884 136046 597980 136102
rect -1916 135978 597980 136046
rect -1916 135922 -1820 135978
rect -1764 135922 -1696 135978
rect -1640 135922 -1572 135978
rect -1516 135922 -1448 135978
rect -1392 135922 9234 135978
rect 9290 135922 9358 135978
rect 9414 135922 9482 135978
rect 9538 135922 9606 135978
rect 9662 135922 39954 135978
rect 40010 135922 40078 135978
rect 40134 135922 40202 135978
rect 40258 135922 40326 135978
rect 40382 135922 70674 135978
rect 70730 135922 70798 135978
rect 70854 135922 70922 135978
rect 70978 135922 71046 135978
rect 71102 135922 101394 135978
rect 101450 135922 101518 135978
rect 101574 135922 101642 135978
rect 101698 135922 101766 135978
rect 101822 135922 132114 135978
rect 132170 135922 132238 135978
rect 132294 135922 132362 135978
rect 132418 135922 132486 135978
rect 132542 135922 162834 135978
rect 162890 135922 162958 135978
rect 163014 135922 163082 135978
rect 163138 135922 163206 135978
rect 163262 135922 193554 135978
rect 193610 135922 193678 135978
rect 193734 135922 193802 135978
rect 193858 135922 193926 135978
rect 193982 135922 224274 135978
rect 224330 135922 224398 135978
rect 224454 135922 224522 135978
rect 224578 135922 224646 135978
rect 224702 135922 254994 135978
rect 255050 135922 255118 135978
rect 255174 135922 255242 135978
rect 255298 135922 255366 135978
rect 255422 135922 285714 135978
rect 285770 135922 285838 135978
rect 285894 135922 285962 135978
rect 286018 135922 286086 135978
rect 286142 135922 316434 135978
rect 316490 135922 316558 135978
rect 316614 135922 316682 135978
rect 316738 135922 316806 135978
rect 316862 135922 347154 135978
rect 347210 135922 347278 135978
rect 347334 135922 347402 135978
rect 347458 135922 347526 135978
rect 347582 135922 377874 135978
rect 377930 135922 377998 135978
rect 378054 135922 378122 135978
rect 378178 135922 378246 135978
rect 378302 135922 408594 135978
rect 408650 135922 408718 135978
rect 408774 135922 408842 135978
rect 408898 135922 408966 135978
rect 409022 135922 439314 135978
rect 439370 135922 439438 135978
rect 439494 135922 439562 135978
rect 439618 135922 439686 135978
rect 439742 135922 470034 135978
rect 470090 135922 470158 135978
rect 470214 135922 470282 135978
rect 470338 135922 470406 135978
rect 470462 135922 500754 135978
rect 500810 135922 500878 135978
rect 500934 135922 501002 135978
rect 501058 135922 501126 135978
rect 501182 135922 531474 135978
rect 531530 135922 531598 135978
rect 531654 135922 531722 135978
rect 531778 135922 531846 135978
rect 531902 135922 562194 135978
rect 562250 135922 562318 135978
rect 562374 135922 562442 135978
rect 562498 135922 562566 135978
rect 562622 135922 592914 135978
rect 592970 135922 593038 135978
rect 593094 135922 593162 135978
rect 593218 135922 593286 135978
rect 593342 135922 597456 135978
rect 597512 135922 597580 135978
rect 597636 135922 597704 135978
rect 597760 135922 597828 135978
rect 597884 135922 597980 135978
rect -1916 135826 597980 135922
rect -1916 130350 597980 130446
rect -1916 130294 -860 130350
rect -804 130294 -736 130350
rect -680 130294 -612 130350
rect -556 130294 -488 130350
rect -432 130294 5514 130350
rect 5570 130294 5638 130350
rect 5694 130294 5762 130350
rect 5818 130294 5886 130350
rect 5942 130294 36234 130350
rect 36290 130294 36358 130350
rect 36414 130294 36482 130350
rect 36538 130294 36606 130350
rect 36662 130294 66954 130350
rect 67010 130294 67078 130350
rect 67134 130294 67202 130350
rect 67258 130294 67326 130350
rect 67382 130294 97674 130350
rect 97730 130294 97798 130350
rect 97854 130294 97922 130350
rect 97978 130294 98046 130350
rect 98102 130294 128394 130350
rect 128450 130294 128518 130350
rect 128574 130294 128642 130350
rect 128698 130294 128766 130350
rect 128822 130294 159114 130350
rect 159170 130294 159238 130350
rect 159294 130294 159362 130350
rect 159418 130294 159486 130350
rect 159542 130294 189834 130350
rect 189890 130294 189958 130350
rect 190014 130294 190082 130350
rect 190138 130294 190206 130350
rect 190262 130294 220554 130350
rect 220610 130294 220678 130350
rect 220734 130294 220802 130350
rect 220858 130294 220926 130350
rect 220982 130294 251274 130350
rect 251330 130294 251398 130350
rect 251454 130294 251522 130350
rect 251578 130294 251646 130350
rect 251702 130294 281994 130350
rect 282050 130294 282118 130350
rect 282174 130294 282242 130350
rect 282298 130294 282366 130350
rect 282422 130294 312714 130350
rect 312770 130294 312838 130350
rect 312894 130294 312962 130350
rect 313018 130294 313086 130350
rect 313142 130294 343434 130350
rect 343490 130294 343558 130350
rect 343614 130294 343682 130350
rect 343738 130294 343806 130350
rect 343862 130294 374154 130350
rect 374210 130294 374278 130350
rect 374334 130294 374402 130350
rect 374458 130294 374526 130350
rect 374582 130294 404874 130350
rect 404930 130294 404998 130350
rect 405054 130294 405122 130350
rect 405178 130294 405246 130350
rect 405302 130294 435594 130350
rect 435650 130294 435718 130350
rect 435774 130294 435842 130350
rect 435898 130294 435966 130350
rect 436022 130294 466314 130350
rect 466370 130294 466438 130350
rect 466494 130294 466562 130350
rect 466618 130294 466686 130350
rect 466742 130294 497034 130350
rect 497090 130294 497158 130350
rect 497214 130294 497282 130350
rect 497338 130294 497406 130350
rect 497462 130294 527754 130350
rect 527810 130294 527878 130350
rect 527934 130294 528002 130350
rect 528058 130294 528126 130350
rect 528182 130294 558474 130350
rect 558530 130294 558598 130350
rect 558654 130294 558722 130350
rect 558778 130294 558846 130350
rect 558902 130294 589194 130350
rect 589250 130294 589318 130350
rect 589374 130294 589442 130350
rect 589498 130294 589566 130350
rect 589622 130294 596496 130350
rect 596552 130294 596620 130350
rect 596676 130294 596744 130350
rect 596800 130294 596868 130350
rect 596924 130294 597980 130350
rect -1916 130226 597980 130294
rect -1916 130170 -860 130226
rect -804 130170 -736 130226
rect -680 130170 -612 130226
rect -556 130170 -488 130226
rect -432 130170 5514 130226
rect 5570 130170 5638 130226
rect 5694 130170 5762 130226
rect 5818 130170 5886 130226
rect 5942 130170 36234 130226
rect 36290 130170 36358 130226
rect 36414 130170 36482 130226
rect 36538 130170 36606 130226
rect 36662 130170 66954 130226
rect 67010 130170 67078 130226
rect 67134 130170 67202 130226
rect 67258 130170 67326 130226
rect 67382 130170 97674 130226
rect 97730 130170 97798 130226
rect 97854 130170 97922 130226
rect 97978 130170 98046 130226
rect 98102 130170 128394 130226
rect 128450 130170 128518 130226
rect 128574 130170 128642 130226
rect 128698 130170 128766 130226
rect 128822 130170 159114 130226
rect 159170 130170 159238 130226
rect 159294 130170 159362 130226
rect 159418 130170 159486 130226
rect 159542 130170 189834 130226
rect 189890 130170 189958 130226
rect 190014 130170 190082 130226
rect 190138 130170 190206 130226
rect 190262 130170 220554 130226
rect 220610 130170 220678 130226
rect 220734 130170 220802 130226
rect 220858 130170 220926 130226
rect 220982 130170 251274 130226
rect 251330 130170 251398 130226
rect 251454 130170 251522 130226
rect 251578 130170 251646 130226
rect 251702 130170 281994 130226
rect 282050 130170 282118 130226
rect 282174 130170 282242 130226
rect 282298 130170 282366 130226
rect 282422 130170 312714 130226
rect 312770 130170 312838 130226
rect 312894 130170 312962 130226
rect 313018 130170 313086 130226
rect 313142 130170 343434 130226
rect 343490 130170 343558 130226
rect 343614 130170 343682 130226
rect 343738 130170 343806 130226
rect 343862 130170 374154 130226
rect 374210 130170 374278 130226
rect 374334 130170 374402 130226
rect 374458 130170 374526 130226
rect 374582 130170 404874 130226
rect 404930 130170 404998 130226
rect 405054 130170 405122 130226
rect 405178 130170 405246 130226
rect 405302 130170 435594 130226
rect 435650 130170 435718 130226
rect 435774 130170 435842 130226
rect 435898 130170 435966 130226
rect 436022 130170 466314 130226
rect 466370 130170 466438 130226
rect 466494 130170 466562 130226
rect 466618 130170 466686 130226
rect 466742 130170 497034 130226
rect 497090 130170 497158 130226
rect 497214 130170 497282 130226
rect 497338 130170 497406 130226
rect 497462 130170 527754 130226
rect 527810 130170 527878 130226
rect 527934 130170 528002 130226
rect 528058 130170 528126 130226
rect 528182 130170 558474 130226
rect 558530 130170 558598 130226
rect 558654 130170 558722 130226
rect 558778 130170 558846 130226
rect 558902 130170 589194 130226
rect 589250 130170 589318 130226
rect 589374 130170 589442 130226
rect 589498 130170 589566 130226
rect 589622 130170 596496 130226
rect 596552 130170 596620 130226
rect 596676 130170 596744 130226
rect 596800 130170 596868 130226
rect 596924 130170 597980 130226
rect -1916 130102 597980 130170
rect -1916 130046 -860 130102
rect -804 130046 -736 130102
rect -680 130046 -612 130102
rect -556 130046 -488 130102
rect -432 130046 5514 130102
rect 5570 130046 5638 130102
rect 5694 130046 5762 130102
rect 5818 130046 5886 130102
rect 5942 130046 36234 130102
rect 36290 130046 36358 130102
rect 36414 130046 36482 130102
rect 36538 130046 36606 130102
rect 36662 130046 66954 130102
rect 67010 130046 67078 130102
rect 67134 130046 67202 130102
rect 67258 130046 67326 130102
rect 67382 130046 97674 130102
rect 97730 130046 97798 130102
rect 97854 130046 97922 130102
rect 97978 130046 98046 130102
rect 98102 130046 128394 130102
rect 128450 130046 128518 130102
rect 128574 130046 128642 130102
rect 128698 130046 128766 130102
rect 128822 130046 159114 130102
rect 159170 130046 159238 130102
rect 159294 130046 159362 130102
rect 159418 130046 159486 130102
rect 159542 130046 189834 130102
rect 189890 130046 189958 130102
rect 190014 130046 190082 130102
rect 190138 130046 190206 130102
rect 190262 130046 220554 130102
rect 220610 130046 220678 130102
rect 220734 130046 220802 130102
rect 220858 130046 220926 130102
rect 220982 130046 251274 130102
rect 251330 130046 251398 130102
rect 251454 130046 251522 130102
rect 251578 130046 251646 130102
rect 251702 130046 281994 130102
rect 282050 130046 282118 130102
rect 282174 130046 282242 130102
rect 282298 130046 282366 130102
rect 282422 130046 312714 130102
rect 312770 130046 312838 130102
rect 312894 130046 312962 130102
rect 313018 130046 313086 130102
rect 313142 130046 343434 130102
rect 343490 130046 343558 130102
rect 343614 130046 343682 130102
rect 343738 130046 343806 130102
rect 343862 130046 374154 130102
rect 374210 130046 374278 130102
rect 374334 130046 374402 130102
rect 374458 130046 374526 130102
rect 374582 130046 404874 130102
rect 404930 130046 404998 130102
rect 405054 130046 405122 130102
rect 405178 130046 405246 130102
rect 405302 130046 435594 130102
rect 435650 130046 435718 130102
rect 435774 130046 435842 130102
rect 435898 130046 435966 130102
rect 436022 130046 466314 130102
rect 466370 130046 466438 130102
rect 466494 130046 466562 130102
rect 466618 130046 466686 130102
rect 466742 130046 497034 130102
rect 497090 130046 497158 130102
rect 497214 130046 497282 130102
rect 497338 130046 497406 130102
rect 497462 130046 527754 130102
rect 527810 130046 527878 130102
rect 527934 130046 528002 130102
rect 528058 130046 528126 130102
rect 528182 130046 558474 130102
rect 558530 130046 558598 130102
rect 558654 130046 558722 130102
rect 558778 130046 558846 130102
rect 558902 130046 589194 130102
rect 589250 130046 589318 130102
rect 589374 130046 589442 130102
rect 589498 130046 589566 130102
rect 589622 130046 596496 130102
rect 596552 130046 596620 130102
rect 596676 130046 596744 130102
rect 596800 130046 596868 130102
rect 596924 130046 597980 130102
rect -1916 129978 597980 130046
rect -1916 129922 -860 129978
rect -804 129922 -736 129978
rect -680 129922 -612 129978
rect -556 129922 -488 129978
rect -432 129922 5514 129978
rect 5570 129922 5638 129978
rect 5694 129922 5762 129978
rect 5818 129922 5886 129978
rect 5942 129922 36234 129978
rect 36290 129922 36358 129978
rect 36414 129922 36482 129978
rect 36538 129922 36606 129978
rect 36662 129922 66954 129978
rect 67010 129922 67078 129978
rect 67134 129922 67202 129978
rect 67258 129922 67326 129978
rect 67382 129922 97674 129978
rect 97730 129922 97798 129978
rect 97854 129922 97922 129978
rect 97978 129922 98046 129978
rect 98102 129922 128394 129978
rect 128450 129922 128518 129978
rect 128574 129922 128642 129978
rect 128698 129922 128766 129978
rect 128822 129922 159114 129978
rect 159170 129922 159238 129978
rect 159294 129922 159362 129978
rect 159418 129922 159486 129978
rect 159542 129922 189834 129978
rect 189890 129922 189958 129978
rect 190014 129922 190082 129978
rect 190138 129922 190206 129978
rect 190262 129922 220554 129978
rect 220610 129922 220678 129978
rect 220734 129922 220802 129978
rect 220858 129922 220926 129978
rect 220982 129922 251274 129978
rect 251330 129922 251398 129978
rect 251454 129922 251522 129978
rect 251578 129922 251646 129978
rect 251702 129922 281994 129978
rect 282050 129922 282118 129978
rect 282174 129922 282242 129978
rect 282298 129922 282366 129978
rect 282422 129922 312714 129978
rect 312770 129922 312838 129978
rect 312894 129922 312962 129978
rect 313018 129922 313086 129978
rect 313142 129922 343434 129978
rect 343490 129922 343558 129978
rect 343614 129922 343682 129978
rect 343738 129922 343806 129978
rect 343862 129922 374154 129978
rect 374210 129922 374278 129978
rect 374334 129922 374402 129978
rect 374458 129922 374526 129978
rect 374582 129922 404874 129978
rect 404930 129922 404998 129978
rect 405054 129922 405122 129978
rect 405178 129922 405246 129978
rect 405302 129922 435594 129978
rect 435650 129922 435718 129978
rect 435774 129922 435842 129978
rect 435898 129922 435966 129978
rect 436022 129922 466314 129978
rect 466370 129922 466438 129978
rect 466494 129922 466562 129978
rect 466618 129922 466686 129978
rect 466742 129922 497034 129978
rect 497090 129922 497158 129978
rect 497214 129922 497282 129978
rect 497338 129922 497406 129978
rect 497462 129922 527754 129978
rect 527810 129922 527878 129978
rect 527934 129922 528002 129978
rect 528058 129922 528126 129978
rect 528182 129922 558474 129978
rect 558530 129922 558598 129978
rect 558654 129922 558722 129978
rect 558778 129922 558846 129978
rect 558902 129922 589194 129978
rect 589250 129922 589318 129978
rect 589374 129922 589442 129978
rect 589498 129922 589566 129978
rect 589622 129922 596496 129978
rect 596552 129922 596620 129978
rect 596676 129922 596744 129978
rect 596800 129922 596868 129978
rect 596924 129922 597980 129978
rect -1916 129826 597980 129922
rect -1916 118350 597980 118446
rect -1916 118294 -1820 118350
rect -1764 118294 -1696 118350
rect -1640 118294 -1572 118350
rect -1516 118294 -1448 118350
rect -1392 118294 9234 118350
rect 9290 118294 9358 118350
rect 9414 118294 9482 118350
rect 9538 118294 9606 118350
rect 9662 118294 39954 118350
rect 40010 118294 40078 118350
rect 40134 118294 40202 118350
rect 40258 118294 40326 118350
rect 40382 118294 70674 118350
rect 70730 118294 70798 118350
rect 70854 118294 70922 118350
rect 70978 118294 71046 118350
rect 71102 118294 101394 118350
rect 101450 118294 101518 118350
rect 101574 118294 101642 118350
rect 101698 118294 101766 118350
rect 101822 118294 132114 118350
rect 132170 118294 132238 118350
rect 132294 118294 132362 118350
rect 132418 118294 132486 118350
rect 132542 118294 162834 118350
rect 162890 118294 162958 118350
rect 163014 118294 163082 118350
rect 163138 118294 163206 118350
rect 163262 118294 193554 118350
rect 193610 118294 193678 118350
rect 193734 118294 193802 118350
rect 193858 118294 193926 118350
rect 193982 118294 224274 118350
rect 224330 118294 224398 118350
rect 224454 118294 224522 118350
rect 224578 118294 224646 118350
rect 224702 118294 254994 118350
rect 255050 118294 255118 118350
rect 255174 118294 255242 118350
rect 255298 118294 255366 118350
rect 255422 118294 285714 118350
rect 285770 118294 285838 118350
rect 285894 118294 285962 118350
rect 286018 118294 286086 118350
rect 286142 118294 316434 118350
rect 316490 118294 316558 118350
rect 316614 118294 316682 118350
rect 316738 118294 316806 118350
rect 316862 118294 347154 118350
rect 347210 118294 347278 118350
rect 347334 118294 347402 118350
rect 347458 118294 347526 118350
rect 347582 118294 377874 118350
rect 377930 118294 377998 118350
rect 378054 118294 378122 118350
rect 378178 118294 378246 118350
rect 378302 118294 408594 118350
rect 408650 118294 408718 118350
rect 408774 118294 408842 118350
rect 408898 118294 408966 118350
rect 409022 118294 439314 118350
rect 439370 118294 439438 118350
rect 439494 118294 439562 118350
rect 439618 118294 439686 118350
rect 439742 118294 470034 118350
rect 470090 118294 470158 118350
rect 470214 118294 470282 118350
rect 470338 118294 470406 118350
rect 470462 118294 500754 118350
rect 500810 118294 500878 118350
rect 500934 118294 501002 118350
rect 501058 118294 501126 118350
rect 501182 118294 531474 118350
rect 531530 118294 531598 118350
rect 531654 118294 531722 118350
rect 531778 118294 531846 118350
rect 531902 118294 562194 118350
rect 562250 118294 562318 118350
rect 562374 118294 562442 118350
rect 562498 118294 562566 118350
rect 562622 118294 592914 118350
rect 592970 118294 593038 118350
rect 593094 118294 593162 118350
rect 593218 118294 593286 118350
rect 593342 118294 597456 118350
rect 597512 118294 597580 118350
rect 597636 118294 597704 118350
rect 597760 118294 597828 118350
rect 597884 118294 597980 118350
rect -1916 118226 597980 118294
rect -1916 118170 -1820 118226
rect -1764 118170 -1696 118226
rect -1640 118170 -1572 118226
rect -1516 118170 -1448 118226
rect -1392 118170 9234 118226
rect 9290 118170 9358 118226
rect 9414 118170 9482 118226
rect 9538 118170 9606 118226
rect 9662 118170 39954 118226
rect 40010 118170 40078 118226
rect 40134 118170 40202 118226
rect 40258 118170 40326 118226
rect 40382 118170 70674 118226
rect 70730 118170 70798 118226
rect 70854 118170 70922 118226
rect 70978 118170 71046 118226
rect 71102 118170 101394 118226
rect 101450 118170 101518 118226
rect 101574 118170 101642 118226
rect 101698 118170 101766 118226
rect 101822 118170 132114 118226
rect 132170 118170 132238 118226
rect 132294 118170 132362 118226
rect 132418 118170 132486 118226
rect 132542 118170 162834 118226
rect 162890 118170 162958 118226
rect 163014 118170 163082 118226
rect 163138 118170 163206 118226
rect 163262 118170 193554 118226
rect 193610 118170 193678 118226
rect 193734 118170 193802 118226
rect 193858 118170 193926 118226
rect 193982 118170 224274 118226
rect 224330 118170 224398 118226
rect 224454 118170 224522 118226
rect 224578 118170 224646 118226
rect 224702 118170 254994 118226
rect 255050 118170 255118 118226
rect 255174 118170 255242 118226
rect 255298 118170 255366 118226
rect 255422 118170 285714 118226
rect 285770 118170 285838 118226
rect 285894 118170 285962 118226
rect 286018 118170 286086 118226
rect 286142 118170 316434 118226
rect 316490 118170 316558 118226
rect 316614 118170 316682 118226
rect 316738 118170 316806 118226
rect 316862 118170 347154 118226
rect 347210 118170 347278 118226
rect 347334 118170 347402 118226
rect 347458 118170 347526 118226
rect 347582 118170 377874 118226
rect 377930 118170 377998 118226
rect 378054 118170 378122 118226
rect 378178 118170 378246 118226
rect 378302 118170 408594 118226
rect 408650 118170 408718 118226
rect 408774 118170 408842 118226
rect 408898 118170 408966 118226
rect 409022 118170 439314 118226
rect 439370 118170 439438 118226
rect 439494 118170 439562 118226
rect 439618 118170 439686 118226
rect 439742 118170 470034 118226
rect 470090 118170 470158 118226
rect 470214 118170 470282 118226
rect 470338 118170 470406 118226
rect 470462 118170 500754 118226
rect 500810 118170 500878 118226
rect 500934 118170 501002 118226
rect 501058 118170 501126 118226
rect 501182 118170 531474 118226
rect 531530 118170 531598 118226
rect 531654 118170 531722 118226
rect 531778 118170 531846 118226
rect 531902 118170 562194 118226
rect 562250 118170 562318 118226
rect 562374 118170 562442 118226
rect 562498 118170 562566 118226
rect 562622 118170 592914 118226
rect 592970 118170 593038 118226
rect 593094 118170 593162 118226
rect 593218 118170 593286 118226
rect 593342 118170 597456 118226
rect 597512 118170 597580 118226
rect 597636 118170 597704 118226
rect 597760 118170 597828 118226
rect 597884 118170 597980 118226
rect -1916 118102 597980 118170
rect -1916 118046 -1820 118102
rect -1764 118046 -1696 118102
rect -1640 118046 -1572 118102
rect -1516 118046 -1448 118102
rect -1392 118046 9234 118102
rect 9290 118046 9358 118102
rect 9414 118046 9482 118102
rect 9538 118046 9606 118102
rect 9662 118046 39954 118102
rect 40010 118046 40078 118102
rect 40134 118046 40202 118102
rect 40258 118046 40326 118102
rect 40382 118046 70674 118102
rect 70730 118046 70798 118102
rect 70854 118046 70922 118102
rect 70978 118046 71046 118102
rect 71102 118046 101394 118102
rect 101450 118046 101518 118102
rect 101574 118046 101642 118102
rect 101698 118046 101766 118102
rect 101822 118046 132114 118102
rect 132170 118046 132238 118102
rect 132294 118046 132362 118102
rect 132418 118046 132486 118102
rect 132542 118046 162834 118102
rect 162890 118046 162958 118102
rect 163014 118046 163082 118102
rect 163138 118046 163206 118102
rect 163262 118046 193554 118102
rect 193610 118046 193678 118102
rect 193734 118046 193802 118102
rect 193858 118046 193926 118102
rect 193982 118046 224274 118102
rect 224330 118046 224398 118102
rect 224454 118046 224522 118102
rect 224578 118046 224646 118102
rect 224702 118046 254994 118102
rect 255050 118046 255118 118102
rect 255174 118046 255242 118102
rect 255298 118046 255366 118102
rect 255422 118046 285714 118102
rect 285770 118046 285838 118102
rect 285894 118046 285962 118102
rect 286018 118046 286086 118102
rect 286142 118046 316434 118102
rect 316490 118046 316558 118102
rect 316614 118046 316682 118102
rect 316738 118046 316806 118102
rect 316862 118046 347154 118102
rect 347210 118046 347278 118102
rect 347334 118046 347402 118102
rect 347458 118046 347526 118102
rect 347582 118046 377874 118102
rect 377930 118046 377998 118102
rect 378054 118046 378122 118102
rect 378178 118046 378246 118102
rect 378302 118046 408594 118102
rect 408650 118046 408718 118102
rect 408774 118046 408842 118102
rect 408898 118046 408966 118102
rect 409022 118046 439314 118102
rect 439370 118046 439438 118102
rect 439494 118046 439562 118102
rect 439618 118046 439686 118102
rect 439742 118046 470034 118102
rect 470090 118046 470158 118102
rect 470214 118046 470282 118102
rect 470338 118046 470406 118102
rect 470462 118046 500754 118102
rect 500810 118046 500878 118102
rect 500934 118046 501002 118102
rect 501058 118046 501126 118102
rect 501182 118046 531474 118102
rect 531530 118046 531598 118102
rect 531654 118046 531722 118102
rect 531778 118046 531846 118102
rect 531902 118046 562194 118102
rect 562250 118046 562318 118102
rect 562374 118046 562442 118102
rect 562498 118046 562566 118102
rect 562622 118046 592914 118102
rect 592970 118046 593038 118102
rect 593094 118046 593162 118102
rect 593218 118046 593286 118102
rect 593342 118046 597456 118102
rect 597512 118046 597580 118102
rect 597636 118046 597704 118102
rect 597760 118046 597828 118102
rect 597884 118046 597980 118102
rect -1916 117978 597980 118046
rect -1916 117922 -1820 117978
rect -1764 117922 -1696 117978
rect -1640 117922 -1572 117978
rect -1516 117922 -1448 117978
rect -1392 117922 9234 117978
rect 9290 117922 9358 117978
rect 9414 117922 9482 117978
rect 9538 117922 9606 117978
rect 9662 117922 39954 117978
rect 40010 117922 40078 117978
rect 40134 117922 40202 117978
rect 40258 117922 40326 117978
rect 40382 117922 70674 117978
rect 70730 117922 70798 117978
rect 70854 117922 70922 117978
rect 70978 117922 71046 117978
rect 71102 117922 101394 117978
rect 101450 117922 101518 117978
rect 101574 117922 101642 117978
rect 101698 117922 101766 117978
rect 101822 117922 132114 117978
rect 132170 117922 132238 117978
rect 132294 117922 132362 117978
rect 132418 117922 132486 117978
rect 132542 117922 162834 117978
rect 162890 117922 162958 117978
rect 163014 117922 163082 117978
rect 163138 117922 163206 117978
rect 163262 117922 193554 117978
rect 193610 117922 193678 117978
rect 193734 117922 193802 117978
rect 193858 117922 193926 117978
rect 193982 117922 224274 117978
rect 224330 117922 224398 117978
rect 224454 117922 224522 117978
rect 224578 117922 224646 117978
rect 224702 117922 254994 117978
rect 255050 117922 255118 117978
rect 255174 117922 255242 117978
rect 255298 117922 255366 117978
rect 255422 117922 285714 117978
rect 285770 117922 285838 117978
rect 285894 117922 285962 117978
rect 286018 117922 286086 117978
rect 286142 117922 316434 117978
rect 316490 117922 316558 117978
rect 316614 117922 316682 117978
rect 316738 117922 316806 117978
rect 316862 117922 347154 117978
rect 347210 117922 347278 117978
rect 347334 117922 347402 117978
rect 347458 117922 347526 117978
rect 347582 117922 377874 117978
rect 377930 117922 377998 117978
rect 378054 117922 378122 117978
rect 378178 117922 378246 117978
rect 378302 117922 408594 117978
rect 408650 117922 408718 117978
rect 408774 117922 408842 117978
rect 408898 117922 408966 117978
rect 409022 117922 439314 117978
rect 439370 117922 439438 117978
rect 439494 117922 439562 117978
rect 439618 117922 439686 117978
rect 439742 117922 470034 117978
rect 470090 117922 470158 117978
rect 470214 117922 470282 117978
rect 470338 117922 470406 117978
rect 470462 117922 500754 117978
rect 500810 117922 500878 117978
rect 500934 117922 501002 117978
rect 501058 117922 501126 117978
rect 501182 117922 531474 117978
rect 531530 117922 531598 117978
rect 531654 117922 531722 117978
rect 531778 117922 531846 117978
rect 531902 117922 562194 117978
rect 562250 117922 562318 117978
rect 562374 117922 562442 117978
rect 562498 117922 562566 117978
rect 562622 117922 592914 117978
rect 592970 117922 593038 117978
rect 593094 117922 593162 117978
rect 593218 117922 593286 117978
rect 593342 117922 597456 117978
rect 597512 117922 597580 117978
rect 597636 117922 597704 117978
rect 597760 117922 597828 117978
rect 597884 117922 597980 117978
rect -1916 117826 597980 117922
rect -1916 112350 597980 112446
rect -1916 112294 -860 112350
rect -804 112294 -736 112350
rect -680 112294 -612 112350
rect -556 112294 -488 112350
rect -432 112294 5514 112350
rect 5570 112294 5638 112350
rect 5694 112294 5762 112350
rect 5818 112294 5886 112350
rect 5942 112294 36234 112350
rect 36290 112294 36358 112350
rect 36414 112294 36482 112350
rect 36538 112294 36606 112350
rect 36662 112294 66954 112350
rect 67010 112294 67078 112350
rect 67134 112294 67202 112350
rect 67258 112294 67326 112350
rect 67382 112294 97674 112350
rect 97730 112294 97798 112350
rect 97854 112294 97922 112350
rect 97978 112294 98046 112350
rect 98102 112294 128394 112350
rect 128450 112294 128518 112350
rect 128574 112294 128642 112350
rect 128698 112294 128766 112350
rect 128822 112294 159114 112350
rect 159170 112294 159238 112350
rect 159294 112294 159362 112350
rect 159418 112294 159486 112350
rect 159542 112294 189834 112350
rect 189890 112294 189958 112350
rect 190014 112294 190082 112350
rect 190138 112294 190206 112350
rect 190262 112294 220554 112350
rect 220610 112294 220678 112350
rect 220734 112294 220802 112350
rect 220858 112294 220926 112350
rect 220982 112294 251274 112350
rect 251330 112294 251398 112350
rect 251454 112294 251522 112350
rect 251578 112294 251646 112350
rect 251702 112294 281994 112350
rect 282050 112294 282118 112350
rect 282174 112294 282242 112350
rect 282298 112294 282366 112350
rect 282422 112294 312714 112350
rect 312770 112294 312838 112350
rect 312894 112294 312962 112350
rect 313018 112294 313086 112350
rect 313142 112294 343434 112350
rect 343490 112294 343558 112350
rect 343614 112294 343682 112350
rect 343738 112294 343806 112350
rect 343862 112294 374154 112350
rect 374210 112294 374278 112350
rect 374334 112294 374402 112350
rect 374458 112294 374526 112350
rect 374582 112294 404874 112350
rect 404930 112294 404998 112350
rect 405054 112294 405122 112350
rect 405178 112294 405246 112350
rect 405302 112294 435594 112350
rect 435650 112294 435718 112350
rect 435774 112294 435842 112350
rect 435898 112294 435966 112350
rect 436022 112294 466314 112350
rect 466370 112294 466438 112350
rect 466494 112294 466562 112350
rect 466618 112294 466686 112350
rect 466742 112294 497034 112350
rect 497090 112294 497158 112350
rect 497214 112294 497282 112350
rect 497338 112294 497406 112350
rect 497462 112294 527754 112350
rect 527810 112294 527878 112350
rect 527934 112294 528002 112350
rect 528058 112294 528126 112350
rect 528182 112294 558474 112350
rect 558530 112294 558598 112350
rect 558654 112294 558722 112350
rect 558778 112294 558846 112350
rect 558902 112294 589194 112350
rect 589250 112294 589318 112350
rect 589374 112294 589442 112350
rect 589498 112294 589566 112350
rect 589622 112294 596496 112350
rect 596552 112294 596620 112350
rect 596676 112294 596744 112350
rect 596800 112294 596868 112350
rect 596924 112294 597980 112350
rect -1916 112226 597980 112294
rect -1916 112170 -860 112226
rect -804 112170 -736 112226
rect -680 112170 -612 112226
rect -556 112170 -488 112226
rect -432 112170 5514 112226
rect 5570 112170 5638 112226
rect 5694 112170 5762 112226
rect 5818 112170 5886 112226
rect 5942 112170 36234 112226
rect 36290 112170 36358 112226
rect 36414 112170 36482 112226
rect 36538 112170 36606 112226
rect 36662 112170 66954 112226
rect 67010 112170 67078 112226
rect 67134 112170 67202 112226
rect 67258 112170 67326 112226
rect 67382 112170 97674 112226
rect 97730 112170 97798 112226
rect 97854 112170 97922 112226
rect 97978 112170 98046 112226
rect 98102 112170 128394 112226
rect 128450 112170 128518 112226
rect 128574 112170 128642 112226
rect 128698 112170 128766 112226
rect 128822 112170 159114 112226
rect 159170 112170 159238 112226
rect 159294 112170 159362 112226
rect 159418 112170 159486 112226
rect 159542 112170 189834 112226
rect 189890 112170 189958 112226
rect 190014 112170 190082 112226
rect 190138 112170 190206 112226
rect 190262 112170 220554 112226
rect 220610 112170 220678 112226
rect 220734 112170 220802 112226
rect 220858 112170 220926 112226
rect 220982 112170 251274 112226
rect 251330 112170 251398 112226
rect 251454 112170 251522 112226
rect 251578 112170 251646 112226
rect 251702 112170 281994 112226
rect 282050 112170 282118 112226
rect 282174 112170 282242 112226
rect 282298 112170 282366 112226
rect 282422 112170 312714 112226
rect 312770 112170 312838 112226
rect 312894 112170 312962 112226
rect 313018 112170 313086 112226
rect 313142 112170 343434 112226
rect 343490 112170 343558 112226
rect 343614 112170 343682 112226
rect 343738 112170 343806 112226
rect 343862 112170 374154 112226
rect 374210 112170 374278 112226
rect 374334 112170 374402 112226
rect 374458 112170 374526 112226
rect 374582 112170 404874 112226
rect 404930 112170 404998 112226
rect 405054 112170 405122 112226
rect 405178 112170 405246 112226
rect 405302 112170 435594 112226
rect 435650 112170 435718 112226
rect 435774 112170 435842 112226
rect 435898 112170 435966 112226
rect 436022 112170 466314 112226
rect 466370 112170 466438 112226
rect 466494 112170 466562 112226
rect 466618 112170 466686 112226
rect 466742 112170 497034 112226
rect 497090 112170 497158 112226
rect 497214 112170 497282 112226
rect 497338 112170 497406 112226
rect 497462 112170 527754 112226
rect 527810 112170 527878 112226
rect 527934 112170 528002 112226
rect 528058 112170 528126 112226
rect 528182 112170 558474 112226
rect 558530 112170 558598 112226
rect 558654 112170 558722 112226
rect 558778 112170 558846 112226
rect 558902 112170 589194 112226
rect 589250 112170 589318 112226
rect 589374 112170 589442 112226
rect 589498 112170 589566 112226
rect 589622 112170 596496 112226
rect 596552 112170 596620 112226
rect 596676 112170 596744 112226
rect 596800 112170 596868 112226
rect 596924 112170 597980 112226
rect -1916 112102 597980 112170
rect -1916 112046 -860 112102
rect -804 112046 -736 112102
rect -680 112046 -612 112102
rect -556 112046 -488 112102
rect -432 112046 5514 112102
rect 5570 112046 5638 112102
rect 5694 112046 5762 112102
rect 5818 112046 5886 112102
rect 5942 112046 36234 112102
rect 36290 112046 36358 112102
rect 36414 112046 36482 112102
rect 36538 112046 36606 112102
rect 36662 112046 66954 112102
rect 67010 112046 67078 112102
rect 67134 112046 67202 112102
rect 67258 112046 67326 112102
rect 67382 112046 97674 112102
rect 97730 112046 97798 112102
rect 97854 112046 97922 112102
rect 97978 112046 98046 112102
rect 98102 112046 128394 112102
rect 128450 112046 128518 112102
rect 128574 112046 128642 112102
rect 128698 112046 128766 112102
rect 128822 112046 159114 112102
rect 159170 112046 159238 112102
rect 159294 112046 159362 112102
rect 159418 112046 159486 112102
rect 159542 112046 189834 112102
rect 189890 112046 189958 112102
rect 190014 112046 190082 112102
rect 190138 112046 190206 112102
rect 190262 112046 220554 112102
rect 220610 112046 220678 112102
rect 220734 112046 220802 112102
rect 220858 112046 220926 112102
rect 220982 112046 251274 112102
rect 251330 112046 251398 112102
rect 251454 112046 251522 112102
rect 251578 112046 251646 112102
rect 251702 112046 281994 112102
rect 282050 112046 282118 112102
rect 282174 112046 282242 112102
rect 282298 112046 282366 112102
rect 282422 112046 312714 112102
rect 312770 112046 312838 112102
rect 312894 112046 312962 112102
rect 313018 112046 313086 112102
rect 313142 112046 343434 112102
rect 343490 112046 343558 112102
rect 343614 112046 343682 112102
rect 343738 112046 343806 112102
rect 343862 112046 374154 112102
rect 374210 112046 374278 112102
rect 374334 112046 374402 112102
rect 374458 112046 374526 112102
rect 374582 112046 404874 112102
rect 404930 112046 404998 112102
rect 405054 112046 405122 112102
rect 405178 112046 405246 112102
rect 405302 112046 435594 112102
rect 435650 112046 435718 112102
rect 435774 112046 435842 112102
rect 435898 112046 435966 112102
rect 436022 112046 466314 112102
rect 466370 112046 466438 112102
rect 466494 112046 466562 112102
rect 466618 112046 466686 112102
rect 466742 112046 497034 112102
rect 497090 112046 497158 112102
rect 497214 112046 497282 112102
rect 497338 112046 497406 112102
rect 497462 112046 527754 112102
rect 527810 112046 527878 112102
rect 527934 112046 528002 112102
rect 528058 112046 528126 112102
rect 528182 112046 558474 112102
rect 558530 112046 558598 112102
rect 558654 112046 558722 112102
rect 558778 112046 558846 112102
rect 558902 112046 589194 112102
rect 589250 112046 589318 112102
rect 589374 112046 589442 112102
rect 589498 112046 589566 112102
rect 589622 112046 596496 112102
rect 596552 112046 596620 112102
rect 596676 112046 596744 112102
rect 596800 112046 596868 112102
rect 596924 112046 597980 112102
rect -1916 111978 597980 112046
rect -1916 111922 -860 111978
rect -804 111922 -736 111978
rect -680 111922 -612 111978
rect -556 111922 -488 111978
rect -432 111922 5514 111978
rect 5570 111922 5638 111978
rect 5694 111922 5762 111978
rect 5818 111922 5886 111978
rect 5942 111922 36234 111978
rect 36290 111922 36358 111978
rect 36414 111922 36482 111978
rect 36538 111922 36606 111978
rect 36662 111922 66954 111978
rect 67010 111922 67078 111978
rect 67134 111922 67202 111978
rect 67258 111922 67326 111978
rect 67382 111922 97674 111978
rect 97730 111922 97798 111978
rect 97854 111922 97922 111978
rect 97978 111922 98046 111978
rect 98102 111922 128394 111978
rect 128450 111922 128518 111978
rect 128574 111922 128642 111978
rect 128698 111922 128766 111978
rect 128822 111922 159114 111978
rect 159170 111922 159238 111978
rect 159294 111922 159362 111978
rect 159418 111922 159486 111978
rect 159542 111922 189834 111978
rect 189890 111922 189958 111978
rect 190014 111922 190082 111978
rect 190138 111922 190206 111978
rect 190262 111922 220554 111978
rect 220610 111922 220678 111978
rect 220734 111922 220802 111978
rect 220858 111922 220926 111978
rect 220982 111922 251274 111978
rect 251330 111922 251398 111978
rect 251454 111922 251522 111978
rect 251578 111922 251646 111978
rect 251702 111922 281994 111978
rect 282050 111922 282118 111978
rect 282174 111922 282242 111978
rect 282298 111922 282366 111978
rect 282422 111922 312714 111978
rect 312770 111922 312838 111978
rect 312894 111922 312962 111978
rect 313018 111922 313086 111978
rect 313142 111922 343434 111978
rect 343490 111922 343558 111978
rect 343614 111922 343682 111978
rect 343738 111922 343806 111978
rect 343862 111922 374154 111978
rect 374210 111922 374278 111978
rect 374334 111922 374402 111978
rect 374458 111922 374526 111978
rect 374582 111922 404874 111978
rect 404930 111922 404998 111978
rect 405054 111922 405122 111978
rect 405178 111922 405246 111978
rect 405302 111922 435594 111978
rect 435650 111922 435718 111978
rect 435774 111922 435842 111978
rect 435898 111922 435966 111978
rect 436022 111922 466314 111978
rect 466370 111922 466438 111978
rect 466494 111922 466562 111978
rect 466618 111922 466686 111978
rect 466742 111922 497034 111978
rect 497090 111922 497158 111978
rect 497214 111922 497282 111978
rect 497338 111922 497406 111978
rect 497462 111922 527754 111978
rect 527810 111922 527878 111978
rect 527934 111922 528002 111978
rect 528058 111922 528126 111978
rect 528182 111922 558474 111978
rect 558530 111922 558598 111978
rect 558654 111922 558722 111978
rect 558778 111922 558846 111978
rect 558902 111922 589194 111978
rect 589250 111922 589318 111978
rect 589374 111922 589442 111978
rect 589498 111922 589566 111978
rect 589622 111922 596496 111978
rect 596552 111922 596620 111978
rect 596676 111922 596744 111978
rect 596800 111922 596868 111978
rect 596924 111922 597980 111978
rect -1916 111826 597980 111922
rect -1916 100350 597980 100446
rect -1916 100294 -1820 100350
rect -1764 100294 -1696 100350
rect -1640 100294 -1572 100350
rect -1516 100294 -1448 100350
rect -1392 100294 9234 100350
rect 9290 100294 9358 100350
rect 9414 100294 9482 100350
rect 9538 100294 9606 100350
rect 9662 100294 39954 100350
rect 40010 100294 40078 100350
rect 40134 100294 40202 100350
rect 40258 100294 40326 100350
rect 40382 100294 70674 100350
rect 70730 100294 70798 100350
rect 70854 100294 70922 100350
rect 70978 100294 71046 100350
rect 71102 100294 101394 100350
rect 101450 100294 101518 100350
rect 101574 100294 101642 100350
rect 101698 100294 101766 100350
rect 101822 100294 132114 100350
rect 132170 100294 132238 100350
rect 132294 100294 132362 100350
rect 132418 100294 132486 100350
rect 132542 100294 162834 100350
rect 162890 100294 162958 100350
rect 163014 100294 163082 100350
rect 163138 100294 163206 100350
rect 163262 100294 193554 100350
rect 193610 100294 193678 100350
rect 193734 100294 193802 100350
rect 193858 100294 193926 100350
rect 193982 100294 224274 100350
rect 224330 100294 224398 100350
rect 224454 100294 224522 100350
rect 224578 100294 224646 100350
rect 224702 100294 254994 100350
rect 255050 100294 255118 100350
rect 255174 100294 255242 100350
rect 255298 100294 255366 100350
rect 255422 100294 285714 100350
rect 285770 100294 285838 100350
rect 285894 100294 285962 100350
rect 286018 100294 286086 100350
rect 286142 100294 316434 100350
rect 316490 100294 316558 100350
rect 316614 100294 316682 100350
rect 316738 100294 316806 100350
rect 316862 100294 347154 100350
rect 347210 100294 347278 100350
rect 347334 100294 347402 100350
rect 347458 100294 347526 100350
rect 347582 100294 377874 100350
rect 377930 100294 377998 100350
rect 378054 100294 378122 100350
rect 378178 100294 378246 100350
rect 378302 100294 408594 100350
rect 408650 100294 408718 100350
rect 408774 100294 408842 100350
rect 408898 100294 408966 100350
rect 409022 100294 439314 100350
rect 439370 100294 439438 100350
rect 439494 100294 439562 100350
rect 439618 100294 439686 100350
rect 439742 100294 470034 100350
rect 470090 100294 470158 100350
rect 470214 100294 470282 100350
rect 470338 100294 470406 100350
rect 470462 100294 500754 100350
rect 500810 100294 500878 100350
rect 500934 100294 501002 100350
rect 501058 100294 501126 100350
rect 501182 100294 531474 100350
rect 531530 100294 531598 100350
rect 531654 100294 531722 100350
rect 531778 100294 531846 100350
rect 531902 100294 562194 100350
rect 562250 100294 562318 100350
rect 562374 100294 562442 100350
rect 562498 100294 562566 100350
rect 562622 100294 592914 100350
rect 592970 100294 593038 100350
rect 593094 100294 593162 100350
rect 593218 100294 593286 100350
rect 593342 100294 597456 100350
rect 597512 100294 597580 100350
rect 597636 100294 597704 100350
rect 597760 100294 597828 100350
rect 597884 100294 597980 100350
rect -1916 100226 597980 100294
rect -1916 100170 -1820 100226
rect -1764 100170 -1696 100226
rect -1640 100170 -1572 100226
rect -1516 100170 -1448 100226
rect -1392 100170 9234 100226
rect 9290 100170 9358 100226
rect 9414 100170 9482 100226
rect 9538 100170 9606 100226
rect 9662 100170 39954 100226
rect 40010 100170 40078 100226
rect 40134 100170 40202 100226
rect 40258 100170 40326 100226
rect 40382 100170 70674 100226
rect 70730 100170 70798 100226
rect 70854 100170 70922 100226
rect 70978 100170 71046 100226
rect 71102 100170 101394 100226
rect 101450 100170 101518 100226
rect 101574 100170 101642 100226
rect 101698 100170 101766 100226
rect 101822 100170 132114 100226
rect 132170 100170 132238 100226
rect 132294 100170 132362 100226
rect 132418 100170 132486 100226
rect 132542 100170 162834 100226
rect 162890 100170 162958 100226
rect 163014 100170 163082 100226
rect 163138 100170 163206 100226
rect 163262 100170 193554 100226
rect 193610 100170 193678 100226
rect 193734 100170 193802 100226
rect 193858 100170 193926 100226
rect 193982 100170 224274 100226
rect 224330 100170 224398 100226
rect 224454 100170 224522 100226
rect 224578 100170 224646 100226
rect 224702 100170 254994 100226
rect 255050 100170 255118 100226
rect 255174 100170 255242 100226
rect 255298 100170 255366 100226
rect 255422 100170 285714 100226
rect 285770 100170 285838 100226
rect 285894 100170 285962 100226
rect 286018 100170 286086 100226
rect 286142 100170 316434 100226
rect 316490 100170 316558 100226
rect 316614 100170 316682 100226
rect 316738 100170 316806 100226
rect 316862 100170 347154 100226
rect 347210 100170 347278 100226
rect 347334 100170 347402 100226
rect 347458 100170 347526 100226
rect 347582 100170 377874 100226
rect 377930 100170 377998 100226
rect 378054 100170 378122 100226
rect 378178 100170 378246 100226
rect 378302 100170 408594 100226
rect 408650 100170 408718 100226
rect 408774 100170 408842 100226
rect 408898 100170 408966 100226
rect 409022 100170 439314 100226
rect 439370 100170 439438 100226
rect 439494 100170 439562 100226
rect 439618 100170 439686 100226
rect 439742 100170 470034 100226
rect 470090 100170 470158 100226
rect 470214 100170 470282 100226
rect 470338 100170 470406 100226
rect 470462 100170 500754 100226
rect 500810 100170 500878 100226
rect 500934 100170 501002 100226
rect 501058 100170 501126 100226
rect 501182 100170 531474 100226
rect 531530 100170 531598 100226
rect 531654 100170 531722 100226
rect 531778 100170 531846 100226
rect 531902 100170 562194 100226
rect 562250 100170 562318 100226
rect 562374 100170 562442 100226
rect 562498 100170 562566 100226
rect 562622 100170 592914 100226
rect 592970 100170 593038 100226
rect 593094 100170 593162 100226
rect 593218 100170 593286 100226
rect 593342 100170 597456 100226
rect 597512 100170 597580 100226
rect 597636 100170 597704 100226
rect 597760 100170 597828 100226
rect 597884 100170 597980 100226
rect -1916 100102 597980 100170
rect -1916 100046 -1820 100102
rect -1764 100046 -1696 100102
rect -1640 100046 -1572 100102
rect -1516 100046 -1448 100102
rect -1392 100046 9234 100102
rect 9290 100046 9358 100102
rect 9414 100046 9482 100102
rect 9538 100046 9606 100102
rect 9662 100046 39954 100102
rect 40010 100046 40078 100102
rect 40134 100046 40202 100102
rect 40258 100046 40326 100102
rect 40382 100046 70674 100102
rect 70730 100046 70798 100102
rect 70854 100046 70922 100102
rect 70978 100046 71046 100102
rect 71102 100046 101394 100102
rect 101450 100046 101518 100102
rect 101574 100046 101642 100102
rect 101698 100046 101766 100102
rect 101822 100046 132114 100102
rect 132170 100046 132238 100102
rect 132294 100046 132362 100102
rect 132418 100046 132486 100102
rect 132542 100046 162834 100102
rect 162890 100046 162958 100102
rect 163014 100046 163082 100102
rect 163138 100046 163206 100102
rect 163262 100046 193554 100102
rect 193610 100046 193678 100102
rect 193734 100046 193802 100102
rect 193858 100046 193926 100102
rect 193982 100046 224274 100102
rect 224330 100046 224398 100102
rect 224454 100046 224522 100102
rect 224578 100046 224646 100102
rect 224702 100046 254994 100102
rect 255050 100046 255118 100102
rect 255174 100046 255242 100102
rect 255298 100046 255366 100102
rect 255422 100046 285714 100102
rect 285770 100046 285838 100102
rect 285894 100046 285962 100102
rect 286018 100046 286086 100102
rect 286142 100046 316434 100102
rect 316490 100046 316558 100102
rect 316614 100046 316682 100102
rect 316738 100046 316806 100102
rect 316862 100046 347154 100102
rect 347210 100046 347278 100102
rect 347334 100046 347402 100102
rect 347458 100046 347526 100102
rect 347582 100046 377874 100102
rect 377930 100046 377998 100102
rect 378054 100046 378122 100102
rect 378178 100046 378246 100102
rect 378302 100046 408594 100102
rect 408650 100046 408718 100102
rect 408774 100046 408842 100102
rect 408898 100046 408966 100102
rect 409022 100046 439314 100102
rect 439370 100046 439438 100102
rect 439494 100046 439562 100102
rect 439618 100046 439686 100102
rect 439742 100046 470034 100102
rect 470090 100046 470158 100102
rect 470214 100046 470282 100102
rect 470338 100046 470406 100102
rect 470462 100046 500754 100102
rect 500810 100046 500878 100102
rect 500934 100046 501002 100102
rect 501058 100046 501126 100102
rect 501182 100046 531474 100102
rect 531530 100046 531598 100102
rect 531654 100046 531722 100102
rect 531778 100046 531846 100102
rect 531902 100046 562194 100102
rect 562250 100046 562318 100102
rect 562374 100046 562442 100102
rect 562498 100046 562566 100102
rect 562622 100046 592914 100102
rect 592970 100046 593038 100102
rect 593094 100046 593162 100102
rect 593218 100046 593286 100102
rect 593342 100046 597456 100102
rect 597512 100046 597580 100102
rect 597636 100046 597704 100102
rect 597760 100046 597828 100102
rect 597884 100046 597980 100102
rect -1916 99978 597980 100046
rect -1916 99922 -1820 99978
rect -1764 99922 -1696 99978
rect -1640 99922 -1572 99978
rect -1516 99922 -1448 99978
rect -1392 99922 9234 99978
rect 9290 99922 9358 99978
rect 9414 99922 9482 99978
rect 9538 99922 9606 99978
rect 9662 99922 39954 99978
rect 40010 99922 40078 99978
rect 40134 99922 40202 99978
rect 40258 99922 40326 99978
rect 40382 99922 70674 99978
rect 70730 99922 70798 99978
rect 70854 99922 70922 99978
rect 70978 99922 71046 99978
rect 71102 99922 101394 99978
rect 101450 99922 101518 99978
rect 101574 99922 101642 99978
rect 101698 99922 101766 99978
rect 101822 99922 132114 99978
rect 132170 99922 132238 99978
rect 132294 99922 132362 99978
rect 132418 99922 132486 99978
rect 132542 99922 162834 99978
rect 162890 99922 162958 99978
rect 163014 99922 163082 99978
rect 163138 99922 163206 99978
rect 163262 99922 193554 99978
rect 193610 99922 193678 99978
rect 193734 99922 193802 99978
rect 193858 99922 193926 99978
rect 193982 99922 224274 99978
rect 224330 99922 224398 99978
rect 224454 99922 224522 99978
rect 224578 99922 224646 99978
rect 224702 99922 254994 99978
rect 255050 99922 255118 99978
rect 255174 99922 255242 99978
rect 255298 99922 255366 99978
rect 255422 99922 285714 99978
rect 285770 99922 285838 99978
rect 285894 99922 285962 99978
rect 286018 99922 286086 99978
rect 286142 99922 316434 99978
rect 316490 99922 316558 99978
rect 316614 99922 316682 99978
rect 316738 99922 316806 99978
rect 316862 99922 347154 99978
rect 347210 99922 347278 99978
rect 347334 99922 347402 99978
rect 347458 99922 347526 99978
rect 347582 99922 377874 99978
rect 377930 99922 377998 99978
rect 378054 99922 378122 99978
rect 378178 99922 378246 99978
rect 378302 99922 408594 99978
rect 408650 99922 408718 99978
rect 408774 99922 408842 99978
rect 408898 99922 408966 99978
rect 409022 99922 439314 99978
rect 439370 99922 439438 99978
rect 439494 99922 439562 99978
rect 439618 99922 439686 99978
rect 439742 99922 470034 99978
rect 470090 99922 470158 99978
rect 470214 99922 470282 99978
rect 470338 99922 470406 99978
rect 470462 99922 500754 99978
rect 500810 99922 500878 99978
rect 500934 99922 501002 99978
rect 501058 99922 501126 99978
rect 501182 99922 531474 99978
rect 531530 99922 531598 99978
rect 531654 99922 531722 99978
rect 531778 99922 531846 99978
rect 531902 99922 562194 99978
rect 562250 99922 562318 99978
rect 562374 99922 562442 99978
rect 562498 99922 562566 99978
rect 562622 99922 592914 99978
rect 592970 99922 593038 99978
rect 593094 99922 593162 99978
rect 593218 99922 593286 99978
rect 593342 99922 597456 99978
rect 597512 99922 597580 99978
rect 597636 99922 597704 99978
rect 597760 99922 597828 99978
rect 597884 99922 597980 99978
rect -1916 99826 597980 99922
rect -1916 94350 597980 94446
rect -1916 94294 -860 94350
rect -804 94294 -736 94350
rect -680 94294 -612 94350
rect -556 94294 -488 94350
rect -432 94294 5514 94350
rect 5570 94294 5638 94350
rect 5694 94294 5762 94350
rect 5818 94294 5886 94350
rect 5942 94294 36234 94350
rect 36290 94294 36358 94350
rect 36414 94294 36482 94350
rect 36538 94294 36606 94350
rect 36662 94294 66954 94350
rect 67010 94294 67078 94350
rect 67134 94294 67202 94350
rect 67258 94294 67326 94350
rect 67382 94294 97674 94350
rect 97730 94294 97798 94350
rect 97854 94294 97922 94350
rect 97978 94294 98046 94350
rect 98102 94294 128394 94350
rect 128450 94294 128518 94350
rect 128574 94294 128642 94350
rect 128698 94294 128766 94350
rect 128822 94294 159114 94350
rect 159170 94294 159238 94350
rect 159294 94294 159362 94350
rect 159418 94294 159486 94350
rect 159542 94294 189834 94350
rect 189890 94294 189958 94350
rect 190014 94294 190082 94350
rect 190138 94294 190206 94350
rect 190262 94294 220554 94350
rect 220610 94294 220678 94350
rect 220734 94294 220802 94350
rect 220858 94294 220926 94350
rect 220982 94294 251274 94350
rect 251330 94294 251398 94350
rect 251454 94294 251522 94350
rect 251578 94294 251646 94350
rect 251702 94294 281994 94350
rect 282050 94294 282118 94350
rect 282174 94294 282242 94350
rect 282298 94294 282366 94350
rect 282422 94294 312714 94350
rect 312770 94294 312838 94350
rect 312894 94294 312962 94350
rect 313018 94294 313086 94350
rect 313142 94294 343434 94350
rect 343490 94294 343558 94350
rect 343614 94294 343682 94350
rect 343738 94294 343806 94350
rect 343862 94294 374154 94350
rect 374210 94294 374278 94350
rect 374334 94294 374402 94350
rect 374458 94294 374526 94350
rect 374582 94294 404874 94350
rect 404930 94294 404998 94350
rect 405054 94294 405122 94350
rect 405178 94294 405246 94350
rect 405302 94294 435594 94350
rect 435650 94294 435718 94350
rect 435774 94294 435842 94350
rect 435898 94294 435966 94350
rect 436022 94294 466314 94350
rect 466370 94294 466438 94350
rect 466494 94294 466562 94350
rect 466618 94294 466686 94350
rect 466742 94294 497034 94350
rect 497090 94294 497158 94350
rect 497214 94294 497282 94350
rect 497338 94294 497406 94350
rect 497462 94294 527754 94350
rect 527810 94294 527878 94350
rect 527934 94294 528002 94350
rect 528058 94294 528126 94350
rect 528182 94294 558474 94350
rect 558530 94294 558598 94350
rect 558654 94294 558722 94350
rect 558778 94294 558846 94350
rect 558902 94294 589194 94350
rect 589250 94294 589318 94350
rect 589374 94294 589442 94350
rect 589498 94294 589566 94350
rect 589622 94294 596496 94350
rect 596552 94294 596620 94350
rect 596676 94294 596744 94350
rect 596800 94294 596868 94350
rect 596924 94294 597980 94350
rect -1916 94226 597980 94294
rect -1916 94170 -860 94226
rect -804 94170 -736 94226
rect -680 94170 -612 94226
rect -556 94170 -488 94226
rect -432 94170 5514 94226
rect 5570 94170 5638 94226
rect 5694 94170 5762 94226
rect 5818 94170 5886 94226
rect 5942 94170 36234 94226
rect 36290 94170 36358 94226
rect 36414 94170 36482 94226
rect 36538 94170 36606 94226
rect 36662 94170 66954 94226
rect 67010 94170 67078 94226
rect 67134 94170 67202 94226
rect 67258 94170 67326 94226
rect 67382 94170 97674 94226
rect 97730 94170 97798 94226
rect 97854 94170 97922 94226
rect 97978 94170 98046 94226
rect 98102 94170 128394 94226
rect 128450 94170 128518 94226
rect 128574 94170 128642 94226
rect 128698 94170 128766 94226
rect 128822 94170 159114 94226
rect 159170 94170 159238 94226
rect 159294 94170 159362 94226
rect 159418 94170 159486 94226
rect 159542 94170 189834 94226
rect 189890 94170 189958 94226
rect 190014 94170 190082 94226
rect 190138 94170 190206 94226
rect 190262 94170 220554 94226
rect 220610 94170 220678 94226
rect 220734 94170 220802 94226
rect 220858 94170 220926 94226
rect 220982 94170 251274 94226
rect 251330 94170 251398 94226
rect 251454 94170 251522 94226
rect 251578 94170 251646 94226
rect 251702 94170 281994 94226
rect 282050 94170 282118 94226
rect 282174 94170 282242 94226
rect 282298 94170 282366 94226
rect 282422 94170 312714 94226
rect 312770 94170 312838 94226
rect 312894 94170 312962 94226
rect 313018 94170 313086 94226
rect 313142 94170 343434 94226
rect 343490 94170 343558 94226
rect 343614 94170 343682 94226
rect 343738 94170 343806 94226
rect 343862 94170 374154 94226
rect 374210 94170 374278 94226
rect 374334 94170 374402 94226
rect 374458 94170 374526 94226
rect 374582 94170 404874 94226
rect 404930 94170 404998 94226
rect 405054 94170 405122 94226
rect 405178 94170 405246 94226
rect 405302 94170 435594 94226
rect 435650 94170 435718 94226
rect 435774 94170 435842 94226
rect 435898 94170 435966 94226
rect 436022 94170 466314 94226
rect 466370 94170 466438 94226
rect 466494 94170 466562 94226
rect 466618 94170 466686 94226
rect 466742 94170 497034 94226
rect 497090 94170 497158 94226
rect 497214 94170 497282 94226
rect 497338 94170 497406 94226
rect 497462 94170 527754 94226
rect 527810 94170 527878 94226
rect 527934 94170 528002 94226
rect 528058 94170 528126 94226
rect 528182 94170 558474 94226
rect 558530 94170 558598 94226
rect 558654 94170 558722 94226
rect 558778 94170 558846 94226
rect 558902 94170 589194 94226
rect 589250 94170 589318 94226
rect 589374 94170 589442 94226
rect 589498 94170 589566 94226
rect 589622 94170 596496 94226
rect 596552 94170 596620 94226
rect 596676 94170 596744 94226
rect 596800 94170 596868 94226
rect 596924 94170 597980 94226
rect -1916 94102 597980 94170
rect -1916 94046 -860 94102
rect -804 94046 -736 94102
rect -680 94046 -612 94102
rect -556 94046 -488 94102
rect -432 94046 5514 94102
rect 5570 94046 5638 94102
rect 5694 94046 5762 94102
rect 5818 94046 5886 94102
rect 5942 94046 36234 94102
rect 36290 94046 36358 94102
rect 36414 94046 36482 94102
rect 36538 94046 36606 94102
rect 36662 94046 66954 94102
rect 67010 94046 67078 94102
rect 67134 94046 67202 94102
rect 67258 94046 67326 94102
rect 67382 94046 97674 94102
rect 97730 94046 97798 94102
rect 97854 94046 97922 94102
rect 97978 94046 98046 94102
rect 98102 94046 128394 94102
rect 128450 94046 128518 94102
rect 128574 94046 128642 94102
rect 128698 94046 128766 94102
rect 128822 94046 159114 94102
rect 159170 94046 159238 94102
rect 159294 94046 159362 94102
rect 159418 94046 159486 94102
rect 159542 94046 189834 94102
rect 189890 94046 189958 94102
rect 190014 94046 190082 94102
rect 190138 94046 190206 94102
rect 190262 94046 220554 94102
rect 220610 94046 220678 94102
rect 220734 94046 220802 94102
rect 220858 94046 220926 94102
rect 220982 94046 251274 94102
rect 251330 94046 251398 94102
rect 251454 94046 251522 94102
rect 251578 94046 251646 94102
rect 251702 94046 281994 94102
rect 282050 94046 282118 94102
rect 282174 94046 282242 94102
rect 282298 94046 282366 94102
rect 282422 94046 312714 94102
rect 312770 94046 312838 94102
rect 312894 94046 312962 94102
rect 313018 94046 313086 94102
rect 313142 94046 343434 94102
rect 343490 94046 343558 94102
rect 343614 94046 343682 94102
rect 343738 94046 343806 94102
rect 343862 94046 374154 94102
rect 374210 94046 374278 94102
rect 374334 94046 374402 94102
rect 374458 94046 374526 94102
rect 374582 94046 404874 94102
rect 404930 94046 404998 94102
rect 405054 94046 405122 94102
rect 405178 94046 405246 94102
rect 405302 94046 435594 94102
rect 435650 94046 435718 94102
rect 435774 94046 435842 94102
rect 435898 94046 435966 94102
rect 436022 94046 466314 94102
rect 466370 94046 466438 94102
rect 466494 94046 466562 94102
rect 466618 94046 466686 94102
rect 466742 94046 497034 94102
rect 497090 94046 497158 94102
rect 497214 94046 497282 94102
rect 497338 94046 497406 94102
rect 497462 94046 527754 94102
rect 527810 94046 527878 94102
rect 527934 94046 528002 94102
rect 528058 94046 528126 94102
rect 528182 94046 558474 94102
rect 558530 94046 558598 94102
rect 558654 94046 558722 94102
rect 558778 94046 558846 94102
rect 558902 94046 589194 94102
rect 589250 94046 589318 94102
rect 589374 94046 589442 94102
rect 589498 94046 589566 94102
rect 589622 94046 596496 94102
rect 596552 94046 596620 94102
rect 596676 94046 596744 94102
rect 596800 94046 596868 94102
rect 596924 94046 597980 94102
rect -1916 93978 597980 94046
rect -1916 93922 -860 93978
rect -804 93922 -736 93978
rect -680 93922 -612 93978
rect -556 93922 -488 93978
rect -432 93922 5514 93978
rect 5570 93922 5638 93978
rect 5694 93922 5762 93978
rect 5818 93922 5886 93978
rect 5942 93922 36234 93978
rect 36290 93922 36358 93978
rect 36414 93922 36482 93978
rect 36538 93922 36606 93978
rect 36662 93922 66954 93978
rect 67010 93922 67078 93978
rect 67134 93922 67202 93978
rect 67258 93922 67326 93978
rect 67382 93922 97674 93978
rect 97730 93922 97798 93978
rect 97854 93922 97922 93978
rect 97978 93922 98046 93978
rect 98102 93922 128394 93978
rect 128450 93922 128518 93978
rect 128574 93922 128642 93978
rect 128698 93922 128766 93978
rect 128822 93922 159114 93978
rect 159170 93922 159238 93978
rect 159294 93922 159362 93978
rect 159418 93922 159486 93978
rect 159542 93922 189834 93978
rect 189890 93922 189958 93978
rect 190014 93922 190082 93978
rect 190138 93922 190206 93978
rect 190262 93922 220554 93978
rect 220610 93922 220678 93978
rect 220734 93922 220802 93978
rect 220858 93922 220926 93978
rect 220982 93922 251274 93978
rect 251330 93922 251398 93978
rect 251454 93922 251522 93978
rect 251578 93922 251646 93978
rect 251702 93922 281994 93978
rect 282050 93922 282118 93978
rect 282174 93922 282242 93978
rect 282298 93922 282366 93978
rect 282422 93922 312714 93978
rect 312770 93922 312838 93978
rect 312894 93922 312962 93978
rect 313018 93922 313086 93978
rect 313142 93922 343434 93978
rect 343490 93922 343558 93978
rect 343614 93922 343682 93978
rect 343738 93922 343806 93978
rect 343862 93922 374154 93978
rect 374210 93922 374278 93978
rect 374334 93922 374402 93978
rect 374458 93922 374526 93978
rect 374582 93922 404874 93978
rect 404930 93922 404998 93978
rect 405054 93922 405122 93978
rect 405178 93922 405246 93978
rect 405302 93922 435594 93978
rect 435650 93922 435718 93978
rect 435774 93922 435842 93978
rect 435898 93922 435966 93978
rect 436022 93922 466314 93978
rect 466370 93922 466438 93978
rect 466494 93922 466562 93978
rect 466618 93922 466686 93978
rect 466742 93922 497034 93978
rect 497090 93922 497158 93978
rect 497214 93922 497282 93978
rect 497338 93922 497406 93978
rect 497462 93922 527754 93978
rect 527810 93922 527878 93978
rect 527934 93922 528002 93978
rect 528058 93922 528126 93978
rect 528182 93922 558474 93978
rect 558530 93922 558598 93978
rect 558654 93922 558722 93978
rect 558778 93922 558846 93978
rect 558902 93922 589194 93978
rect 589250 93922 589318 93978
rect 589374 93922 589442 93978
rect 589498 93922 589566 93978
rect 589622 93922 596496 93978
rect 596552 93922 596620 93978
rect 596676 93922 596744 93978
rect 596800 93922 596868 93978
rect 596924 93922 597980 93978
rect -1916 93826 597980 93922
rect -1916 82350 597980 82446
rect -1916 82294 -1820 82350
rect -1764 82294 -1696 82350
rect -1640 82294 -1572 82350
rect -1516 82294 -1448 82350
rect -1392 82294 9234 82350
rect 9290 82294 9358 82350
rect 9414 82294 9482 82350
rect 9538 82294 9606 82350
rect 9662 82294 39954 82350
rect 40010 82294 40078 82350
rect 40134 82294 40202 82350
rect 40258 82294 40326 82350
rect 40382 82294 70674 82350
rect 70730 82294 70798 82350
rect 70854 82294 70922 82350
rect 70978 82294 71046 82350
rect 71102 82294 101394 82350
rect 101450 82294 101518 82350
rect 101574 82294 101642 82350
rect 101698 82294 101766 82350
rect 101822 82294 132114 82350
rect 132170 82294 132238 82350
rect 132294 82294 132362 82350
rect 132418 82294 132486 82350
rect 132542 82294 162834 82350
rect 162890 82294 162958 82350
rect 163014 82294 163082 82350
rect 163138 82294 163206 82350
rect 163262 82294 193554 82350
rect 193610 82294 193678 82350
rect 193734 82294 193802 82350
rect 193858 82294 193926 82350
rect 193982 82294 224274 82350
rect 224330 82294 224398 82350
rect 224454 82294 224522 82350
rect 224578 82294 224646 82350
rect 224702 82294 254994 82350
rect 255050 82294 255118 82350
rect 255174 82294 255242 82350
rect 255298 82294 255366 82350
rect 255422 82294 285714 82350
rect 285770 82294 285838 82350
rect 285894 82294 285962 82350
rect 286018 82294 286086 82350
rect 286142 82294 316434 82350
rect 316490 82294 316558 82350
rect 316614 82294 316682 82350
rect 316738 82294 316806 82350
rect 316862 82294 347154 82350
rect 347210 82294 347278 82350
rect 347334 82294 347402 82350
rect 347458 82294 347526 82350
rect 347582 82294 377874 82350
rect 377930 82294 377998 82350
rect 378054 82294 378122 82350
rect 378178 82294 378246 82350
rect 378302 82294 408594 82350
rect 408650 82294 408718 82350
rect 408774 82294 408842 82350
rect 408898 82294 408966 82350
rect 409022 82294 439314 82350
rect 439370 82294 439438 82350
rect 439494 82294 439562 82350
rect 439618 82294 439686 82350
rect 439742 82294 470034 82350
rect 470090 82294 470158 82350
rect 470214 82294 470282 82350
rect 470338 82294 470406 82350
rect 470462 82294 500754 82350
rect 500810 82294 500878 82350
rect 500934 82294 501002 82350
rect 501058 82294 501126 82350
rect 501182 82294 531474 82350
rect 531530 82294 531598 82350
rect 531654 82294 531722 82350
rect 531778 82294 531846 82350
rect 531902 82294 562194 82350
rect 562250 82294 562318 82350
rect 562374 82294 562442 82350
rect 562498 82294 562566 82350
rect 562622 82294 592914 82350
rect 592970 82294 593038 82350
rect 593094 82294 593162 82350
rect 593218 82294 593286 82350
rect 593342 82294 597456 82350
rect 597512 82294 597580 82350
rect 597636 82294 597704 82350
rect 597760 82294 597828 82350
rect 597884 82294 597980 82350
rect -1916 82226 597980 82294
rect -1916 82170 -1820 82226
rect -1764 82170 -1696 82226
rect -1640 82170 -1572 82226
rect -1516 82170 -1448 82226
rect -1392 82170 9234 82226
rect 9290 82170 9358 82226
rect 9414 82170 9482 82226
rect 9538 82170 9606 82226
rect 9662 82170 39954 82226
rect 40010 82170 40078 82226
rect 40134 82170 40202 82226
rect 40258 82170 40326 82226
rect 40382 82170 70674 82226
rect 70730 82170 70798 82226
rect 70854 82170 70922 82226
rect 70978 82170 71046 82226
rect 71102 82170 101394 82226
rect 101450 82170 101518 82226
rect 101574 82170 101642 82226
rect 101698 82170 101766 82226
rect 101822 82170 132114 82226
rect 132170 82170 132238 82226
rect 132294 82170 132362 82226
rect 132418 82170 132486 82226
rect 132542 82170 162834 82226
rect 162890 82170 162958 82226
rect 163014 82170 163082 82226
rect 163138 82170 163206 82226
rect 163262 82170 193554 82226
rect 193610 82170 193678 82226
rect 193734 82170 193802 82226
rect 193858 82170 193926 82226
rect 193982 82170 224274 82226
rect 224330 82170 224398 82226
rect 224454 82170 224522 82226
rect 224578 82170 224646 82226
rect 224702 82170 254994 82226
rect 255050 82170 255118 82226
rect 255174 82170 255242 82226
rect 255298 82170 255366 82226
rect 255422 82170 285714 82226
rect 285770 82170 285838 82226
rect 285894 82170 285962 82226
rect 286018 82170 286086 82226
rect 286142 82170 316434 82226
rect 316490 82170 316558 82226
rect 316614 82170 316682 82226
rect 316738 82170 316806 82226
rect 316862 82170 347154 82226
rect 347210 82170 347278 82226
rect 347334 82170 347402 82226
rect 347458 82170 347526 82226
rect 347582 82170 377874 82226
rect 377930 82170 377998 82226
rect 378054 82170 378122 82226
rect 378178 82170 378246 82226
rect 378302 82170 408594 82226
rect 408650 82170 408718 82226
rect 408774 82170 408842 82226
rect 408898 82170 408966 82226
rect 409022 82170 439314 82226
rect 439370 82170 439438 82226
rect 439494 82170 439562 82226
rect 439618 82170 439686 82226
rect 439742 82170 470034 82226
rect 470090 82170 470158 82226
rect 470214 82170 470282 82226
rect 470338 82170 470406 82226
rect 470462 82170 500754 82226
rect 500810 82170 500878 82226
rect 500934 82170 501002 82226
rect 501058 82170 501126 82226
rect 501182 82170 531474 82226
rect 531530 82170 531598 82226
rect 531654 82170 531722 82226
rect 531778 82170 531846 82226
rect 531902 82170 562194 82226
rect 562250 82170 562318 82226
rect 562374 82170 562442 82226
rect 562498 82170 562566 82226
rect 562622 82170 592914 82226
rect 592970 82170 593038 82226
rect 593094 82170 593162 82226
rect 593218 82170 593286 82226
rect 593342 82170 597456 82226
rect 597512 82170 597580 82226
rect 597636 82170 597704 82226
rect 597760 82170 597828 82226
rect 597884 82170 597980 82226
rect -1916 82102 597980 82170
rect -1916 82046 -1820 82102
rect -1764 82046 -1696 82102
rect -1640 82046 -1572 82102
rect -1516 82046 -1448 82102
rect -1392 82046 9234 82102
rect 9290 82046 9358 82102
rect 9414 82046 9482 82102
rect 9538 82046 9606 82102
rect 9662 82046 39954 82102
rect 40010 82046 40078 82102
rect 40134 82046 40202 82102
rect 40258 82046 40326 82102
rect 40382 82046 70674 82102
rect 70730 82046 70798 82102
rect 70854 82046 70922 82102
rect 70978 82046 71046 82102
rect 71102 82046 101394 82102
rect 101450 82046 101518 82102
rect 101574 82046 101642 82102
rect 101698 82046 101766 82102
rect 101822 82046 132114 82102
rect 132170 82046 132238 82102
rect 132294 82046 132362 82102
rect 132418 82046 132486 82102
rect 132542 82046 162834 82102
rect 162890 82046 162958 82102
rect 163014 82046 163082 82102
rect 163138 82046 163206 82102
rect 163262 82046 193554 82102
rect 193610 82046 193678 82102
rect 193734 82046 193802 82102
rect 193858 82046 193926 82102
rect 193982 82046 224274 82102
rect 224330 82046 224398 82102
rect 224454 82046 224522 82102
rect 224578 82046 224646 82102
rect 224702 82046 254994 82102
rect 255050 82046 255118 82102
rect 255174 82046 255242 82102
rect 255298 82046 255366 82102
rect 255422 82046 285714 82102
rect 285770 82046 285838 82102
rect 285894 82046 285962 82102
rect 286018 82046 286086 82102
rect 286142 82046 316434 82102
rect 316490 82046 316558 82102
rect 316614 82046 316682 82102
rect 316738 82046 316806 82102
rect 316862 82046 347154 82102
rect 347210 82046 347278 82102
rect 347334 82046 347402 82102
rect 347458 82046 347526 82102
rect 347582 82046 377874 82102
rect 377930 82046 377998 82102
rect 378054 82046 378122 82102
rect 378178 82046 378246 82102
rect 378302 82046 408594 82102
rect 408650 82046 408718 82102
rect 408774 82046 408842 82102
rect 408898 82046 408966 82102
rect 409022 82046 439314 82102
rect 439370 82046 439438 82102
rect 439494 82046 439562 82102
rect 439618 82046 439686 82102
rect 439742 82046 470034 82102
rect 470090 82046 470158 82102
rect 470214 82046 470282 82102
rect 470338 82046 470406 82102
rect 470462 82046 500754 82102
rect 500810 82046 500878 82102
rect 500934 82046 501002 82102
rect 501058 82046 501126 82102
rect 501182 82046 531474 82102
rect 531530 82046 531598 82102
rect 531654 82046 531722 82102
rect 531778 82046 531846 82102
rect 531902 82046 562194 82102
rect 562250 82046 562318 82102
rect 562374 82046 562442 82102
rect 562498 82046 562566 82102
rect 562622 82046 592914 82102
rect 592970 82046 593038 82102
rect 593094 82046 593162 82102
rect 593218 82046 593286 82102
rect 593342 82046 597456 82102
rect 597512 82046 597580 82102
rect 597636 82046 597704 82102
rect 597760 82046 597828 82102
rect 597884 82046 597980 82102
rect -1916 81978 597980 82046
rect -1916 81922 -1820 81978
rect -1764 81922 -1696 81978
rect -1640 81922 -1572 81978
rect -1516 81922 -1448 81978
rect -1392 81922 9234 81978
rect 9290 81922 9358 81978
rect 9414 81922 9482 81978
rect 9538 81922 9606 81978
rect 9662 81922 39954 81978
rect 40010 81922 40078 81978
rect 40134 81922 40202 81978
rect 40258 81922 40326 81978
rect 40382 81922 70674 81978
rect 70730 81922 70798 81978
rect 70854 81922 70922 81978
rect 70978 81922 71046 81978
rect 71102 81922 101394 81978
rect 101450 81922 101518 81978
rect 101574 81922 101642 81978
rect 101698 81922 101766 81978
rect 101822 81922 132114 81978
rect 132170 81922 132238 81978
rect 132294 81922 132362 81978
rect 132418 81922 132486 81978
rect 132542 81922 162834 81978
rect 162890 81922 162958 81978
rect 163014 81922 163082 81978
rect 163138 81922 163206 81978
rect 163262 81922 193554 81978
rect 193610 81922 193678 81978
rect 193734 81922 193802 81978
rect 193858 81922 193926 81978
rect 193982 81922 224274 81978
rect 224330 81922 224398 81978
rect 224454 81922 224522 81978
rect 224578 81922 224646 81978
rect 224702 81922 254994 81978
rect 255050 81922 255118 81978
rect 255174 81922 255242 81978
rect 255298 81922 255366 81978
rect 255422 81922 285714 81978
rect 285770 81922 285838 81978
rect 285894 81922 285962 81978
rect 286018 81922 286086 81978
rect 286142 81922 316434 81978
rect 316490 81922 316558 81978
rect 316614 81922 316682 81978
rect 316738 81922 316806 81978
rect 316862 81922 347154 81978
rect 347210 81922 347278 81978
rect 347334 81922 347402 81978
rect 347458 81922 347526 81978
rect 347582 81922 377874 81978
rect 377930 81922 377998 81978
rect 378054 81922 378122 81978
rect 378178 81922 378246 81978
rect 378302 81922 408594 81978
rect 408650 81922 408718 81978
rect 408774 81922 408842 81978
rect 408898 81922 408966 81978
rect 409022 81922 439314 81978
rect 439370 81922 439438 81978
rect 439494 81922 439562 81978
rect 439618 81922 439686 81978
rect 439742 81922 470034 81978
rect 470090 81922 470158 81978
rect 470214 81922 470282 81978
rect 470338 81922 470406 81978
rect 470462 81922 500754 81978
rect 500810 81922 500878 81978
rect 500934 81922 501002 81978
rect 501058 81922 501126 81978
rect 501182 81922 531474 81978
rect 531530 81922 531598 81978
rect 531654 81922 531722 81978
rect 531778 81922 531846 81978
rect 531902 81922 562194 81978
rect 562250 81922 562318 81978
rect 562374 81922 562442 81978
rect 562498 81922 562566 81978
rect 562622 81922 592914 81978
rect 592970 81922 593038 81978
rect 593094 81922 593162 81978
rect 593218 81922 593286 81978
rect 593342 81922 597456 81978
rect 597512 81922 597580 81978
rect 597636 81922 597704 81978
rect 597760 81922 597828 81978
rect 597884 81922 597980 81978
rect -1916 81826 597980 81922
rect 3036 80038 99220 80054
rect 3036 79982 3052 80038
rect 3108 79982 99148 80038
rect 99204 79982 99220 80038
rect 3036 79966 99220 79982
rect 6508 79858 341140 79874
rect 6508 79802 6524 79858
rect 6580 79802 341068 79858
rect 341124 79802 341140 79858
rect 6508 79786 341140 79802
rect 85916 79318 446980 79334
rect 85916 79262 85932 79318
rect 85988 79262 446908 79318
rect 446964 79262 446980 79318
rect 85916 79246 446980 79262
rect 89724 79138 480580 79154
rect 89724 79082 89740 79138
rect 89796 79082 480508 79138
rect 480564 79082 480580 79138
rect 89724 79066 480580 79082
rect 8076 78418 121060 78434
rect 8076 78362 8092 78418
rect 8148 78362 120988 78418
rect 121044 78362 121060 78418
rect 8076 78346 121060 78362
rect 6620 78238 297460 78254
rect 6620 78182 6636 78238
rect 6692 78182 297388 78238
rect 297444 78182 297460 78238
rect 6620 78166 297460 78182
rect 11436 78058 590564 78074
rect 11436 78002 11452 78058
rect 11508 78002 590492 78058
rect 590548 78002 590564 78058
rect 11436 77986 590564 78002
rect 92300 77338 497716 77354
rect 92300 77282 92316 77338
rect 92372 77282 497644 77338
rect 497700 77282 497716 77338
rect 92300 77266 497716 77282
rect -1916 76350 597980 76446
rect -1916 76294 -860 76350
rect -804 76294 -736 76350
rect -680 76294 -612 76350
rect -556 76294 -488 76350
rect -432 76294 5514 76350
rect 5570 76294 5638 76350
rect 5694 76294 5762 76350
rect 5818 76294 5886 76350
rect 5942 76294 36234 76350
rect 36290 76294 36358 76350
rect 36414 76294 36482 76350
rect 36538 76294 36606 76350
rect 36662 76294 66954 76350
rect 67010 76294 67078 76350
rect 67134 76294 67202 76350
rect 67258 76294 67326 76350
rect 67382 76294 97674 76350
rect 97730 76294 97798 76350
rect 97854 76294 97922 76350
rect 97978 76294 98046 76350
rect 98102 76294 128394 76350
rect 128450 76294 128518 76350
rect 128574 76294 128642 76350
rect 128698 76294 128766 76350
rect 128822 76294 159114 76350
rect 159170 76294 159238 76350
rect 159294 76294 159362 76350
rect 159418 76294 159486 76350
rect 159542 76294 189834 76350
rect 189890 76294 189958 76350
rect 190014 76294 190082 76350
rect 190138 76294 190206 76350
rect 190262 76294 220554 76350
rect 220610 76294 220678 76350
rect 220734 76294 220802 76350
rect 220858 76294 220926 76350
rect 220982 76294 251274 76350
rect 251330 76294 251398 76350
rect 251454 76294 251522 76350
rect 251578 76294 251646 76350
rect 251702 76294 281994 76350
rect 282050 76294 282118 76350
rect 282174 76294 282242 76350
rect 282298 76294 282366 76350
rect 282422 76294 312714 76350
rect 312770 76294 312838 76350
rect 312894 76294 312962 76350
rect 313018 76294 313086 76350
rect 313142 76294 343434 76350
rect 343490 76294 343558 76350
rect 343614 76294 343682 76350
rect 343738 76294 343806 76350
rect 343862 76294 374154 76350
rect 374210 76294 374278 76350
rect 374334 76294 374402 76350
rect 374458 76294 374526 76350
rect 374582 76294 404874 76350
rect 404930 76294 404998 76350
rect 405054 76294 405122 76350
rect 405178 76294 405246 76350
rect 405302 76294 435594 76350
rect 435650 76294 435718 76350
rect 435774 76294 435842 76350
rect 435898 76294 435966 76350
rect 436022 76294 466314 76350
rect 466370 76294 466438 76350
rect 466494 76294 466562 76350
rect 466618 76294 466686 76350
rect 466742 76294 497034 76350
rect 497090 76294 497158 76350
rect 497214 76294 497282 76350
rect 497338 76294 497406 76350
rect 497462 76294 527754 76350
rect 527810 76294 527878 76350
rect 527934 76294 528002 76350
rect 528058 76294 528126 76350
rect 528182 76294 558474 76350
rect 558530 76294 558598 76350
rect 558654 76294 558722 76350
rect 558778 76294 558846 76350
rect 558902 76294 589194 76350
rect 589250 76294 589318 76350
rect 589374 76294 589442 76350
rect 589498 76294 589566 76350
rect 589622 76294 596496 76350
rect 596552 76294 596620 76350
rect 596676 76294 596744 76350
rect 596800 76294 596868 76350
rect 596924 76294 597980 76350
rect -1916 76226 597980 76294
rect -1916 76170 -860 76226
rect -804 76170 -736 76226
rect -680 76170 -612 76226
rect -556 76170 -488 76226
rect -432 76170 5514 76226
rect 5570 76170 5638 76226
rect 5694 76170 5762 76226
rect 5818 76170 5886 76226
rect 5942 76170 36234 76226
rect 36290 76170 36358 76226
rect 36414 76170 36482 76226
rect 36538 76170 36606 76226
rect 36662 76170 66954 76226
rect 67010 76170 67078 76226
rect 67134 76170 67202 76226
rect 67258 76170 67326 76226
rect 67382 76170 97674 76226
rect 97730 76170 97798 76226
rect 97854 76170 97922 76226
rect 97978 76170 98046 76226
rect 98102 76170 128394 76226
rect 128450 76170 128518 76226
rect 128574 76170 128642 76226
rect 128698 76170 128766 76226
rect 128822 76170 159114 76226
rect 159170 76170 159238 76226
rect 159294 76170 159362 76226
rect 159418 76170 159486 76226
rect 159542 76170 189834 76226
rect 189890 76170 189958 76226
rect 190014 76170 190082 76226
rect 190138 76170 190206 76226
rect 190262 76170 220554 76226
rect 220610 76170 220678 76226
rect 220734 76170 220802 76226
rect 220858 76170 220926 76226
rect 220982 76170 251274 76226
rect 251330 76170 251398 76226
rect 251454 76170 251522 76226
rect 251578 76170 251646 76226
rect 251702 76170 281994 76226
rect 282050 76170 282118 76226
rect 282174 76170 282242 76226
rect 282298 76170 282366 76226
rect 282422 76170 312714 76226
rect 312770 76170 312838 76226
rect 312894 76170 312962 76226
rect 313018 76170 313086 76226
rect 313142 76170 343434 76226
rect 343490 76170 343558 76226
rect 343614 76170 343682 76226
rect 343738 76170 343806 76226
rect 343862 76170 374154 76226
rect 374210 76170 374278 76226
rect 374334 76170 374402 76226
rect 374458 76170 374526 76226
rect 374582 76170 404874 76226
rect 404930 76170 404998 76226
rect 405054 76170 405122 76226
rect 405178 76170 405246 76226
rect 405302 76170 435594 76226
rect 435650 76170 435718 76226
rect 435774 76170 435842 76226
rect 435898 76170 435966 76226
rect 436022 76170 466314 76226
rect 466370 76170 466438 76226
rect 466494 76170 466562 76226
rect 466618 76170 466686 76226
rect 466742 76170 497034 76226
rect 497090 76170 497158 76226
rect 497214 76170 497282 76226
rect 497338 76170 497406 76226
rect 497462 76170 527754 76226
rect 527810 76170 527878 76226
rect 527934 76170 528002 76226
rect 528058 76170 528126 76226
rect 528182 76170 558474 76226
rect 558530 76170 558598 76226
rect 558654 76170 558722 76226
rect 558778 76170 558846 76226
rect 558902 76170 589194 76226
rect 589250 76170 589318 76226
rect 589374 76170 589442 76226
rect 589498 76170 589566 76226
rect 589622 76170 596496 76226
rect 596552 76170 596620 76226
rect 596676 76170 596744 76226
rect 596800 76170 596868 76226
rect 596924 76170 597980 76226
rect -1916 76102 597980 76170
rect -1916 76046 -860 76102
rect -804 76046 -736 76102
rect -680 76046 -612 76102
rect -556 76046 -488 76102
rect -432 76046 5514 76102
rect 5570 76046 5638 76102
rect 5694 76046 5762 76102
rect 5818 76046 5886 76102
rect 5942 76046 36234 76102
rect 36290 76046 36358 76102
rect 36414 76046 36482 76102
rect 36538 76046 36606 76102
rect 36662 76046 66954 76102
rect 67010 76046 67078 76102
rect 67134 76046 67202 76102
rect 67258 76046 67326 76102
rect 67382 76046 97674 76102
rect 97730 76046 97798 76102
rect 97854 76046 97922 76102
rect 97978 76046 98046 76102
rect 98102 76046 128394 76102
rect 128450 76046 128518 76102
rect 128574 76046 128642 76102
rect 128698 76046 128766 76102
rect 128822 76046 159114 76102
rect 159170 76046 159238 76102
rect 159294 76046 159362 76102
rect 159418 76046 159486 76102
rect 159542 76046 189834 76102
rect 189890 76046 189958 76102
rect 190014 76046 190082 76102
rect 190138 76046 190206 76102
rect 190262 76046 220554 76102
rect 220610 76046 220678 76102
rect 220734 76046 220802 76102
rect 220858 76046 220926 76102
rect 220982 76046 251274 76102
rect 251330 76046 251398 76102
rect 251454 76046 251522 76102
rect 251578 76046 251646 76102
rect 251702 76046 281994 76102
rect 282050 76046 282118 76102
rect 282174 76046 282242 76102
rect 282298 76046 282366 76102
rect 282422 76046 312714 76102
rect 312770 76046 312838 76102
rect 312894 76046 312962 76102
rect 313018 76046 313086 76102
rect 313142 76046 343434 76102
rect 343490 76046 343558 76102
rect 343614 76046 343682 76102
rect 343738 76046 343806 76102
rect 343862 76046 374154 76102
rect 374210 76046 374278 76102
rect 374334 76046 374402 76102
rect 374458 76046 374526 76102
rect 374582 76046 404874 76102
rect 404930 76046 404998 76102
rect 405054 76046 405122 76102
rect 405178 76046 405246 76102
rect 405302 76046 435594 76102
rect 435650 76046 435718 76102
rect 435774 76046 435842 76102
rect 435898 76046 435966 76102
rect 436022 76046 466314 76102
rect 466370 76046 466438 76102
rect 466494 76046 466562 76102
rect 466618 76046 466686 76102
rect 466742 76046 497034 76102
rect 497090 76046 497158 76102
rect 497214 76046 497282 76102
rect 497338 76046 497406 76102
rect 497462 76046 527754 76102
rect 527810 76046 527878 76102
rect 527934 76046 528002 76102
rect 528058 76046 528126 76102
rect 528182 76046 558474 76102
rect 558530 76046 558598 76102
rect 558654 76046 558722 76102
rect 558778 76046 558846 76102
rect 558902 76046 589194 76102
rect 589250 76046 589318 76102
rect 589374 76046 589442 76102
rect 589498 76046 589566 76102
rect 589622 76046 596496 76102
rect 596552 76046 596620 76102
rect 596676 76046 596744 76102
rect 596800 76046 596868 76102
rect 596924 76046 597980 76102
rect -1916 75978 597980 76046
rect -1916 75922 -860 75978
rect -804 75922 -736 75978
rect -680 75922 -612 75978
rect -556 75922 -488 75978
rect -432 75922 5514 75978
rect 5570 75922 5638 75978
rect 5694 75922 5762 75978
rect 5818 75922 5886 75978
rect 5942 75922 36234 75978
rect 36290 75922 36358 75978
rect 36414 75922 36482 75978
rect 36538 75922 36606 75978
rect 36662 75922 66954 75978
rect 67010 75922 67078 75978
rect 67134 75922 67202 75978
rect 67258 75922 67326 75978
rect 67382 75922 97674 75978
rect 97730 75922 97798 75978
rect 97854 75922 97922 75978
rect 97978 75922 98046 75978
rect 98102 75922 128394 75978
rect 128450 75922 128518 75978
rect 128574 75922 128642 75978
rect 128698 75922 128766 75978
rect 128822 75922 159114 75978
rect 159170 75922 159238 75978
rect 159294 75922 159362 75978
rect 159418 75922 159486 75978
rect 159542 75922 189834 75978
rect 189890 75922 189958 75978
rect 190014 75922 190082 75978
rect 190138 75922 190206 75978
rect 190262 75922 220554 75978
rect 220610 75922 220678 75978
rect 220734 75922 220802 75978
rect 220858 75922 220926 75978
rect 220982 75922 251274 75978
rect 251330 75922 251398 75978
rect 251454 75922 251522 75978
rect 251578 75922 251646 75978
rect 251702 75922 281994 75978
rect 282050 75922 282118 75978
rect 282174 75922 282242 75978
rect 282298 75922 282366 75978
rect 282422 75922 312714 75978
rect 312770 75922 312838 75978
rect 312894 75922 312962 75978
rect 313018 75922 313086 75978
rect 313142 75922 343434 75978
rect 343490 75922 343558 75978
rect 343614 75922 343682 75978
rect 343738 75922 343806 75978
rect 343862 75922 374154 75978
rect 374210 75922 374278 75978
rect 374334 75922 374402 75978
rect 374458 75922 374526 75978
rect 374582 75922 404874 75978
rect 404930 75922 404998 75978
rect 405054 75922 405122 75978
rect 405178 75922 405246 75978
rect 405302 75922 435594 75978
rect 435650 75922 435718 75978
rect 435774 75922 435842 75978
rect 435898 75922 435966 75978
rect 436022 75922 466314 75978
rect 466370 75922 466438 75978
rect 466494 75922 466562 75978
rect 466618 75922 466686 75978
rect 466742 75922 497034 75978
rect 497090 75922 497158 75978
rect 497214 75922 497282 75978
rect 497338 75922 497406 75978
rect 497462 75922 527754 75978
rect 527810 75922 527878 75978
rect 527934 75922 528002 75978
rect 528058 75922 528126 75978
rect 528182 75922 558474 75978
rect 558530 75922 558598 75978
rect 558654 75922 558722 75978
rect 558778 75922 558846 75978
rect 558902 75922 589194 75978
rect 589250 75922 589318 75978
rect 589374 75922 589442 75978
rect 589498 75922 589566 75978
rect 589622 75922 596496 75978
rect 596552 75922 596620 75978
rect 596676 75922 596744 75978
rect 596800 75922 596868 75978
rect 596924 75922 597980 75978
rect -1916 75826 597980 75922
rect 7964 74998 164740 75014
rect 7964 74942 7980 74998
rect 8036 74942 164668 74998
rect 164724 74942 164740 74998
rect 7964 74926 164740 74942
rect 11548 74818 186580 74834
rect 11548 74762 11564 74818
rect 11620 74762 186508 74818
rect 186564 74762 186580 74818
rect 11548 74746 186580 74762
rect 99916 74278 123860 74294
rect 99916 74222 99932 74278
rect 99988 74222 123788 74278
rect 123844 74222 123860 74278
rect 99916 74206 123860 74222
rect 87260 74098 452020 74114
rect 87260 74042 87276 74098
rect 87332 74042 451948 74098
rect 452004 74042 452020 74098
rect 87260 74026 452020 74042
rect 80092 72658 383140 72674
rect 80092 72602 80108 72658
rect 80164 72602 383068 72658
rect 383124 72602 383140 72658
rect 80092 72586 383140 72602
rect 84572 72478 435220 72494
rect 84572 72422 84588 72478
rect 84644 72422 435148 72478
rect 435204 72422 435220 72478
rect 84572 72406 435220 72422
rect 88940 72298 468820 72314
rect 88940 72242 88956 72298
rect 89012 72242 468748 72298
rect 468804 72242 468820 72298
rect 88940 72226 468820 72242
rect 8972 72118 15220 72134
rect 8972 72062 8988 72118
rect 9044 72062 15148 72118
rect 15204 72062 15220 72118
rect 8972 72046 15220 72062
rect 94876 71398 206740 71414
rect 94876 71342 94892 71398
rect 94948 71342 206668 71398
rect 206724 71342 206740 71398
rect 94876 71326 206740 71342
rect 89836 71218 248740 71234
rect 89836 71162 89852 71218
rect 89908 71162 248668 71218
rect 248724 71162 248740 71218
rect 89836 71146 248740 71162
rect 88268 71038 263860 71054
rect 88268 70982 88284 71038
rect 88340 70982 263788 71038
rect 263844 70982 263860 71038
rect 88268 70966 263860 70982
rect 68668 70858 289060 70874
rect 68668 70802 68684 70858
rect 68740 70802 288988 70858
rect 289044 70802 289060 70858
rect 68668 70786 289060 70802
rect 65196 70678 295780 70694
rect 65196 70622 65212 70678
rect 65268 70622 295708 70678
rect 295764 70622 295780 70678
rect 65196 70606 295780 70622
rect 56124 69418 238660 69434
rect 56124 69362 56140 69418
rect 56196 69362 238588 69418
rect 238644 69362 238660 69418
rect 56124 69346 238660 69362
rect 83116 69238 286372 69254
rect 83116 69182 83132 69238
rect 83188 69182 286300 69238
rect 286356 69182 286372 69238
rect 83116 69166 286372 69182
rect 12668 69058 16004 69074
rect 12668 69002 12684 69058
rect 12740 69002 15932 69058
rect 15988 69002 16004 69058
rect 12668 68986 16004 69002
rect 70124 69058 302500 69074
rect 70124 69002 70140 69058
rect 70196 69002 302428 69058
rect 302484 69002 302500 69058
rect 70124 68986 302500 69002
rect 8860 68878 13540 68894
rect 8860 68822 8876 68878
rect 8932 68822 13468 68878
rect 13524 68822 13540 68878
rect 8860 68806 13540 68822
rect 91628 67978 223540 67994
rect 91628 67922 91644 67978
rect 91700 67922 223468 67978
rect 223524 67922 223540 67978
rect 91628 67906 223540 67922
rect 83340 67798 305860 67814
rect 83340 67742 83356 67798
rect 83412 67742 305788 67798
rect 305844 67742 305860 67798
rect 83340 67726 305860 67742
rect 66540 67618 294100 67634
rect 66540 67562 66556 67618
rect 66612 67562 294028 67618
rect 294084 67562 294100 67618
rect 66540 67546 294100 67562
rect 84124 67438 431860 67454
rect 84124 67382 84140 67438
rect 84196 67382 431788 67438
rect 431844 67382 431860 67438
rect 84124 67366 431860 67382
rect 100588 67258 572980 67274
rect 100588 67202 100604 67258
rect 100660 67202 572908 67258
rect 572964 67202 572980 67258
rect 100588 67186 572980 67202
rect 12668 67078 29444 67094
rect 12668 67022 12684 67078
rect 12740 67022 29372 67078
rect 29428 67022 29444 67078
rect 12668 67006 29444 67022
rect 91740 66358 235300 66374
rect 91740 66302 91756 66358
rect 91812 66302 235228 66358
rect 235284 66302 235300 66358
rect 91740 66286 235300 66302
rect 87372 66178 258820 66194
rect 87372 66122 87388 66178
rect 87444 66122 258748 66178
rect 258804 66122 258820 66178
rect 87372 66106 258820 66122
rect 84908 65998 317620 66014
rect 84908 65942 84924 65998
rect 84980 65942 317548 65998
rect 317604 65942 317620 65998
rect 84908 65926 317620 65942
rect 81212 65818 406660 65834
rect 81212 65762 81228 65818
rect 81284 65762 406588 65818
rect 406644 65762 406660 65818
rect 81212 65746 406660 65762
rect 102044 65638 576340 65654
rect 102044 65582 102060 65638
rect 102116 65582 576268 65638
rect 576324 65582 576340 65638
rect 102044 65566 576340 65582
rect 12444 65458 76484 65474
rect 12444 65402 12460 65458
rect 12516 65402 76412 65458
rect 76468 65402 76484 65458
rect 12444 65386 76484 65402
rect 84684 64918 252100 64934
rect 84684 64862 84700 64918
rect 84756 64862 252028 64918
rect 252084 64862 252100 64918
rect 84684 64846 252100 64862
rect 78412 64738 253780 64754
rect 78412 64682 78428 64738
rect 78484 64682 253708 64738
rect 253764 64682 253780 64738
rect 78412 64666 253780 64682
rect -1916 64350 597980 64446
rect -1916 64294 -1820 64350
rect -1764 64294 -1696 64350
rect -1640 64294 -1572 64350
rect -1516 64294 -1448 64350
rect -1392 64294 9234 64350
rect 9290 64294 9358 64350
rect 9414 64294 9482 64350
rect 9538 64294 9606 64350
rect 9662 64294 31878 64350
rect 31934 64294 32002 64350
rect 32058 64294 39954 64350
rect 40010 64294 40078 64350
rect 40134 64294 40202 64350
rect 40258 64294 40326 64350
rect 40382 64294 62598 64350
rect 62654 64294 62722 64350
rect 62778 64294 70674 64350
rect 70730 64294 70798 64350
rect 70854 64294 70922 64350
rect 70978 64294 71046 64350
rect 71102 64294 93318 64350
rect 93374 64294 93442 64350
rect 93498 64294 101394 64350
rect 101450 64294 101518 64350
rect 101574 64294 101642 64350
rect 101698 64294 101766 64350
rect 101822 64294 132114 64350
rect 132170 64294 132238 64350
rect 132294 64294 132362 64350
rect 132418 64294 132486 64350
rect 132542 64294 162834 64350
rect 162890 64294 162958 64350
rect 163014 64294 163082 64350
rect 163138 64294 163206 64350
rect 163262 64294 193554 64350
rect 193610 64294 193678 64350
rect 193734 64294 193802 64350
rect 193858 64294 193926 64350
rect 193982 64294 224274 64350
rect 224330 64294 224398 64350
rect 224454 64294 224522 64350
rect 224578 64294 224646 64350
rect 224702 64294 254994 64350
rect 255050 64294 255118 64350
rect 255174 64294 255242 64350
rect 255298 64294 255366 64350
rect 255422 64294 285714 64350
rect 285770 64294 285838 64350
rect 285894 64294 285962 64350
rect 286018 64294 286086 64350
rect 286142 64294 316434 64350
rect 316490 64294 316558 64350
rect 316614 64294 316682 64350
rect 316738 64294 316806 64350
rect 316862 64294 347154 64350
rect 347210 64294 347278 64350
rect 347334 64294 347402 64350
rect 347458 64294 347526 64350
rect 347582 64294 377874 64350
rect 377930 64294 377998 64350
rect 378054 64294 378122 64350
rect 378178 64294 378246 64350
rect 378302 64294 408594 64350
rect 408650 64294 408718 64350
rect 408774 64294 408842 64350
rect 408898 64294 408966 64350
rect 409022 64294 439314 64350
rect 439370 64294 439438 64350
rect 439494 64294 439562 64350
rect 439618 64294 439686 64350
rect 439742 64294 470034 64350
rect 470090 64294 470158 64350
rect 470214 64294 470282 64350
rect 470338 64294 470406 64350
rect 470462 64294 500754 64350
rect 500810 64294 500878 64350
rect 500934 64294 501002 64350
rect 501058 64294 501126 64350
rect 501182 64294 531474 64350
rect 531530 64294 531598 64350
rect 531654 64294 531722 64350
rect 531778 64294 531846 64350
rect 531902 64294 562194 64350
rect 562250 64294 562318 64350
rect 562374 64294 562442 64350
rect 562498 64294 562566 64350
rect 562622 64294 592914 64350
rect 592970 64294 593038 64350
rect 593094 64294 593162 64350
rect 593218 64294 593286 64350
rect 593342 64294 597456 64350
rect 597512 64294 597580 64350
rect 597636 64294 597704 64350
rect 597760 64294 597828 64350
rect 597884 64294 597980 64350
rect -1916 64226 597980 64294
rect -1916 64170 -1820 64226
rect -1764 64170 -1696 64226
rect -1640 64170 -1572 64226
rect -1516 64170 -1448 64226
rect -1392 64170 9234 64226
rect 9290 64170 9358 64226
rect 9414 64170 9482 64226
rect 9538 64170 9606 64226
rect 9662 64170 31878 64226
rect 31934 64170 32002 64226
rect 32058 64170 39954 64226
rect 40010 64170 40078 64226
rect 40134 64170 40202 64226
rect 40258 64170 40326 64226
rect 40382 64170 62598 64226
rect 62654 64170 62722 64226
rect 62778 64170 70674 64226
rect 70730 64170 70798 64226
rect 70854 64170 70922 64226
rect 70978 64170 71046 64226
rect 71102 64170 93318 64226
rect 93374 64170 93442 64226
rect 93498 64170 101394 64226
rect 101450 64170 101518 64226
rect 101574 64170 101642 64226
rect 101698 64170 101766 64226
rect 101822 64170 132114 64226
rect 132170 64170 132238 64226
rect 132294 64170 132362 64226
rect 132418 64170 132486 64226
rect 132542 64170 162834 64226
rect 162890 64170 162958 64226
rect 163014 64170 163082 64226
rect 163138 64170 163206 64226
rect 163262 64170 193554 64226
rect 193610 64170 193678 64226
rect 193734 64170 193802 64226
rect 193858 64170 193926 64226
rect 193982 64170 224274 64226
rect 224330 64170 224398 64226
rect 224454 64170 224522 64226
rect 224578 64170 224646 64226
rect 224702 64170 254994 64226
rect 255050 64170 255118 64226
rect 255174 64170 255242 64226
rect 255298 64170 255366 64226
rect 255422 64170 285714 64226
rect 285770 64170 285838 64226
rect 285894 64170 285962 64226
rect 286018 64170 286086 64226
rect 286142 64170 316434 64226
rect 316490 64170 316558 64226
rect 316614 64170 316682 64226
rect 316738 64170 316806 64226
rect 316862 64170 347154 64226
rect 347210 64170 347278 64226
rect 347334 64170 347402 64226
rect 347458 64170 347526 64226
rect 347582 64170 377874 64226
rect 377930 64170 377998 64226
rect 378054 64170 378122 64226
rect 378178 64170 378246 64226
rect 378302 64170 408594 64226
rect 408650 64170 408718 64226
rect 408774 64170 408842 64226
rect 408898 64170 408966 64226
rect 409022 64170 439314 64226
rect 439370 64170 439438 64226
rect 439494 64170 439562 64226
rect 439618 64170 439686 64226
rect 439742 64170 470034 64226
rect 470090 64170 470158 64226
rect 470214 64170 470282 64226
rect 470338 64170 470406 64226
rect 470462 64170 500754 64226
rect 500810 64170 500878 64226
rect 500934 64170 501002 64226
rect 501058 64170 501126 64226
rect 501182 64170 531474 64226
rect 531530 64170 531598 64226
rect 531654 64170 531722 64226
rect 531778 64170 531846 64226
rect 531902 64170 562194 64226
rect 562250 64170 562318 64226
rect 562374 64170 562442 64226
rect 562498 64170 562566 64226
rect 562622 64170 592914 64226
rect 592970 64170 593038 64226
rect 593094 64170 593162 64226
rect 593218 64170 593286 64226
rect 593342 64170 597456 64226
rect 597512 64170 597580 64226
rect 597636 64170 597704 64226
rect 597760 64170 597828 64226
rect 597884 64170 597980 64226
rect -1916 64102 597980 64170
rect -1916 64046 -1820 64102
rect -1764 64046 -1696 64102
rect -1640 64046 -1572 64102
rect -1516 64046 -1448 64102
rect -1392 64046 9234 64102
rect 9290 64046 9358 64102
rect 9414 64046 9482 64102
rect 9538 64046 9606 64102
rect 9662 64046 31878 64102
rect 31934 64046 32002 64102
rect 32058 64046 39954 64102
rect 40010 64046 40078 64102
rect 40134 64046 40202 64102
rect 40258 64046 40326 64102
rect 40382 64046 62598 64102
rect 62654 64046 62722 64102
rect 62778 64046 70674 64102
rect 70730 64046 70798 64102
rect 70854 64046 70922 64102
rect 70978 64046 71046 64102
rect 71102 64046 93318 64102
rect 93374 64046 93442 64102
rect 93498 64046 101394 64102
rect 101450 64046 101518 64102
rect 101574 64046 101642 64102
rect 101698 64046 101766 64102
rect 101822 64046 132114 64102
rect 132170 64046 132238 64102
rect 132294 64046 132362 64102
rect 132418 64046 132486 64102
rect 132542 64046 162834 64102
rect 162890 64046 162958 64102
rect 163014 64046 163082 64102
rect 163138 64046 163206 64102
rect 163262 64046 193554 64102
rect 193610 64046 193678 64102
rect 193734 64046 193802 64102
rect 193858 64046 193926 64102
rect 193982 64046 224274 64102
rect 224330 64046 224398 64102
rect 224454 64046 224522 64102
rect 224578 64046 224646 64102
rect 224702 64046 254994 64102
rect 255050 64046 255118 64102
rect 255174 64046 255242 64102
rect 255298 64046 255366 64102
rect 255422 64046 285714 64102
rect 285770 64046 285838 64102
rect 285894 64046 285962 64102
rect 286018 64046 286086 64102
rect 286142 64046 316434 64102
rect 316490 64046 316558 64102
rect 316614 64046 316682 64102
rect 316738 64046 316806 64102
rect 316862 64046 347154 64102
rect 347210 64046 347278 64102
rect 347334 64046 347402 64102
rect 347458 64046 347526 64102
rect 347582 64046 377874 64102
rect 377930 64046 377998 64102
rect 378054 64046 378122 64102
rect 378178 64046 378246 64102
rect 378302 64046 408594 64102
rect 408650 64046 408718 64102
rect 408774 64046 408842 64102
rect 408898 64046 408966 64102
rect 409022 64046 439314 64102
rect 439370 64046 439438 64102
rect 439494 64046 439562 64102
rect 439618 64046 439686 64102
rect 439742 64046 470034 64102
rect 470090 64046 470158 64102
rect 470214 64046 470282 64102
rect 470338 64046 470406 64102
rect 470462 64046 500754 64102
rect 500810 64046 500878 64102
rect 500934 64046 501002 64102
rect 501058 64046 501126 64102
rect 501182 64046 531474 64102
rect 531530 64046 531598 64102
rect 531654 64046 531722 64102
rect 531778 64046 531846 64102
rect 531902 64046 562194 64102
rect 562250 64046 562318 64102
rect 562374 64046 562442 64102
rect 562498 64046 562566 64102
rect 562622 64046 592914 64102
rect 592970 64046 593038 64102
rect 593094 64046 593162 64102
rect 593218 64046 593286 64102
rect 593342 64046 597456 64102
rect 597512 64046 597580 64102
rect 597636 64046 597704 64102
rect 597760 64046 597828 64102
rect 597884 64046 597980 64102
rect -1916 63978 597980 64046
rect -1916 63922 -1820 63978
rect -1764 63922 -1696 63978
rect -1640 63922 -1572 63978
rect -1516 63922 -1448 63978
rect -1392 63922 9234 63978
rect 9290 63922 9358 63978
rect 9414 63922 9482 63978
rect 9538 63922 9606 63978
rect 9662 63922 31878 63978
rect 31934 63922 32002 63978
rect 32058 63922 39954 63978
rect 40010 63922 40078 63978
rect 40134 63922 40202 63978
rect 40258 63922 40326 63978
rect 40382 63922 62598 63978
rect 62654 63922 62722 63978
rect 62778 63922 70674 63978
rect 70730 63922 70798 63978
rect 70854 63922 70922 63978
rect 70978 63922 71046 63978
rect 71102 63922 93318 63978
rect 93374 63922 93442 63978
rect 93498 63922 101394 63978
rect 101450 63922 101518 63978
rect 101574 63922 101642 63978
rect 101698 63922 101766 63978
rect 101822 63922 132114 63978
rect 132170 63922 132238 63978
rect 132294 63922 132362 63978
rect 132418 63922 132486 63978
rect 132542 63922 162834 63978
rect 162890 63922 162958 63978
rect 163014 63922 163082 63978
rect 163138 63922 163206 63978
rect 163262 63922 193554 63978
rect 193610 63922 193678 63978
rect 193734 63922 193802 63978
rect 193858 63922 193926 63978
rect 193982 63922 224274 63978
rect 224330 63922 224398 63978
rect 224454 63922 224522 63978
rect 224578 63922 224646 63978
rect 224702 63922 254994 63978
rect 255050 63922 255118 63978
rect 255174 63922 255242 63978
rect 255298 63922 255366 63978
rect 255422 63922 285714 63978
rect 285770 63922 285838 63978
rect 285894 63922 285962 63978
rect 286018 63922 286086 63978
rect 286142 63922 316434 63978
rect 316490 63922 316558 63978
rect 316614 63922 316682 63978
rect 316738 63922 316806 63978
rect 316862 63922 347154 63978
rect 347210 63922 347278 63978
rect 347334 63922 347402 63978
rect 347458 63922 347526 63978
rect 347582 63922 377874 63978
rect 377930 63922 377998 63978
rect 378054 63922 378122 63978
rect 378178 63922 378246 63978
rect 378302 63922 408594 63978
rect 408650 63922 408718 63978
rect 408774 63922 408842 63978
rect 408898 63922 408966 63978
rect 409022 63922 439314 63978
rect 439370 63922 439438 63978
rect 439494 63922 439562 63978
rect 439618 63922 439686 63978
rect 439742 63922 470034 63978
rect 470090 63922 470158 63978
rect 470214 63922 470282 63978
rect 470338 63922 470406 63978
rect 470462 63922 500754 63978
rect 500810 63922 500878 63978
rect 500934 63922 501002 63978
rect 501058 63922 501126 63978
rect 501182 63922 531474 63978
rect 531530 63922 531598 63978
rect 531654 63922 531722 63978
rect 531778 63922 531846 63978
rect 531902 63922 562194 63978
rect 562250 63922 562318 63978
rect 562374 63922 562442 63978
rect 562498 63922 562566 63978
rect 562622 63922 592914 63978
rect 592970 63922 593038 63978
rect 593094 63922 593162 63978
rect 593218 63922 593286 63978
rect 593342 63922 597456 63978
rect 597512 63922 597580 63978
rect 597636 63922 597704 63978
rect 597760 63922 597828 63978
rect 597884 63922 597980 63978
rect -1916 63826 597980 63922
rect 12444 63658 86564 63674
rect 12444 63602 12460 63658
rect 12516 63602 86492 63658
rect 86548 63602 86564 63658
rect 12444 63586 86564 63602
rect 63180 62938 87460 62954
rect 63180 62882 63196 62938
rect 63252 62882 87388 62938
rect 87444 62882 87460 62938
rect 63180 62866 87460 62882
rect 76396 62578 324340 62594
rect 76396 62522 76412 62578
rect 76468 62522 324268 62578
rect 324324 62522 324340 62578
rect 76396 62506 324340 62522
rect 88828 62398 472180 62414
rect 88828 62342 88844 62398
rect 88900 62342 472108 62398
rect 472164 62342 472180 62398
rect 88828 62326 472180 62342
rect 95660 62218 525940 62234
rect 95660 62162 95676 62218
rect 95732 62162 525868 62218
rect 525924 62162 525940 62218
rect 95660 62146 525940 62162
rect 12668 62038 21044 62054
rect 12668 61982 12684 62038
rect 12740 61982 20972 62038
rect 21028 61982 21044 62038
rect 12668 61966 21044 61982
rect 80540 61318 166420 61334
rect 80540 61262 80556 61318
rect 80612 61262 166348 61318
rect 166404 61262 166420 61318
rect 80540 61246 166420 61262
rect 58700 61138 216820 61154
rect 58700 61082 58716 61138
rect 58772 61082 216748 61138
rect 216804 61082 216820 61138
rect 58700 61066 216820 61082
rect 83228 60958 396580 60974
rect 83228 60902 83244 60958
rect 83300 60902 396508 60958
rect 396564 60902 396580 60958
rect 83228 60886 396580 60902
rect 12668 60778 14324 60794
rect 12668 60722 12684 60778
rect 12740 60722 14252 60778
rect 14308 60722 14324 60778
rect 12668 60706 14324 60722
rect 90620 60778 482260 60794
rect 90620 60722 90636 60778
rect 90692 60722 482188 60778
rect 482244 60722 482260 60778
rect 90620 60706 482260 60722
rect 92860 60598 515860 60614
rect 92860 60542 92876 60598
rect 92932 60542 515788 60598
rect 515844 60542 515860 60598
rect 92860 60526 515860 60542
rect 12444 60418 31124 60434
rect 12444 60362 12460 60418
rect 12516 60362 31052 60418
rect 31108 60362 31124 60418
rect 12444 60346 31124 60362
rect 79868 60418 89924 60434
rect 79868 60362 79884 60418
rect 79940 60362 89852 60418
rect 89908 60362 89924 60418
rect 79868 60346 89924 60362
rect 63628 60058 84772 60074
rect 63628 60002 63644 60058
rect 63700 60002 84700 60058
rect 84756 60002 84772 60058
rect 63628 59986 84772 60002
rect 54556 59878 80628 59894
rect 54556 59822 54572 59878
rect 54628 59822 80556 59878
rect 80612 59822 80628 59878
rect 54556 59806 80628 59822
rect 73148 59698 273940 59714
rect 73148 59642 73164 59698
rect 73220 59642 273868 59698
rect 273924 59642 273940 59698
rect 73148 59626 273940 59642
rect 74828 59518 322660 59534
rect 74828 59462 74844 59518
rect 74900 59462 322588 59518
rect 322644 59462 322660 59518
rect 74828 59446 322660 59462
rect 87148 59338 458740 59354
rect 87148 59282 87164 59338
rect 87220 59282 458668 59338
rect 458724 59282 458740 59338
rect 87148 59266 458740 59282
rect 89500 59158 477220 59174
rect 89500 59102 89516 59158
rect 89572 59102 477148 59158
rect 477204 59102 477220 59158
rect 89500 59086 477220 59102
rect 95548 58978 520900 58994
rect 95548 58922 95564 58978
rect 95620 58922 520828 58978
rect 520884 58922 520900 58978
rect 95548 58906 520900 58922
rect -1916 58350 597980 58446
rect -1916 58294 -860 58350
rect -804 58294 -736 58350
rect -680 58294 -612 58350
rect -556 58294 -488 58350
rect -432 58294 5514 58350
rect 5570 58294 5638 58350
rect 5694 58294 5762 58350
rect 5818 58294 5886 58350
rect 5942 58294 16518 58350
rect 16574 58294 16642 58350
rect 16698 58294 36234 58350
rect 36290 58294 36358 58350
rect 36414 58294 36482 58350
rect 36538 58294 36606 58350
rect 36662 58294 47238 58350
rect 47294 58294 47362 58350
rect 47418 58294 66954 58350
rect 67010 58294 67078 58350
rect 67134 58294 67202 58350
rect 67258 58294 67326 58350
rect 67382 58294 77958 58350
rect 78014 58294 78082 58350
rect 78138 58294 97674 58350
rect 97730 58294 97798 58350
rect 97854 58294 97922 58350
rect 97978 58294 98046 58350
rect 98102 58294 108678 58350
rect 108734 58294 108802 58350
rect 108858 58294 128394 58350
rect 128450 58294 128518 58350
rect 128574 58294 128642 58350
rect 128698 58294 128766 58350
rect 128822 58294 159114 58350
rect 159170 58294 159238 58350
rect 159294 58294 159362 58350
rect 159418 58294 159486 58350
rect 159542 58294 189834 58350
rect 189890 58294 189958 58350
rect 190014 58294 190082 58350
rect 190138 58294 190206 58350
rect 190262 58294 220554 58350
rect 220610 58294 220678 58350
rect 220734 58294 220802 58350
rect 220858 58294 220926 58350
rect 220982 58294 251274 58350
rect 251330 58294 251398 58350
rect 251454 58294 251522 58350
rect 251578 58294 251646 58350
rect 251702 58294 281994 58350
rect 282050 58294 282118 58350
rect 282174 58294 282242 58350
rect 282298 58294 282366 58350
rect 282422 58294 312714 58350
rect 312770 58294 312838 58350
rect 312894 58294 312962 58350
rect 313018 58294 313086 58350
rect 313142 58294 343434 58350
rect 343490 58294 343558 58350
rect 343614 58294 343682 58350
rect 343738 58294 343806 58350
rect 343862 58294 374154 58350
rect 374210 58294 374278 58350
rect 374334 58294 374402 58350
rect 374458 58294 374526 58350
rect 374582 58294 404874 58350
rect 404930 58294 404998 58350
rect 405054 58294 405122 58350
rect 405178 58294 405246 58350
rect 405302 58294 435594 58350
rect 435650 58294 435718 58350
rect 435774 58294 435842 58350
rect 435898 58294 435966 58350
rect 436022 58294 466314 58350
rect 466370 58294 466438 58350
rect 466494 58294 466562 58350
rect 466618 58294 466686 58350
rect 466742 58294 497034 58350
rect 497090 58294 497158 58350
rect 497214 58294 497282 58350
rect 497338 58294 497406 58350
rect 497462 58294 527754 58350
rect 527810 58294 527878 58350
rect 527934 58294 528002 58350
rect 528058 58294 528126 58350
rect 528182 58294 558474 58350
rect 558530 58294 558598 58350
rect 558654 58294 558722 58350
rect 558778 58294 558846 58350
rect 558902 58294 589194 58350
rect 589250 58294 589318 58350
rect 589374 58294 589442 58350
rect 589498 58294 589566 58350
rect 589622 58294 596496 58350
rect 596552 58294 596620 58350
rect 596676 58294 596744 58350
rect 596800 58294 596868 58350
rect 596924 58294 597980 58350
rect -1916 58226 597980 58294
rect -1916 58170 -860 58226
rect -804 58170 -736 58226
rect -680 58170 -612 58226
rect -556 58170 -488 58226
rect -432 58170 5514 58226
rect 5570 58170 5638 58226
rect 5694 58170 5762 58226
rect 5818 58170 5886 58226
rect 5942 58170 16518 58226
rect 16574 58170 16642 58226
rect 16698 58170 36234 58226
rect 36290 58170 36358 58226
rect 36414 58170 36482 58226
rect 36538 58170 36606 58226
rect 36662 58170 47238 58226
rect 47294 58170 47362 58226
rect 47418 58170 66954 58226
rect 67010 58170 67078 58226
rect 67134 58170 67202 58226
rect 67258 58170 67326 58226
rect 67382 58170 77958 58226
rect 78014 58170 78082 58226
rect 78138 58170 97674 58226
rect 97730 58170 97798 58226
rect 97854 58170 97922 58226
rect 97978 58170 98046 58226
rect 98102 58170 108678 58226
rect 108734 58170 108802 58226
rect 108858 58170 128394 58226
rect 128450 58170 128518 58226
rect 128574 58170 128642 58226
rect 128698 58170 128766 58226
rect 128822 58170 159114 58226
rect 159170 58170 159238 58226
rect 159294 58170 159362 58226
rect 159418 58170 159486 58226
rect 159542 58170 189834 58226
rect 189890 58170 189958 58226
rect 190014 58170 190082 58226
rect 190138 58170 190206 58226
rect 190262 58170 220554 58226
rect 220610 58170 220678 58226
rect 220734 58170 220802 58226
rect 220858 58170 220926 58226
rect 220982 58170 251274 58226
rect 251330 58170 251398 58226
rect 251454 58170 251522 58226
rect 251578 58170 251646 58226
rect 251702 58170 281994 58226
rect 282050 58170 282118 58226
rect 282174 58170 282242 58226
rect 282298 58170 282366 58226
rect 282422 58170 312714 58226
rect 312770 58170 312838 58226
rect 312894 58170 312962 58226
rect 313018 58170 313086 58226
rect 313142 58170 343434 58226
rect 343490 58170 343558 58226
rect 343614 58170 343682 58226
rect 343738 58170 343806 58226
rect 343862 58170 374154 58226
rect 374210 58170 374278 58226
rect 374334 58170 374402 58226
rect 374458 58170 374526 58226
rect 374582 58170 404874 58226
rect 404930 58170 404998 58226
rect 405054 58170 405122 58226
rect 405178 58170 405246 58226
rect 405302 58170 435594 58226
rect 435650 58170 435718 58226
rect 435774 58170 435842 58226
rect 435898 58170 435966 58226
rect 436022 58170 466314 58226
rect 466370 58170 466438 58226
rect 466494 58170 466562 58226
rect 466618 58170 466686 58226
rect 466742 58170 497034 58226
rect 497090 58170 497158 58226
rect 497214 58170 497282 58226
rect 497338 58170 497406 58226
rect 497462 58170 527754 58226
rect 527810 58170 527878 58226
rect 527934 58170 528002 58226
rect 528058 58170 528126 58226
rect 528182 58170 558474 58226
rect 558530 58170 558598 58226
rect 558654 58170 558722 58226
rect 558778 58170 558846 58226
rect 558902 58170 589194 58226
rect 589250 58170 589318 58226
rect 589374 58170 589442 58226
rect 589498 58170 589566 58226
rect 589622 58170 596496 58226
rect 596552 58170 596620 58226
rect 596676 58170 596744 58226
rect 596800 58170 596868 58226
rect 596924 58170 597980 58226
rect -1916 58102 597980 58170
rect -1916 58046 -860 58102
rect -804 58046 -736 58102
rect -680 58046 -612 58102
rect -556 58046 -488 58102
rect -432 58046 5514 58102
rect 5570 58046 5638 58102
rect 5694 58046 5762 58102
rect 5818 58046 5886 58102
rect 5942 58046 16518 58102
rect 16574 58046 16642 58102
rect 16698 58046 36234 58102
rect 36290 58046 36358 58102
rect 36414 58046 36482 58102
rect 36538 58046 36606 58102
rect 36662 58046 47238 58102
rect 47294 58046 47362 58102
rect 47418 58046 66954 58102
rect 67010 58046 67078 58102
rect 67134 58046 67202 58102
rect 67258 58046 67326 58102
rect 67382 58046 77958 58102
rect 78014 58046 78082 58102
rect 78138 58046 97674 58102
rect 97730 58046 97798 58102
rect 97854 58046 97922 58102
rect 97978 58046 98046 58102
rect 98102 58046 108678 58102
rect 108734 58046 108802 58102
rect 108858 58046 128394 58102
rect 128450 58046 128518 58102
rect 128574 58046 128642 58102
rect 128698 58046 128766 58102
rect 128822 58046 159114 58102
rect 159170 58046 159238 58102
rect 159294 58046 159362 58102
rect 159418 58046 159486 58102
rect 159542 58046 189834 58102
rect 189890 58046 189958 58102
rect 190014 58046 190082 58102
rect 190138 58046 190206 58102
rect 190262 58046 220554 58102
rect 220610 58046 220678 58102
rect 220734 58046 220802 58102
rect 220858 58046 220926 58102
rect 220982 58046 251274 58102
rect 251330 58046 251398 58102
rect 251454 58046 251522 58102
rect 251578 58046 251646 58102
rect 251702 58046 281994 58102
rect 282050 58046 282118 58102
rect 282174 58046 282242 58102
rect 282298 58046 282366 58102
rect 282422 58046 312714 58102
rect 312770 58046 312838 58102
rect 312894 58046 312962 58102
rect 313018 58046 313086 58102
rect 313142 58046 343434 58102
rect 343490 58046 343558 58102
rect 343614 58046 343682 58102
rect 343738 58046 343806 58102
rect 343862 58046 374154 58102
rect 374210 58046 374278 58102
rect 374334 58046 374402 58102
rect 374458 58046 374526 58102
rect 374582 58046 404874 58102
rect 404930 58046 404998 58102
rect 405054 58046 405122 58102
rect 405178 58046 405246 58102
rect 405302 58046 435594 58102
rect 435650 58046 435718 58102
rect 435774 58046 435842 58102
rect 435898 58046 435966 58102
rect 436022 58046 466314 58102
rect 466370 58046 466438 58102
rect 466494 58046 466562 58102
rect 466618 58046 466686 58102
rect 466742 58046 497034 58102
rect 497090 58046 497158 58102
rect 497214 58046 497282 58102
rect 497338 58046 497406 58102
rect 497462 58046 527754 58102
rect 527810 58046 527878 58102
rect 527934 58046 528002 58102
rect 528058 58046 528126 58102
rect 528182 58046 558474 58102
rect 558530 58046 558598 58102
rect 558654 58046 558722 58102
rect 558778 58046 558846 58102
rect 558902 58046 589194 58102
rect 589250 58046 589318 58102
rect 589374 58046 589442 58102
rect 589498 58046 589566 58102
rect 589622 58046 596496 58102
rect 596552 58046 596620 58102
rect 596676 58046 596744 58102
rect 596800 58046 596868 58102
rect 596924 58046 597980 58102
rect -1916 57978 597980 58046
rect -1916 57922 -860 57978
rect -804 57922 -736 57978
rect -680 57922 -612 57978
rect -556 57922 -488 57978
rect -432 57922 5514 57978
rect 5570 57922 5638 57978
rect 5694 57922 5762 57978
rect 5818 57922 5886 57978
rect 5942 57922 16518 57978
rect 16574 57922 16642 57978
rect 16698 57922 36234 57978
rect 36290 57922 36358 57978
rect 36414 57922 36482 57978
rect 36538 57922 36606 57978
rect 36662 57922 47238 57978
rect 47294 57922 47362 57978
rect 47418 57922 66954 57978
rect 67010 57922 67078 57978
rect 67134 57922 67202 57978
rect 67258 57922 67326 57978
rect 67382 57922 77958 57978
rect 78014 57922 78082 57978
rect 78138 57922 97674 57978
rect 97730 57922 97798 57978
rect 97854 57922 97922 57978
rect 97978 57922 98046 57978
rect 98102 57922 108678 57978
rect 108734 57922 108802 57978
rect 108858 57922 128394 57978
rect 128450 57922 128518 57978
rect 128574 57922 128642 57978
rect 128698 57922 128766 57978
rect 128822 57922 159114 57978
rect 159170 57922 159238 57978
rect 159294 57922 159362 57978
rect 159418 57922 159486 57978
rect 159542 57922 189834 57978
rect 189890 57922 189958 57978
rect 190014 57922 190082 57978
rect 190138 57922 190206 57978
rect 190262 57922 220554 57978
rect 220610 57922 220678 57978
rect 220734 57922 220802 57978
rect 220858 57922 220926 57978
rect 220982 57922 251274 57978
rect 251330 57922 251398 57978
rect 251454 57922 251522 57978
rect 251578 57922 251646 57978
rect 251702 57922 281994 57978
rect 282050 57922 282118 57978
rect 282174 57922 282242 57978
rect 282298 57922 282366 57978
rect 282422 57922 312714 57978
rect 312770 57922 312838 57978
rect 312894 57922 312962 57978
rect 313018 57922 313086 57978
rect 313142 57922 343434 57978
rect 343490 57922 343558 57978
rect 343614 57922 343682 57978
rect 343738 57922 343806 57978
rect 343862 57922 374154 57978
rect 374210 57922 374278 57978
rect 374334 57922 374402 57978
rect 374458 57922 374526 57978
rect 374582 57922 404874 57978
rect 404930 57922 404998 57978
rect 405054 57922 405122 57978
rect 405178 57922 405246 57978
rect 405302 57922 435594 57978
rect 435650 57922 435718 57978
rect 435774 57922 435842 57978
rect 435898 57922 435966 57978
rect 436022 57922 466314 57978
rect 466370 57922 466438 57978
rect 466494 57922 466562 57978
rect 466618 57922 466686 57978
rect 466742 57922 497034 57978
rect 497090 57922 497158 57978
rect 497214 57922 497282 57978
rect 497338 57922 497406 57978
rect 497462 57922 527754 57978
rect 527810 57922 527878 57978
rect 527934 57922 528002 57978
rect 528058 57922 528126 57978
rect 528182 57922 558474 57978
rect 558530 57922 558598 57978
rect 558654 57922 558722 57978
rect 558778 57922 558846 57978
rect 558902 57922 589194 57978
rect 589250 57922 589318 57978
rect 589374 57922 589442 57978
rect 589498 57922 589566 57978
rect 589622 57922 596496 57978
rect 596552 57922 596620 57978
rect 596676 57922 596744 57978
rect 596800 57922 596868 57978
rect 596924 57922 597980 57978
rect -1916 57826 597980 57922
rect 92748 57358 509140 57374
rect 92748 57302 92764 57358
rect 92820 57302 509068 57358
rect 509124 57302 509140 57358
rect 92748 57286 509140 57302
rect 96444 57178 539380 57194
rect 96444 57122 96460 57178
rect 96516 57122 539308 57178
rect 539364 57122 539380 57178
rect 96444 57106 539380 57122
rect 12332 56998 24404 57014
rect 12332 56942 12348 56998
rect 12404 56942 24332 56998
rect 24388 56942 24404 56998
rect 12332 56926 24404 56942
rect 66428 56458 110868 56474
rect 66428 56402 66444 56458
rect 66500 56402 110796 56458
rect 110852 56402 110868 56458
rect 66428 56386 110868 56402
rect 53660 56278 91716 56294
rect 53660 56222 53676 56278
rect 53732 56222 91644 56278
rect 91700 56222 91716 56278
rect 53660 56206 91716 56222
rect 91628 56098 265540 56114
rect 91628 56042 91644 56098
rect 91700 56042 265468 56098
rect 265524 56042 265540 56098
rect 91628 56026 265540 56042
rect 79980 55918 376420 55934
rect 79980 55862 79996 55918
rect 80052 55862 376348 55918
rect 376404 55862 376420 55918
rect 79980 55846 376420 55862
rect 95436 55738 522580 55754
rect 95436 55682 95452 55738
rect 95508 55682 522508 55738
rect 522564 55682 522580 55738
rect 95436 55666 522580 55682
rect 99356 55558 561220 55574
rect 99356 55502 99372 55558
rect 99428 55502 561148 55558
rect 561204 55502 561220 55558
rect 99356 55486 561220 55502
rect 78524 55018 83204 55034
rect 78524 54962 78540 55018
rect 78596 54962 83132 55018
rect 83188 54962 83204 55018
rect 78524 54946 83204 54962
rect 69452 54838 83428 54854
rect 69452 54782 69468 54838
rect 69524 54782 83356 54838
rect 83412 54782 83428 54838
rect 69452 54766 83428 54782
rect 12332 54658 26084 54674
rect 12332 54602 12348 54658
rect 12404 54602 26012 54658
rect 26068 54602 26084 54658
rect 12332 54586 26084 54602
rect 57692 54658 94964 54674
rect 57692 54602 57708 54658
rect 57764 54602 94892 54658
rect 94948 54602 94964 54658
rect 57692 54586 94964 54602
rect 96556 54658 120164 54674
rect 96556 54602 96572 54658
rect 96628 54602 120092 54658
rect 120148 54602 120164 54658
rect 96556 54586 120164 54602
rect 87036 54478 453700 54494
rect 87036 54422 87052 54478
rect 87108 54422 453628 54478
rect 453684 54422 453700 54478
rect 87036 54406 453700 54422
rect 90396 54298 487300 54314
rect 90396 54242 90412 54298
rect 90468 54242 487228 54298
rect 487284 54242 487300 54298
rect 90396 54226 487300 54242
rect 94876 54118 510820 54134
rect 94876 54062 94892 54118
rect 94948 54062 510748 54118
rect 510804 54062 510820 54118
rect 94876 54046 510820 54062
rect 100476 53938 566260 53954
rect 100476 53882 100492 53938
rect 100548 53882 566188 53938
rect 566244 53882 566260 53938
rect 100476 53866 566260 53882
rect 12668 53758 17684 53774
rect 12668 53702 12684 53758
rect 12740 53702 17612 53758
rect 17668 53702 17684 53758
rect 12668 53686 17684 53702
rect 79756 53038 96644 53054
rect 79756 52982 79772 53038
rect 79828 52982 96572 53038
rect 96628 52982 96644 53038
rect 79756 52966 96644 52982
rect 61052 52858 91828 52874
rect 61052 52802 61068 52858
rect 61124 52802 91756 52858
rect 91812 52802 91828 52858
rect 61052 52786 91828 52802
rect 68556 52678 290740 52694
rect 68556 52622 68572 52678
rect 68628 52622 290668 52678
rect 290724 52622 290740 52678
rect 68556 52606 290740 52622
rect 88716 52498 465460 52514
rect 88716 52442 88732 52498
rect 88788 52442 465388 52498
rect 465444 52442 465460 52498
rect 88716 52426 465460 52442
rect 94204 52318 517540 52334
rect 94204 52262 94220 52318
rect 94276 52262 517468 52318
rect 517524 52262 517540 52318
rect 94204 52246 517540 52262
rect 98572 52138 554500 52154
rect 98572 52082 98588 52138
rect 98644 52082 554428 52138
rect 554484 52082 554500 52138
rect 98572 52066 554500 52082
rect 12332 51958 22724 51974
rect 12332 51902 12348 51958
rect 12404 51902 22652 51958
rect 22708 51902 22724 51958
rect 12332 51886 22724 51902
rect 72028 51598 84996 51614
rect 72028 51542 72044 51598
rect 72100 51542 84924 51598
rect 84980 51542 84996 51598
rect 72028 51526 84996 51542
rect 57020 51418 78500 51434
rect 57020 51362 57036 51418
rect 57092 51362 78428 51418
rect 78484 51362 78500 51418
rect 57020 51346 78500 51362
rect 73932 51238 134500 51254
rect 73932 51182 73948 51238
rect 74004 51182 134428 51238
rect 134484 51182 134500 51238
rect 73932 51166 134500 51182
rect 85468 51058 436900 51074
rect 85468 51002 85484 51058
rect 85540 51002 436828 51058
rect 436884 51002 436900 51058
rect 85468 50986 436900 51002
rect 89276 50878 475540 50894
rect 89276 50822 89292 50878
rect 89348 50822 475468 50878
rect 475524 50822 475540 50878
rect 89276 50806 475540 50822
rect 96220 50698 534340 50714
rect 96220 50642 96236 50698
rect 96292 50642 534268 50698
rect 534324 50642 534340 50698
rect 96220 50626 534340 50642
rect 97340 50518 537700 50534
rect 97340 50462 97356 50518
rect 97412 50462 537628 50518
rect 537684 50462 537700 50518
rect 97340 50446 537700 50462
rect 9980 49618 27764 49634
rect 9980 49562 9996 49618
rect 10052 49562 27692 49618
rect 27748 49562 27764 49618
rect 9980 49546 27764 49562
rect 64412 49618 88356 49634
rect 64412 49562 64428 49618
rect 64484 49562 88284 49618
rect 88340 49562 88356 49618
rect 64412 49546 88356 49562
rect 110780 49618 282676 49634
rect 110780 49562 110796 49618
rect 110852 49562 282604 49618
rect 282660 49562 282676 49618
rect 110780 49546 282676 49562
rect 88156 49078 443620 49094
rect 88156 49022 88172 49078
rect 88228 49022 443548 49078
rect 443604 49022 443620 49078
rect 88156 49006 443620 49022
rect 98684 48898 549460 48914
rect 98684 48842 98700 48898
rect 98756 48842 549388 48898
rect 549444 48842 549460 48898
rect 98684 48826 549460 48842
rect 12668 48718 19364 48734
rect 12668 48662 12684 48718
rect 12740 48662 19292 48718
rect 19348 48662 19364 48718
rect 12668 48646 19364 48662
rect 78412 48718 81636 48734
rect 78412 48662 78428 48718
rect 78484 48662 81564 48718
rect 81620 48662 81636 48718
rect 78412 48646 81636 48662
rect 49180 47818 74020 47834
rect 49180 47762 49196 47818
rect 49252 47762 73948 47818
rect 74004 47762 74020 47818
rect 49180 47746 74020 47762
rect 59484 47638 221860 47654
rect 59484 47582 59500 47638
rect 59556 47582 221788 47638
rect 221844 47582 221860 47638
rect 59484 47566 221860 47582
rect 86140 47458 448660 47474
rect 86140 47402 86156 47458
rect 86212 47402 448588 47458
rect 448644 47402 448660 47458
rect 86140 47386 448660 47402
rect 90844 47278 488980 47294
rect 90844 47222 90860 47278
rect 90916 47222 488908 47278
rect 488964 47222 488980 47278
rect 90844 47206 488980 47222
rect 95996 47098 532660 47114
rect 95996 47042 96012 47098
rect 96068 47042 532588 47098
rect 532644 47042 532660 47098
rect 95996 47026 532660 47042
rect -1916 46350 597980 46446
rect -1916 46294 -1820 46350
rect -1764 46294 -1696 46350
rect -1640 46294 -1572 46350
rect -1516 46294 -1448 46350
rect -1392 46294 9234 46350
rect 9290 46294 9358 46350
rect 9414 46294 9482 46350
rect 9538 46294 9606 46350
rect 9662 46294 31878 46350
rect 31934 46294 32002 46350
rect 32058 46294 39954 46350
rect 40010 46294 40078 46350
rect 40134 46294 40202 46350
rect 40258 46294 40326 46350
rect 40382 46294 62598 46350
rect 62654 46294 62722 46350
rect 62778 46294 70674 46350
rect 70730 46294 70798 46350
rect 70854 46294 70922 46350
rect 70978 46294 71046 46350
rect 71102 46294 93318 46350
rect 93374 46294 93442 46350
rect 93498 46294 101394 46350
rect 101450 46294 101518 46350
rect 101574 46294 101642 46350
rect 101698 46294 101766 46350
rect 101822 46294 132114 46350
rect 132170 46294 132238 46350
rect 132294 46294 132362 46350
rect 132418 46294 132486 46350
rect 132542 46294 162834 46350
rect 162890 46294 162958 46350
rect 163014 46294 163082 46350
rect 163138 46294 163206 46350
rect 163262 46294 193554 46350
rect 193610 46294 193678 46350
rect 193734 46294 193802 46350
rect 193858 46294 193926 46350
rect 193982 46294 224274 46350
rect 224330 46294 224398 46350
rect 224454 46294 224522 46350
rect 224578 46294 224646 46350
rect 224702 46294 254994 46350
rect 255050 46294 255118 46350
rect 255174 46294 255242 46350
rect 255298 46294 255366 46350
rect 255422 46294 285714 46350
rect 285770 46294 285838 46350
rect 285894 46294 285962 46350
rect 286018 46294 286086 46350
rect 286142 46294 316434 46350
rect 316490 46294 316558 46350
rect 316614 46294 316682 46350
rect 316738 46294 316806 46350
rect 316862 46294 347154 46350
rect 347210 46294 347278 46350
rect 347334 46294 347402 46350
rect 347458 46294 347526 46350
rect 347582 46294 377874 46350
rect 377930 46294 377998 46350
rect 378054 46294 378122 46350
rect 378178 46294 378246 46350
rect 378302 46294 408594 46350
rect 408650 46294 408718 46350
rect 408774 46294 408842 46350
rect 408898 46294 408966 46350
rect 409022 46294 439314 46350
rect 439370 46294 439438 46350
rect 439494 46294 439562 46350
rect 439618 46294 439686 46350
rect 439742 46294 470034 46350
rect 470090 46294 470158 46350
rect 470214 46294 470282 46350
rect 470338 46294 470406 46350
rect 470462 46294 500754 46350
rect 500810 46294 500878 46350
rect 500934 46294 501002 46350
rect 501058 46294 501126 46350
rect 501182 46294 531474 46350
rect 531530 46294 531598 46350
rect 531654 46294 531722 46350
rect 531778 46294 531846 46350
rect 531902 46294 562194 46350
rect 562250 46294 562318 46350
rect 562374 46294 562442 46350
rect 562498 46294 562566 46350
rect 562622 46294 592914 46350
rect 592970 46294 593038 46350
rect 593094 46294 593162 46350
rect 593218 46294 593286 46350
rect 593342 46294 597456 46350
rect 597512 46294 597580 46350
rect 597636 46294 597704 46350
rect 597760 46294 597828 46350
rect 597884 46294 597980 46350
rect -1916 46226 597980 46294
rect -1916 46170 -1820 46226
rect -1764 46170 -1696 46226
rect -1640 46170 -1572 46226
rect -1516 46170 -1448 46226
rect -1392 46170 9234 46226
rect 9290 46170 9358 46226
rect 9414 46170 9482 46226
rect 9538 46170 9606 46226
rect 9662 46170 31878 46226
rect 31934 46170 32002 46226
rect 32058 46170 39954 46226
rect 40010 46170 40078 46226
rect 40134 46170 40202 46226
rect 40258 46170 40326 46226
rect 40382 46170 62598 46226
rect 62654 46170 62722 46226
rect 62778 46170 70674 46226
rect 70730 46170 70798 46226
rect 70854 46170 70922 46226
rect 70978 46170 71046 46226
rect 71102 46170 93318 46226
rect 93374 46170 93442 46226
rect 93498 46170 101394 46226
rect 101450 46170 101518 46226
rect 101574 46170 101642 46226
rect 101698 46170 101766 46226
rect 101822 46170 132114 46226
rect 132170 46170 132238 46226
rect 132294 46170 132362 46226
rect 132418 46170 132486 46226
rect 132542 46170 162834 46226
rect 162890 46170 162958 46226
rect 163014 46170 163082 46226
rect 163138 46170 163206 46226
rect 163262 46170 193554 46226
rect 193610 46170 193678 46226
rect 193734 46170 193802 46226
rect 193858 46170 193926 46226
rect 193982 46170 224274 46226
rect 224330 46170 224398 46226
rect 224454 46170 224522 46226
rect 224578 46170 224646 46226
rect 224702 46170 254994 46226
rect 255050 46170 255118 46226
rect 255174 46170 255242 46226
rect 255298 46170 255366 46226
rect 255422 46170 285714 46226
rect 285770 46170 285838 46226
rect 285894 46170 285962 46226
rect 286018 46170 286086 46226
rect 286142 46170 316434 46226
rect 316490 46170 316558 46226
rect 316614 46170 316682 46226
rect 316738 46170 316806 46226
rect 316862 46170 347154 46226
rect 347210 46170 347278 46226
rect 347334 46170 347402 46226
rect 347458 46170 347526 46226
rect 347582 46170 377874 46226
rect 377930 46170 377998 46226
rect 378054 46170 378122 46226
rect 378178 46170 378246 46226
rect 378302 46170 408594 46226
rect 408650 46170 408718 46226
rect 408774 46170 408842 46226
rect 408898 46170 408966 46226
rect 409022 46170 439314 46226
rect 439370 46170 439438 46226
rect 439494 46170 439562 46226
rect 439618 46170 439686 46226
rect 439742 46170 470034 46226
rect 470090 46170 470158 46226
rect 470214 46170 470282 46226
rect 470338 46170 470406 46226
rect 470462 46170 500754 46226
rect 500810 46170 500878 46226
rect 500934 46170 501002 46226
rect 501058 46170 501126 46226
rect 501182 46170 531474 46226
rect 531530 46170 531598 46226
rect 531654 46170 531722 46226
rect 531778 46170 531846 46226
rect 531902 46170 562194 46226
rect 562250 46170 562318 46226
rect 562374 46170 562442 46226
rect 562498 46170 562566 46226
rect 562622 46170 592914 46226
rect 592970 46170 593038 46226
rect 593094 46170 593162 46226
rect 593218 46170 593286 46226
rect 593342 46170 597456 46226
rect 597512 46170 597580 46226
rect 597636 46170 597704 46226
rect 597760 46170 597828 46226
rect 597884 46170 597980 46226
rect -1916 46102 597980 46170
rect -1916 46046 -1820 46102
rect -1764 46046 -1696 46102
rect -1640 46046 -1572 46102
rect -1516 46046 -1448 46102
rect -1392 46046 9234 46102
rect 9290 46046 9358 46102
rect 9414 46046 9482 46102
rect 9538 46046 9606 46102
rect 9662 46046 31878 46102
rect 31934 46046 32002 46102
rect 32058 46046 39954 46102
rect 40010 46046 40078 46102
rect 40134 46046 40202 46102
rect 40258 46046 40326 46102
rect 40382 46046 62598 46102
rect 62654 46046 62722 46102
rect 62778 46046 70674 46102
rect 70730 46046 70798 46102
rect 70854 46046 70922 46102
rect 70978 46046 71046 46102
rect 71102 46046 93318 46102
rect 93374 46046 93442 46102
rect 93498 46046 101394 46102
rect 101450 46046 101518 46102
rect 101574 46046 101642 46102
rect 101698 46046 101766 46102
rect 101822 46046 132114 46102
rect 132170 46046 132238 46102
rect 132294 46046 132362 46102
rect 132418 46046 132486 46102
rect 132542 46046 162834 46102
rect 162890 46046 162958 46102
rect 163014 46046 163082 46102
rect 163138 46046 163206 46102
rect 163262 46046 193554 46102
rect 193610 46046 193678 46102
rect 193734 46046 193802 46102
rect 193858 46046 193926 46102
rect 193982 46046 224274 46102
rect 224330 46046 224398 46102
rect 224454 46046 224522 46102
rect 224578 46046 224646 46102
rect 224702 46046 254994 46102
rect 255050 46046 255118 46102
rect 255174 46046 255242 46102
rect 255298 46046 255366 46102
rect 255422 46046 285714 46102
rect 285770 46046 285838 46102
rect 285894 46046 285962 46102
rect 286018 46046 286086 46102
rect 286142 46046 316434 46102
rect 316490 46046 316558 46102
rect 316614 46046 316682 46102
rect 316738 46046 316806 46102
rect 316862 46046 347154 46102
rect 347210 46046 347278 46102
rect 347334 46046 347402 46102
rect 347458 46046 347526 46102
rect 347582 46046 377874 46102
rect 377930 46046 377998 46102
rect 378054 46046 378122 46102
rect 378178 46046 378246 46102
rect 378302 46046 408594 46102
rect 408650 46046 408718 46102
rect 408774 46046 408842 46102
rect 408898 46046 408966 46102
rect 409022 46046 439314 46102
rect 439370 46046 439438 46102
rect 439494 46046 439562 46102
rect 439618 46046 439686 46102
rect 439742 46046 470034 46102
rect 470090 46046 470158 46102
rect 470214 46046 470282 46102
rect 470338 46046 470406 46102
rect 470462 46046 500754 46102
rect 500810 46046 500878 46102
rect 500934 46046 501002 46102
rect 501058 46046 501126 46102
rect 501182 46046 531474 46102
rect 531530 46046 531598 46102
rect 531654 46046 531722 46102
rect 531778 46046 531846 46102
rect 531902 46046 562194 46102
rect 562250 46046 562318 46102
rect 562374 46046 562442 46102
rect 562498 46046 562566 46102
rect 562622 46046 592914 46102
rect 592970 46046 593038 46102
rect 593094 46046 593162 46102
rect 593218 46046 593286 46102
rect 593342 46046 597456 46102
rect 597512 46046 597580 46102
rect 597636 46046 597704 46102
rect 597760 46046 597828 46102
rect 597884 46046 597980 46102
rect -1916 45978 597980 46046
rect -1916 45922 -1820 45978
rect -1764 45922 -1696 45978
rect -1640 45922 -1572 45978
rect -1516 45922 -1448 45978
rect -1392 45922 9234 45978
rect 9290 45922 9358 45978
rect 9414 45922 9482 45978
rect 9538 45922 9606 45978
rect 9662 45922 31878 45978
rect 31934 45922 32002 45978
rect 32058 45922 39954 45978
rect 40010 45922 40078 45978
rect 40134 45922 40202 45978
rect 40258 45922 40326 45978
rect 40382 45922 62598 45978
rect 62654 45922 62722 45978
rect 62778 45922 70674 45978
rect 70730 45922 70798 45978
rect 70854 45922 70922 45978
rect 70978 45922 71046 45978
rect 71102 45922 93318 45978
rect 93374 45922 93442 45978
rect 93498 45922 101394 45978
rect 101450 45922 101518 45978
rect 101574 45922 101642 45978
rect 101698 45922 101766 45978
rect 101822 45922 132114 45978
rect 132170 45922 132238 45978
rect 132294 45922 132362 45978
rect 132418 45922 132486 45978
rect 132542 45922 162834 45978
rect 162890 45922 162958 45978
rect 163014 45922 163082 45978
rect 163138 45922 163206 45978
rect 163262 45922 193554 45978
rect 193610 45922 193678 45978
rect 193734 45922 193802 45978
rect 193858 45922 193926 45978
rect 193982 45922 224274 45978
rect 224330 45922 224398 45978
rect 224454 45922 224522 45978
rect 224578 45922 224646 45978
rect 224702 45922 254994 45978
rect 255050 45922 255118 45978
rect 255174 45922 255242 45978
rect 255298 45922 255366 45978
rect 255422 45922 285714 45978
rect 285770 45922 285838 45978
rect 285894 45922 285962 45978
rect 286018 45922 286086 45978
rect 286142 45922 316434 45978
rect 316490 45922 316558 45978
rect 316614 45922 316682 45978
rect 316738 45922 316806 45978
rect 316862 45922 347154 45978
rect 347210 45922 347278 45978
rect 347334 45922 347402 45978
rect 347458 45922 347526 45978
rect 347582 45922 377874 45978
rect 377930 45922 377998 45978
rect 378054 45922 378122 45978
rect 378178 45922 378246 45978
rect 378302 45922 408594 45978
rect 408650 45922 408718 45978
rect 408774 45922 408842 45978
rect 408898 45922 408966 45978
rect 409022 45922 439314 45978
rect 439370 45922 439438 45978
rect 439494 45922 439562 45978
rect 439618 45922 439686 45978
rect 439742 45922 470034 45978
rect 470090 45922 470158 45978
rect 470214 45922 470282 45978
rect 470338 45922 470406 45978
rect 470462 45922 500754 45978
rect 500810 45922 500878 45978
rect 500934 45922 501002 45978
rect 501058 45922 501126 45978
rect 501182 45922 531474 45978
rect 531530 45922 531598 45978
rect 531654 45922 531722 45978
rect 531778 45922 531846 45978
rect 531902 45922 562194 45978
rect 562250 45922 562318 45978
rect 562374 45922 562442 45978
rect 562498 45922 562566 45978
rect 562622 45922 592914 45978
rect 592970 45922 593038 45978
rect 593094 45922 593162 45978
rect 593218 45922 593286 45978
rect 593342 45922 597456 45978
rect 597512 45922 597580 45978
rect 597636 45922 597704 45978
rect 597760 45922 597828 45978
rect 597884 45922 597980 45978
rect -1916 45826 597980 45922
rect 75500 45658 126100 45674
rect 75500 45602 75516 45658
rect 75572 45602 126028 45658
rect 126084 45602 126100 45658
rect 75500 45586 126100 45602
rect 90732 45478 190500 45494
rect 90732 45422 90748 45478
rect 90804 45422 190428 45478
rect 190484 45422 190500 45478
rect 90732 45406 190500 45422
rect 63516 44758 79956 44774
rect 63516 44702 63532 44758
rect 63588 44702 79884 44758
rect 79940 44702 79956 44758
rect 63516 44686 79956 44702
rect 48956 44578 132820 44594
rect 48956 44522 48972 44578
rect 49028 44522 132748 44578
rect 132804 44522 132820 44578
rect 48956 44506 132820 44522
rect 83116 44398 319300 44414
rect 83116 44342 83132 44398
rect 83188 44342 319228 44398
rect 319284 44342 319300 44398
rect 83116 44326 319300 44342
rect 95324 44218 364660 44234
rect 95324 44162 95340 44218
rect 95396 44162 364588 44218
rect 364644 44162 364660 44218
rect 95324 44146 364660 44162
rect 81660 44038 352900 44054
rect 81660 43982 81676 44038
rect 81732 43982 352828 44038
rect 352884 43982 352900 44038
rect 81660 43966 352900 43982
rect 75276 43858 351220 43874
rect 75276 43802 75292 43858
rect 75348 43802 351148 43858
rect 351204 43802 351220 43858
rect 75276 43786 351220 43802
rect 55676 42778 90820 42794
rect 55676 42722 55692 42778
rect 55748 42722 90748 42778
rect 90804 42722 90820 42778
rect 55676 42706 90820 42722
rect 120076 42778 346180 42794
rect 120076 42722 120092 42778
rect 120148 42722 346108 42778
rect 346164 42722 346180 42778
rect 120076 42706 346180 42722
rect 72924 42418 260500 42434
rect 72924 42362 72940 42418
rect 72996 42362 260428 42418
rect 260484 42362 260500 42418
rect 72924 42346 260500 42362
rect 76060 42238 362980 42254
rect 76060 42182 76076 42238
rect 76132 42182 362908 42238
rect 362964 42182 362980 42238
rect 76060 42166 362980 42182
rect 100028 42058 416740 42074
rect 100028 42002 100044 42058
rect 100100 42002 416668 42058
rect 416724 42002 416740 42058
rect 100028 41986 416740 42002
rect 81548 41338 95412 41354
rect 81548 41282 81564 41338
rect 81620 41282 95340 41338
rect 95396 41282 95412 41338
rect 81548 41266 95412 41282
rect 54108 41158 147940 41174
rect 54108 41102 54124 41158
rect 54180 41102 147868 41158
rect 147924 41102 147940 41158
rect 54108 41086 147940 41102
rect 59260 40978 220180 40994
rect 59260 40922 59276 40978
rect 59332 40922 220108 40978
rect 220164 40922 220180 40978
rect 59260 40906 220180 40922
rect 73708 40798 331060 40814
rect 73708 40742 73724 40798
rect 73780 40742 330988 40798
rect 331044 40742 331060 40798
rect 73708 40726 331060 40742
rect 97228 40618 544420 40634
rect 97228 40562 97244 40618
rect 97300 40562 544348 40618
rect 544404 40562 544420 40618
rect 97228 40546 544420 40562
rect -1916 40350 597980 40446
rect -1916 40294 -860 40350
rect -804 40294 -736 40350
rect -680 40294 -612 40350
rect -556 40294 -488 40350
rect -432 40294 5514 40350
rect 5570 40294 5638 40350
rect 5694 40294 5762 40350
rect 5818 40294 5886 40350
rect 5942 40294 16518 40350
rect 16574 40294 16642 40350
rect 16698 40294 36234 40350
rect 36290 40294 36358 40350
rect 36414 40294 36482 40350
rect 36538 40294 36606 40350
rect 36662 40294 47238 40350
rect 47294 40294 47362 40350
rect 47418 40294 66954 40350
rect 67010 40294 67078 40350
rect 67134 40294 67202 40350
rect 67258 40294 67326 40350
rect 67382 40294 77958 40350
rect 78014 40294 78082 40350
rect 78138 40294 97674 40350
rect 97730 40294 97798 40350
rect 97854 40294 97922 40350
rect 97978 40294 98046 40350
rect 98102 40294 108678 40350
rect 108734 40294 108802 40350
rect 108858 40294 128394 40350
rect 128450 40294 128518 40350
rect 128574 40294 128642 40350
rect 128698 40294 128766 40350
rect 128822 40294 159114 40350
rect 159170 40294 159238 40350
rect 159294 40294 159362 40350
rect 159418 40294 159486 40350
rect 159542 40294 189834 40350
rect 189890 40294 189958 40350
rect 190014 40294 190082 40350
rect 190138 40294 190206 40350
rect 190262 40294 220554 40350
rect 220610 40294 220678 40350
rect 220734 40294 220802 40350
rect 220858 40294 220926 40350
rect 220982 40294 251274 40350
rect 251330 40294 251398 40350
rect 251454 40294 251522 40350
rect 251578 40294 251646 40350
rect 251702 40294 281994 40350
rect 282050 40294 282118 40350
rect 282174 40294 282242 40350
rect 282298 40294 282366 40350
rect 282422 40294 312714 40350
rect 312770 40294 312838 40350
rect 312894 40294 312962 40350
rect 313018 40294 313086 40350
rect 313142 40294 343434 40350
rect 343490 40294 343558 40350
rect 343614 40294 343682 40350
rect 343738 40294 343806 40350
rect 343862 40294 374154 40350
rect 374210 40294 374278 40350
rect 374334 40294 374402 40350
rect 374458 40294 374526 40350
rect 374582 40294 404874 40350
rect 404930 40294 404998 40350
rect 405054 40294 405122 40350
rect 405178 40294 405246 40350
rect 405302 40294 435594 40350
rect 435650 40294 435718 40350
rect 435774 40294 435842 40350
rect 435898 40294 435966 40350
rect 436022 40294 466314 40350
rect 466370 40294 466438 40350
rect 466494 40294 466562 40350
rect 466618 40294 466686 40350
rect 466742 40294 497034 40350
rect 497090 40294 497158 40350
rect 497214 40294 497282 40350
rect 497338 40294 497406 40350
rect 497462 40294 527754 40350
rect 527810 40294 527878 40350
rect 527934 40294 528002 40350
rect 528058 40294 528126 40350
rect 528182 40294 558474 40350
rect 558530 40294 558598 40350
rect 558654 40294 558722 40350
rect 558778 40294 558846 40350
rect 558902 40294 589194 40350
rect 589250 40294 589318 40350
rect 589374 40294 589442 40350
rect 589498 40294 589566 40350
rect 589622 40294 596496 40350
rect 596552 40294 596620 40350
rect 596676 40294 596744 40350
rect 596800 40294 596868 40350
rect 596924 40294 597980 40350
rect -1916 40226 597980 40294
rect -1916 40170 -860 40226
rect -804 40170 -736 40226
rect -680 40170 -612 40226
rect -556 40170 -488 40226
rect -432 40170 5514 40226
rect 5570 40170 5638 40226
rect 5694 40170 5762 40226
rect 5818 40170 5886 40226
rect 5942 40170 16518 40226
rect 16574 40170 16642 40226
rect 16698 40170 36234 40226
rect 36290 40170 36358 40226
rect 36414 40170 36482 40226
rect 36538 40170 36606 40226
rect 36662 40170 47238 40226
rect 47294 40170 47362 40226
rect 47418 40170 66954 40226
rect 67010 40170 67078 40226
rect 67134 40170 67202 40226
rect 67258 40170 67326 40226
rect 67382 40170 77958 40226
rect 78014 40170 78082 40226
rect 78138 40170 97674 40226
rect 97730 40170 97798 40226
rect 97854 40170 97922 40226
rect 97978 40170 98046 40226
rect 98102 40170 108678 40226
rect 108734 40170 108802 40226
rect 108858 40170 128394 40226
rect 128450 40170 128518 40226
rect 128574 40170 128642 40226
rect 128698 40170 128766 40226
rect 128822 40170 159114 40226
rect 159170 40170 159238 40226
rect 159294 40170 159362 40226
rect 159418 40170 159486 40226
rect 159542 40170 189834 40226
rect 189890 40170 189958 40226
rect 190014 40170 190082 40226
rect 190138 40170 190206 40226
rect 190262 40170 220554 40226
rect 220610 40170 220678 40226
rect 220734 40170 220802 40226
rect 220858 40170 220926 40226
rect 220982 40170 251274 40226
rect 251330 40170 251398 40226
rect 251454 40170 251522 40226
rect 251578 40170 251646 40226
rect 251702 40170 281994 40226
rect 282050 40170 282118 40226
rect 282174 40170 282242 40226
rect 282298 40170 282366 40226
rect 282422 40170 312714 40226
rect 312770 40170 312838 40226
rect 312894 40170 312962 40226
rect 313018 40170 313086 40226
rect 313142 40170 343434 40226
rect 343490 40170 343558 40226
rect 343614 40170 343682 40226
rect 343738 40170 343806 40226
rect 343862 40170 374154 40226
rect 374210 40170 374278 40226
rect 374334 40170 374402 40226
rect 374458 40170 374526 40226
rect 374582 40170 404874 40226
rect 404930 40170 404998 40226
rect 405054 40170 405122 40226
rect 405178 40170 405246 40226
rect 405302 40170 435594 40226
rect 435650 40170 435718 40226
rect 435774 40170 435842 40226
rect 435898 40170 435966 40226
rect 436022 40170 466314 40226
rect 466370 40170 466438 40226
rect 466494 40170 466562 40226
rect 466618 40170 466686 40226
rect 466742 40170 497034 40226
rect 497090 40170 497158 40226
rect 497214 40170 497282 40226
rect 497338 40170 497406 40226
rect 497462 40170 527754 40226
rect 527810 40170 527878 40226
rect 527934 40170 528002 40226
rect 528058 40170 528126 40226
rect 528182 40170 558474 40226
rect 558530 40170 558598 40226
rect 558654 40170 558722 40226
rect 558778 40170 558846 40226
rect 558902 40170 589194 40226
rect 589250 40170 589318 40226
rect 589374 40170 589442 40226
rect 589498 40170 589566 40226
rect 589622 40170 596496 40226
rect 596552 40170 596620 40226
rect 596676 40170 596744 40226
rect 596800 40170 596868 40226
rect 596924 40170 597980 40226
rect -1916 40102 597980 40170
rect -1916 40046 -860 40102
rect -804 40046 -736 40102
rect -680 40046 -612 40102
rect -556 40046 -488 40102
rect -432 40046 5514 40102
rect 5570 40046 5638 40102
rect 5694 40046 5762 40102
rect 5818 40046 5886 40102
rect 5942 40046 16518 40102
rect 16574 40046 16642 40102
rect 16698 40046 36234 40102
rect 36290 40046 36358 40102
rect 36414 40046 36482 40102
rect 36538 40046 36606 40102
rect 36662 40046 47238 40102
rect 47294 40046 47362 40102
rect 47418 40046 66954 40102
rect 67010 40046 67078 40102
rect 67134 40046 67202 40102
rect 67258 40046 67326 40102
rect 67382 40046 77958 40102
rect 78014 40046 78082 40102
rect 78138 40046 97674 40102
rect 97730 40046 97798 40102
rect 97854 40046 97922 40102
rect 97978 40046 98046 40102
rect 98102 40046 108678 40102
rect 108734 40046 108802 40102
rect 108858 40046 128394 40102
rect 128450 40046 128518 40102
rect 128574 40046 128642 40102
rect 128698 40046 128766 40102
rect 128822 40046 159114 40102
rect 159170 40046 159238 40102
rect 159294 40046 159362 40102
rect 159418 40046 159486 40102
rect 159542 40046 189834 40102
rect 189890 40046 189958 40102
rect 190014 40046 190082 40102
rect 190138 40046 190206 40102
rect 190262 40046 220554 40102
rect 220610 40046 220678 40102
rect 220734 40046 220802 40102
rect 220858 40046 220926 40102
rect 220982 40046 251274 40102
rect 251330 40046 251398 40102
rect 251454 40046 251522 40102
rect 251578 40046 251646 40102
rect 251702 40046 281994 40102
rect 282050 40046 282118 40102
rect 282174 40046 282242 40102
rect 282298 40046 282366 40102
rect 282422 40046 312714 40102
rect 312770 40046 312838 40102
rect 312894 40046 312962 40102
rect 313018 40046 313086 40102
rect 313142 40046 343434 40102
rect 343490 40046 343558 40102
rect 343614 40046 343682 40102
rect 343738 40046 343806 40102
rect 343862 40046 374154 40102
rect 374210 40046 374278 40102
rect 374334 40046 374402 40102
rect 374458 40046 374526 40102
rect 374582 40046 404874 40102
rect 404930 40046 404998 40102
rect 405054 40046 405122 40102
rect 405178 40046 405246 40102
rect 405302 40046 435594 40102
rect 435650 40046 435718 40102
rect 435774 40046 435842 40102
rect 435898 40046 435966 40102
rect 436022 40046 466314 40102
rect 466370 40046 466438 40102
rect 466494 40046 466562 40102
rect 466618 40046 466686 40102
rect 466742 40046 497034 40102
rect 497090 40046 497158 40102
rect 497214 40046 497282 40102
rect 497338 40046 497406 40102
rect 497462 40046 527754 40102
rect 527810 40046 527878 40102
rect 527934 40046 528002 40102
rect 528058 40046 528126 40102
rect 528182 40046 558474 40102
rect 558530 40046 558598 40102
rect 558654 40046 558722 40102
rect 558778 40046 558846 40102
rect 558902 40046 589194 40102
rect 589250 40046 589318 40102
rect 589374 40046 589442 40102
rect 589498 40046 589566 40102
rect 589622 40046 596496 40102
rect 596552 40046 596620 40102
rect 596676 40046 596744 40102
rect 596800 40046 596868 40102
rect 596924 40046 597980 40102
rect -1916 39978 597980 40046
rect -1916 39922 -860 39978
rect -804 39922 -736 39978
rect -680 39922 -612 39978
rect -556 39922 -488 39978
rect -432 39922 5514 39978
rect 5570 39922 5638 39978
rect 5694 39922 5762 39978
rect 5818 39922 5886 39978
rect 5942 39922 16518 39978
rect 16574 39922 16642 39978
rect 16698 39922 36234 39978
rect 36290 39922 36358 39978
rect 36414 39922 36482 39978
rect 36538 39922 36606 39978
rect 36662 39922 47238 39978
rect 47294 39922 47362 39978
rect 47418 39922 66954 39978
rect 67010 39922 67078 39978
rect 67134 39922 67202 39978
rect 67258 39922 67326 39978
rect 67382 39922 77958 39978
rect 78014 39922 78082 39978
rect 78138 39922 97674 39978
rect 97730 39922 97798 39978
rect 97854 39922 97922 39978
rect 97978 39922 98046 39978
rect 98102 39922 108678 39978
rect 108734 39922 108802 39978
rect 108858 39922 128394 39978
rect 128450 39922 128518 39978
rect 128574 39922 128642 39978
rect 128698 39922 128766 39978
rect 128822 39922 159114 39978
rect 159170 39922 159238 39978
rect 159294 39922 159362 39978
rect 159418 39922 159486 39978
rect 159542 39922 189834 39978
rect 189890 39922 189958 39978
rect 190014 39922 190082 39978
rect 190138 39922 190206 39978
rect 190262 39922 220554 39978
rect 220610 39922 220678 39978
rect 220734 39922 220802 39978
rect 220858 39922 220926 39978
rect 220982 39922 251274 39978
rect 251330 39922 251398 39978
rect 251454 39922 251522 39978
rect 251578 39922 251646 39978
rect 251702 39922 281994 39978
rect 282050 39922 282118 39978
rect 282174 39922 282242 39978
rect 282298 39922 282366 39978
rect 282422 39922 312714 39978
rect 312770 39922 312838 39978
rect 312894 39922 312962 39978
rect 313018 39922 313086 39978
rect 313142 39922 343434 39978
rect 343490 39922 343558 39978
rect 343614 39922 343682 39978
rect 343738 39922 343806 39978
rect 343862 39922 374154 39978
rect 374210 39922 374278 39978
rect 374334 39922 374402 39978
rect 374458 39922 374526 39978
rect 374582 39922 404874 39978
rect 404930 39922 404998 39978
rect 405054 39922 405122 39978
rect 405178 39922 405246 39978
rect 405302 39922 435594 39978
rect 435650 39922 435718 39978
rect 435774 39922 435842 39978
rect 435898 39922 435966 39978
rect 436022 39922 466314 39978
rect 466370 39922 466438 39978
rect 466494 39922 466562 39978
rect 466618 39922 466686 39978
rect 466742 39922 497034 39978
rect 497090 39922 497158 39978
rect 497214 39922 497282 39978
rect 497338 39922 497406 39978
rect 497462 39922 527754 39978
rect 527810 39922 527878 39978
rect 527934 39922 528002 39978
rect 528058 39922 528126 39978
rect 528182 39922 558474 39978
rect 558530 39922 558598 39978
rect 558654 39922 558722 39978
rect 558778 39922 558846 39978
rect 558902 39922 589194 39978
rect 589250 39922 589318 39978
rect 589374 39922 589442 39978
rect 589498 39922 589566 39978
rect 589622 39922 596496 39978
rect 596552 39922 596620 39978
rect 596676 39922 596744 39978
rect 596800 39922 596868 39978
rect 596924 39922 597980 39978
rect -1916 39826 597980 39922
rect 65084 39538 91716 39554
rect 65084 39482 65100 39538
rect 65156 39482 91644 39538
rect 91700 39482 91716 39538
rect 65084 39466 91716 39482
rect 91292 38818 492340 38834
rect 91292 38762 91308 38818
rect 91364 38762 492268 38818
rect 492324 38762 492340 38818
rect 91292 38746 492340 38762
rect 51196 37738 151300 37754
rect 51196 37682 51212 37738
rect 51268 37682 151228 37738
rect 151284 37682 151300 37738
rect 51196 37666 151300 37682
rect 58364 37558 215140 37574
rect 58364 37502 58380 37558
rect 58436 37502 215068 37558
rect 215124 37502 215140 37558
rect 58364 37486 215140 37502
rect 61836 37378 231940 37394
rect 61836 37322 61852 37378
rect 61908 37322 231868 37378
rect 231924 37322 231940 37378
rect 61836 37306 231940 37322
rect 79868 37198 374852 37214
rect 79868 37142 79884 37198
rect 79940 37142 374780 37198
rect 374836 37142 374852 37198
rect 79868 37126 374852 37142
rect 84908 37018 386500 37034
rect 84908 36962 84924 37018
rect 84980 36962 386428 37018
rect 386484 36962 386500 37018
rect 84908 36946 386500 36962
rect 48172 36298 75588 36314
rect 48172 36242 48188 36298
rect 48244 36242 75516 36298
rect 75572 36242 75588 36298
rect 48172 36226 75588 36242
rect 60156 36118 228580 36134
rect 60156 36062 60172 36118
rect 60228 36062 228508 36118
rect 228564 36062 228580 36118
rect 60156 36046 228580 36062
rect 61724 35938 243700 35954
rect 61724 35882 61740 35938
rect 61796 35882 243628 35938
rect 243684 35882 243700 35938
rect 61724 35866 243700 35882
rect 74940 35758 310900 35774
rect 74940 35702 74956 35758
rect 75012 35702 310828 35758
rect 310884 35702 310900 35758
rect 74940 35686 310900 35702
rect 83788 35578 425140 35594
rect 83788 35522 83804 35578
rect 83860 35522 425068 35578
rect 425124 35522 425140 35578
rect 83788 35506 425140 35522
rect 103276 35398 505780 35414
rect 103276 35342 103292 35398
rect 103348 35342 505708 35398
rect 505764 35342 505780 35398
rect 103276 35326 505780 35342
rect 46716 34678 116020 34694
rect 46716 34622 46732 34678
rect 46788 34622 115948 34678
rect 116004 34622 116020 34678
rect 46716 34606 116020 34622
rect 63964 34498 73012 34514
rect 63964 34442 63980 34498
rect 64036 34442 72940 34498
rect 72996 34442 73012 34498
rect 63964 34426 73012 34442
rect 80540 34318 278980 34334
rect 80540 34262 80556 34318
rect 80612 34262 278908 34318
rect 278964 34262 278980 34318
rect 80540 34246 278980 34262
rect 90732 34138 379780 34154
rect 90732 34082 90748 34138
rect 90804 34082 379708 34138
rect 379764 34082 379780 34138
rect 90732 34066 379780 34082
rect 75164 33958 81748 33974
rect 75164 33902 75180 33958
rect 75236 33902 81676 33958
rect 81732 33902 81748 33958
rect 75164 33886 81748 33902
rect 115820 33958 420100 33974
rect 115820 33902 115836 33958
rect 115892 33902 420028 33958
rect 420084 33902 420100 33958
rect 115820 33886 420100 33902
rect 80764 33778 403300 33794
rect 80764 33722 80780 33778
rect 80836 33722 403228 33778
rect 403284 33722 403300 33778
rect 80764 33706 403300 33722
rect 66316 32698 80628 32714
rect 66316 32642 66332 32698
rect 66388 32642 80556 32698
rect 80612 32642 80628 32698
rect 66316 32626 80628 32642
rect 82780 32698 115908 32714
rect 82780 32642 82796 32698
rect 82852 32642 115836 32698
rect 115892 32642 115908 32698
rect 82780 32626 115908 32642
rect 54332 32518 178180 32534
rect 54332 32462 54348 32518
rect 54404 32462 178108 32518
rect 178164 32462 178180 32518
rect 54332 32446 178180 32462
rect 60828 32338 233620 32354
rect 60828 32282 60844 32338
rect 60900 32282 233548 32338
rect 233604 32282 233620 32338
rect 60828 32266 233620 32282
rect 68444 32158 300820 32174
rect 68444 32102 68460 32158
rect 68516 32102 300748 32158
rect 300804 32102 300820 32158
rect 68444 32086 300820 32102
rect 99804 31978 564580 31994
rect 99804 31922 99820 31978
rect 99876 31922 564508 31978
rect 564564 31922 564580 31978
rect 99804 31906 564580 31922
rect 46604 31258 109300 31274
rect 46604 31202 46620 31258
rect 46676 31202 109228 31258
rect 109284 31202 109300 31258
rect 46604 31186 109300 31202
rect 51980 30898 154660 30914
rect 51980 30842 51996 30898
rect 52052 30842 154588 30898
rect 154644 30842 154660 30898
rect 51980 30826 154660 30842
rect 104060 30718 342820 30734
rect 104060 30662 104076 30718
rect 104132 30662 342748 30718
rect 342804 30662 342820 30718
rect 104060 30646 342820 30662
rect 73596 30538 339460 30554
rect 73596 30482 73612 30538
rect 73668 30482 339388 30538
rect 339444 30482 339460 30538
rect 73596 30466 339460 30482
rect 70012 30358 73124 30374
rect 70012 30302 70028 30358
rect 70084 30302 73052 30358
rect 73108 30302 73124 30358
rect 70012 30286 73124 30302
rect 92188 30358 494020 30374
rect 92188 30302 92204 30358
rect 92260 30302 493948 30358
rect 494004 30302 494020 30358
rect 92188 30286 494020 30302
rect 52540 29278 142900 29294
rect 52540 29222 52556 29278
rect 52612 29222 142828 29278
rect 142884 29222 142900 29278
rect 52540 29206 142900 29222
rect 53436 29098 164740 29114
rect 53436 29042 53452 29098
rect 53508 29042 164668 29098
rect 164724 29042 164740 29098
rect 53436 29026 164740 29042
rect 83676 28918 428500 28934
rect 83676 28862 83692 28918
rect 83748 28862 428428 28918
rect 428484 28862 428500 28918
rect 83676 28846 428500 28862
rect 87820 28738 90820 28754
rect 87820 28682 87836 28738
rect 87892 28682 90748 28738
rect 90804 28682 90820 28738
rect 87820 28666 90820 28682
rect 92076 28738 501412 28754
rect 92076 28682 92092 28738
rect 92148 28682 501340 28738
rect 501396 28682 501412 28738
rect 92076 28666 501412 28682
rect -1916 28350 597980 28446
rect -1916 28294 -1820 28350
rect -1764 28294 -1696 28350
rect -1640 28294 -1572 28350
rect -1516 28294 -1448 28350
rect -1392 28294 9234 28350
rect 9290 28294 9358 28350
rect 9414 28294 9482 28350
rect 9538 28294 9606 28350
rect 9662 28294 31878 28350
rect 31934 28294 32002 28350
rect 32058 28294 39954 28350
rect 40010 28294 40078 28350
rect 40134 28294 40202 28350
rect 40258 28294 40326 28350
rect 40382 28294 62598 28350
rect 62654 28294 62722 28350
rect 62778 28294 70674 28350
rect 70730 28294 70798 28350
rect 70854 28294 70922 28350
rect 70978 28294 71046 28350
rect 71102 28294 93318 28350
rect 93374 28294 93442 28350
rect 93498 28294 101394 28350
rect 101450 28294 101518 28350
rect 101574 28294 101642 28350
rect 101698 28294 101766 28350
rect 101822 28294 132114 28350
rect 132170 28294 132238 28350
rect 132294 28294 132362 28350
rect 132418 28294 132486 28350
rect 132542 28294 162834 28350
rect 162890 28294 162958 28350
rect 163014 28294 163082 28350
rect 163138 28294 163206 28350
rect 163262 28294 193554 28350
rect 193610 28294 193678 28350
rect 193734 28294 193802 28350
rect 193858 28294 193926 28350
rect 193982 28294 224274 28350
rect 224330 28294 224398 28350
rect 224454 28294 224522 28350
rect 224578 28294 224646 28350
rect 224702 28294 254994 28350
rect 255050 28294 255118 28350
rect 255174 28294 255242 28350
rect 255298 28294 255366 28350
rect 255422 28294 285714 28350
rect 285770 28294 285838 28350
rect 285894 28294 285962 28350
rect 286018 28294 286086 28350
rect 286142 28294 316434 28350
rect 316490 28294 316558 28350
rect 316614 28294 316682 28350
rect 316738 28294 316806 28350
rect 316862 28294 347154 28350
rect 347210 28294 347278 28350
rect 347334 28294 347402 28350
rect 347458 28294 347526 28350
rect 347582 28294 377874 28350
rect 377930 28294 377998 28350
rect 378054 28294 378122 28350
rect 378178 28294 378246 28350
rect 378302 28294 408594 28350
rect 408650 28294 408718 28350
rect 408774 28294 408842 28350
rect 408898 28294 408966 28350
rect 409022 28294 439314 28350
rect 439370 28294 439438 28350
rect 439494 28294 439562 28350
rect 439618 28294 439686 28350
rect 439742 28294 470034 28350
rect 470090 28294 470158 28350
rect 470214 28294 470282 28350
rect 470338 28294 470406 28350
rect 470462 28294 500754 28350
rect 500810 28294 500878 28350
rect 500934 28294 501002 28350
rect 501058 28294 501126 28350
rect 501182 28294 531474 28350
rect 531530 28294 531598 28350
rect 531654 28294 531722 28350
rect 531778 28294 531846 28350
rect 531902 28294 562194 28350
rect 562250 28294 562318 28350
rect 562374 28294 562442 28350
rect 562498 28294 562566 28350
rect 562622 28294 592914 28350
rect 592970 28294 593038 28350
rect 593094 28294 593162 28350
rect 593218 28294 593286 28350
rect 593342 28294 597456 28350
rect 597512 28294 597580 28350
rect 597636 28294 597704 28350
rect 597760 28294 597828 28350
rect 597884 28294 597980 28350
rect -1916 28226 597980 28294
rect -1916 28170 -1820 28226
rect -1764 28170 -1696 28226
rect -1640 28170 -1572 28226
rect -1516 28170 -1448 28226
rect -1392 28170 9234 28226
rect 9290 28170 9358 28226
rect 9414 28170 9482 28226
rect 9538 28170 9606 28226
rect 9662 28170 31878 28226
rect 31934 28170 32002 28226
rect 32058 28170 39954 28226
rect 40010 28170 40078 28226
rect 40134 28170 40202 28226
rect 40258 28170 40326 28226
rect 40382 28170 62598 28226
rect 62654 28170 62722 28226
rect 62778 28170 70674 28226
rect 70730 28170 70798 28226
rect 70854 28170 70922 28226
rect 70978 28170 71046 28226
rect 71102 28170 93318 28226
rect 93374 28170 93442 28226
rect 93498 28170 101394 28226
rect 101450 28170 101518 28226
rect 101574 28170 101642 28226
rect 101698 28170 101766 28226
rect 101822 28170 132114 28226
rect 132170 28170 132238 28226
rect 132294 28170 132362 28226
rect 132418 28170 132486 28226
rect 132542 28170 162834 28226
rect 162890 28170 162958 28226
rect 163014 28170 163082 28226
rect 163138 28170 163206 28226
rect 163262 28170 193554 28226
rect 193610 28170 193678 28226
rect 193734 28170 193802 28226
rect 193858 28170 193926 28226
rect 193982 28170 224274 28226
rect 224330 28170 224398 28226
rect 224454 28170 224522 28226
rect 224578 28170 224646 28226
rect 224702 28170 254994 28226
rect 255050 28170 255118 28226
rect 255174 28170 255242 28226
rect 255298 28170 255366 28226
rect 255422 28170 285714 28226
rect 285770 28170 285838 28226
rect 285894 28170 285962 28226
rect 286018 28170 286086 28226
rect 286142 28170 316434 28226
rect 316490 28170 316558 28226
rect 316614 28170 316682 28226
rect 316738 28170 316806 28226
rect 316862 28170 347154 28226
rect 347210 28170 347278 28226
rect 347334 28170 347402 28226
rect 347458 28170 347526 28226
rect 347582 28170 377874 28226
rect 377930 28170 377998 28226
rect 378054 28170 378122 28226
rect 378178 28170 378246 28226
rect 378302 28170 408594 28226
rect 408650 28170 408718 28226
rect 408774 28170 408842 28226
rect 408898 28170 408966 28226
rect 409022 28170 439314 28226
rect 439370 28170 439438 28226
rect 439494 28170 439562 28226
rect 439618 28170 439686 28226
rect 439742 28170 470034 28226
rect 470090 28170 470158 28226
rect 470214 28170 470282 28226
rect 470338 28170 470406 28226
rect 470462 28170 500754 28226
rect 500810 28170 500878 28226
rect 500934 28170 501002 28226
rect 501058 28170 501126 28226
rect 501182 28170 531474 28226
rect 531530 28170 531598 28226
rect 531654 28170 531722 28226
rect 531778 28170 531846 28226
rect 531902 28170 562194 28226
rect 562250 28170 562318 28226
rect 562374 28170 562442 28226
rect 562498 28170 562566 28226
rect 562622 28170 592914 28226
rect 592970 28170 593038 28226
rect 593094 28170 593162 28226
rect 593218 28170 593286 28226
rect 593342 28170 597456 28226
rect 597512 28170 597580 28226
rect 597636 28170 597704 28226
rect 597760 28170 597828 28226
rect 597884 28170 597980 28226
rect -1916 28102 597980 28170
rect -1916 28046 -1820 28102
rect -1764 28046 -1696 28102
rect -1640 28046 -1572 28102
rect -1516 28046 -1448 28102
rect -1392 28046 9234 28102
rect 9290 28046 9358 28102
rect 9414 28046 9482 28102
rect 9538 28046 9606 28102
rect 9662 28046 31878 28102
rect 31934 28046 32002 28102
rect 32058 28046 39954 28102
rect 40010 28046 40078 28102
rect 40134 28046 40202 28102
rect 40258 28046 40326 28102
rect 40382 28046 62598 28102
rect 62654 28046 62722 28102
rect 62778 28046 70674 28102
rect 70730 28046 70798 28102
rect 70854 28046 70922 28102
rect 70978 28046 71046 28102
rect 71102 28046 93318 28102
rect 93374 28046 93442 28102
rect 93498 28046 101394 28102
rect 101450 28046 101518 28102
rect 101574 28046 101642 28102
rect 101698 28046 101766 28102
rect 101822 28046 132114 28102
rect 132170 28046 132238 28102
rect 132294 28046 132362 28102
rect 132418 28046 132486 28102
rect 132542 28046 162834 28102
rect 162890 28046 162958 28102
rect 163014 28046 163082 28102
rect 163138 28046 163206 28102
rect 163262 28046 193554 28102
rect 193610 28046 193678 28102
rect 193734 28046 193802 28102
rect 193858 28046 193926 28102
rect 193982 28046 224274 28102
rect 224330 28046 224398 28102
rect 224454 28046 224522 28102
rect 224578 28046 224646 28102
rect 224702 28046 254994 28102
rect 255050 28046 255118 28102
rect 255174 28046 255242 28102
rect 255298 28046 255366 28102
rect 255422 28046 285714 28102
rect 285770 28046 285838 28102
rect 285894 28046 285962 28102
rect 286018 28046 286086 28102
rect 286142 28046 316434 28102
rect 316490 28046 316558 28102
rect 316614 28046 316682 28102
rect 316738 28046 316806 28102
rect 316862 28046 347154 28102
rect 347210 28046 347278 28102
rect 347334 28046 347402 28102
rect 347458 28046 347526 28102
rect 347582 28046 377874 28102
rect 377930 28046 377998 28102
rect 378054 28046 378122 28102
rect 378178 28046 378246 28102
rect 378302 28046 408594 28102
rect 408650 28046 408718 28102
rect 408774 28046 408842 28102
rect 408898 28046 408966 28102
rect 409022 28046 439314 28102
rect 439370 28046 439438 28102
rect 439494 28046 439562 28102
rect 439618 28046 439686 28102
rect 439742 28046 470034 28102
rect 470090 28046 470158 28102
rect 470214 28046 470282 28102
rect 470338 28046 470406 28102
rect 470462 28046 500754 28102
rect 500810 28046 500878 28102
rect 500934 28046 501002 28102
rect 501058 28046 501126 28102
rect 501182 28046 531474 28102
rect 531530 28046 531598 28102
rect 531654 28046 531722 28102
rect 531778 28046 531846 28102
rect 531902 28046 562194 28102
rect 562250 28046 562318 28102
rect 562374 28046 562442 28102
rect 562498 28046 562566 28102
rect 562622 28046 592914 28102
rect 592970 28046 593038 28102
rect 593094 28046 593162 28102
rect 593218 28046 593286 28102
rect 593342 28046 597456 28102
rect 597512 28046 597580 28102
rect 597636 28046 597704 28102
rect 597760 28046 597828 28102
rect 597884 28046 597980 28102
rect -1916 27978 597980 28046
rect -1916 27922 -1820 27978
rect -1764 27922 -1696 27978
rect -1640 27922 -1572 27978
rect -1516 27922 -1448 27978
rect -1392 27922 9234 27978
rect 9290 27922 9358 27978
rect 9414 27922 9482 27978
rect 9538 27922 9606 27978
rect 9662 27922 31878 27978
rect 31934 27922 32002 27978
rect 32058 27922 39954 27978
rect 40010 27922 40078 27978
rect 40134 27922 40202 27978
rect 40258 27922 40326 27978
rect 40382 27922 62598 27978
rect 62654 27922 62722 27978
rect 62778 27922 70674 27978
rect 70730 27922 70798 27978
rect 70854 27922 70922 27978
rect 70978 27922 71046 27978
rect 71102 27922 93318 27978
rect 93374 27922 93442 27978
rect 93498 27922 101394 27978
rect 101450 27922 101518 27978
rect 101574 27922 101642 27978
rect 101698 27922 101766 27978
rect 101822 27922 132114 27978
rect 132170 27922 132238 27978
rect 132294 27922 132362 27978
rect 132418 27922 132486 27978
rect 132542 27922 162834 27978
rect 162890 27922 162958 27978
rect 163014 27922 163082 27978
rect 163138 27922 163206 27978
rect 163262 27922 193554 27978
rect 193610 27922 193678 27978
rect 193734 27922 193802 27978
rect 193858 27922 193926 27978
rect 193982 27922 224274 27978
rect 224330 27922 224398 27978
rect 224454 27922 224522 27978
rect 224578 27922 224646 27978
rect 224702 27922 254994 27978
rect 255050 27922 255118 27978
rect 255174 27922 255242 27978
rect 255298 27922 255366 27978
rect 255422 27922 285714 27978
rect 285770 27922 285838 27978
rect 285894 27922 285962 27978
rect 286018 27922 286086 27978
rect 286142 27922 316434 27978
rect 316490 27922 316558 27978
rect 316614 27922 316682 27978
rect 316738 27922 316806 27978
rect 316862 27922 347154 27978
rect 347210 27922 347278 27978
rect 347334 27922 347402 27978
rect 347458 27922 347526 27978
rect 347582 27922 377874 27978
rect 377930 27922 377998 27978
rect 378054 27922 378122 27978
rect 378178 27922 378246 27978
rect 378302 27922 408594 27978
rect 408650 27922 408718 27978
rect 408774 27922 408842 27978
rect 408898 27922 408966 27978
rect 409022 27922 439314 27978
rect 439370 27922 439438 27978
rect 439494 27922 439562 27978
rect 439618 27922 439686 27978
rect 439742 27922 470034 27978
rect 470090 27922 470158 27978
rect 470214 27922 470282 27978
rect 470338 27922 470406 27978
rect 470462 27922 500754 27978
rect 500810 27922 500878 27978
rect 500934 27922 501002 27978
rect 501058 27922 501126 27978
rect 501182 27922 531474 27978
rect 531530 27922 531598 27978
rect 531654 27922 531722 27978
rect 531778 27922 531846 27978
rect 531902 27922 562194 27978
rect 562250 27922 562318 27978
rect 562374 27922 562442 27978
rect 562498 27922 562566 27978
rect 562622 27922 592914 27978
rect 592970 27922 593038 27978
rect 593094 27922 593162 27978
rect 593218 27922 593286 27978
rect 593342 27922 597456 27978
rect 597512 27922 597580 27978
rect 597636 27922 597704 27978
rect 597760 27922 597828 27978
rect 597884 27922 597980 27978
rect -1916 27826 597980 27922
rect 73036 26938 173140 26954
rect 73036 26882 73052 26938
rect 73108 26882 173068 26938
rect 173124 26882 173140 26938
rect 73036 26866 173140 26882
rect 66204 26218 73236 26234
rect 66204 26162 66220 26218
rect 66276 26162 73164 26218
rect 73220 26162 73236 26218
rect 66204 26146 73236 26162
rect 80540 26218 83316 26234
rect 80540 26162 80556 26218
rect 80612 26162 83244 26218
rect 83300 26162 83316 26218
rect 80540 26146 83316 26162
rect 73484 26038 104148 26054
rect 73484 25982 73500 26038
rect 73556 25982 104076 26038
rect 104132 25982 104148 26038
rect 73484 25966 104148 25982
rect 61276 25858 236980 25874
rect 61276 25802 61292 25858
rect 61348 25802 236908 25858
rect 236964 25802 236980 25858
rect 61276 25786 236980 25802
rect 89836 25678 371380 25694
rect 89836 25622 89852 25678
rect 89908 25622 371308 25678
rect 371364 25622 371380 25678
rect 89836 25606 371380 25622
rect 85020 25498 87908 25514
rect 85020 25442 85036 25498
rect 85092 25442 87836 25498
rect 87892 25442 87908 25498
rect 85020 25426 87908 25442
rect 93868 25498 460420 25514
rect 93868 25442 93884 25498
rect 93940 25442 460348 25498
rect 460404 25442 460420 25498
rect 93868 25426 460420 25442
rect 46492 25318 107620 25334
rect 46492 25262 46508 25318
rect 46564 25262 107548 25318
rect 107604 25262 107620 25318
rect 46492 25246 107620 25262
rect 108316 25318 574660 25334
rect 108316 25262 108332 25318
rect 108388 25262 574588 25318
rect 574644 25262 574660 25318
rect 108316 25246 574660 25262
rect 71916 25138 76708 25154
rect 71916 25082 71932 25138
rect 71988 25082 76636 25138
rect 76692 25082 76708 25138
rect 71916 25066 76708 25082
rect 77628 25138 80068 25154
rect 77628 25082 77644 25138
rect 77700 25082 79996 25138
rect 80052 25082 80068 25138
rect 77628 25066 80068 25082
rect 53324 24598 73124 24614
rect 53324 24542 53340 24598
rect 53396 24542 73052 24598
rect 73108 24542 73124 24598
rect 53324 24526 73124 24542
rect 50300 24418 144580 24434
rect 50300 24362 50316 24418
rect 50372 24362 144508 24418
rect 144564 24362 144580 24418
rect 50300 24346 144580 24362
rect 51868 24238 152980 24254
rect 51868 24182 51884 24238
rect 51940 24182 152908 24238
rect 152964 24182 152980 24238
rect 51868 24166 152980 24182
rect 76844 24058 347860 24074
rect 76844 24002 76860 24058
rect 76916 24002 347788 24058
rect 347844 24002 347860 24058
rect 76844 23986 347860 24002
rect 80428 23878 388180 23894
rect 80428 23822 80444 23878
rect 80500 23822 388108 23878
rect 388164 23822 388180 23878
rect 80428 23806 388180 23822
rect 81660 23698 391540 23714
rect 81660 23642 81676 23698
rect 81732 23642 391468 23698
rect 391524 23642 391540 23698
rect 81660 23626 391540 23642
rect 69900 22798 314260 22814
rect 69900 22742 69916 22798
rect 69972 22742 314188 22798
rect 314244 22742 314260 22798
rect 69900 22726 314260 22742
rect 86924 22618 450340 22634
rect 86924 22562 86940 22618
rect 86996 22562 450268 22618
rect 450324 22562 450340 22618
rect 86924 22546 450340 22562
rect -1916 22350 597980 22446
rect -1916 22294 -860 22350
rect -804 22294 -736 22350
rect -680 22294 -612 22350
rect -556 22294 -488 22350
rect -432 22294 5514 22350
rect 5570 22294 5638 22350
rect 5694 22294 5762 22350
rect 5818 22294 5886 22350
rect 5942 22294 16518 22350
rect 16574 22294 16642 22350
rect 16698 22294 36234 22350
rect 36290 22294 36358 22350
rect 36414 22294 36482 22350
rect 36538 22294 36606 22350
rect 36662 22294 47238 22350
rect 47294 22294 47362 22350
rect 47418 22294 66954 22350
rect 67010 22294 67078 22350
rect 67134 22294 67202 22350
rect 67258 22294 67326 22350
rect 67382 22294 77958 22350
rect 78014 22294 78082 22350
rect 78138 22294 97674 22350
rect 97730 22294 97798 22350
rect 97854 22294 97922 22350
rect 97978 22294 98046 22350
rect 98102 22294 108678 22350
rect 108734 22294 108802 22350
rect 108858 22294 128394 22350
rect 128450 22294 128518 22350
rect 128574 22294 128642 22350
rect 128698 22294 128766 22350
rect 128822 22294 159114 22350
rect 159170 22294 159238 22350
rect 159294 22294 159362 22350
rect 159418 22294 159486 22350
rect 159542 22294 189834 22350
rect 189890 22294 189958 22350
rect 190014 22294 190082 22350
rect 190138 22294 190206 22350
rect 190262 22294 220554 22350
rect 220610 22294 220678 22350
rect 220734 22294 220802 22350
rect 220858 22294 220926 22350
rect 220982 22294 251274 22350
rect 251330 22294 251398 22350
rect 251454 22294 251522 22350
rect 251578 22294 251646 22350
rect 251702 22294 281994 22350
rect 282050 22294 282118 22350
rect 282174 22294 282242 22350
rect 282298 22294 282366 22350
rect 282422 22294 312714 22350
rect 312770 22294 312838 22350
rect 312894 22294 312962 22350
rect 313018 22294 313086 22350
rect 313142 22294 343434 22350
rect 343490 22294 343558 22350
rect 343614 22294 343682 22350
rect 343738 22294 343806 22350
rect 343862 22294 374154 22350
rect 374210 22294 374278 22350
rect 374334 22294 374402 22350
rect 374458 22294 374526 22350
rect 374582 22294 404874 22350
rect 404930 22294 404998 22350
rect 405054 22294 405122 22350
rect 405178 22294 405246 22350
rect 405302 22294 435594 22350
rect 435650 22294 435718 22350
rect 435774 22294 435842 22350
rect 435898 22294 435966 22350
rect 436022 22294 466314 22350
rect 466370 22294 466438 22350
rect 466494 22294 466562 22350
rect 466618 22294 466686 22350
rect 466742 22294 497034 22350
rect 497090 22294 497158 22350
rect 497214 22294 497282 22350
rect 497338 22294 497406 22350
rect 497462 22294 527754 22350
rect 527810 22294 527878 22350
rect 527934 22294 528002 22350
rect 528058 22294 528126 22350
rect 528182 22294 558474 22350
rect 558530 22294 558598 22350
rect 558654 22294 558722 22350
rect 558778 22294 558846 22350
rect 558902 22294 589194 22350
rect 589250 22294 589318 22350
rect 589374 22294 589442 22350
rect 589498 22294 589566 22350
rect 589622 22294 596496 22350
rect 596552 22294 596620 22350
rect 596676 22294 596744 22350
rect 596800 22294 596868 22350
rect 596924 22294 597980 22350
rect -1916 22226 597980 22294
rect -1916 22170 -860 22226
rect -804 22170 -736 22226
rect -680 22170 -612 22226
rect -556 22170 -488 22226
rect -432 22170 5514 22226
rect 5570 22170 5638 22226
rect 5694 22170 5762 22226
rect 5818 22170 5886 22226
rect 5942 22170 16518 22226
rect 16574 22170 16642 22226
rect 16698 22170 36234 22226
rect 36290 22170 36358 22226
rect 36414 22170 36482 22226
rect 36538 22170 36606 22226
rect 36662 22170 47238 22226
rect 47294 22170 47362 22226
rect 47418 22170 66954 22226
rect 67010 22170 67078 22226
rect 67134 22170 67202 22226
rect 67258 22170 67326 22226
rect 67382 22170 77958 22226
rect 78014 22170 78082 22226
rect 78138 22170 97674 22226
rect 97730 22170 97798 22226
rect 97854 22170 97922 22226
rect 97978 22170 98046 22226
rect 98102 22170 108678 22226
rect 108734 22170 108802 22226
rect 108858 22170 128394 22226
rect 128450 22170 128518 22226
rect 128574 22170 128642 22226
rect 128698 22170 128766 22226
rect 128822 22170 159114 22226
rect 159170 22170 159238 22226
rect 159294 22170 159362 22226
rect 159418 22170 159486 22226
rect 159542 22170 189834 22226
rect 189890 22170 189958 22226
rect 190014 22170 190082 22226
rect 190138 22170 190206 22226
rect 190262 22170 220554 22226
rect 220610 22170 220678 22226
rect 220734 22170 220802 22226
rect 220858 22170 220926 22226
rect 220982 22170 251274 22226
rect 251330 22170 251398 22226
rect 251454 22170 251522 22226
rect 251578 22170 251646 22226
rect 251702 22170 281994 22226
rect 282050 22170 282118 22226
rect 282174 22170 282242 22226
rect 282298 22170 282366 22226
rect 282422 22170 312714 22226
rect 312770 22170 312838 22226
rect 312894 22170 312962 22226
rect 313018 22170 313086 22226
rect 313142 22170 343434 22226
rect 343490 22170 343558 22226
rect 343614 22170 343682 22226
rect 343738 22170 343806 22226
rect 343862 22170 374154 22226
rect 374210 22170 374278 22226
rect 374334 22170 374402 22226
rect 374458 22170 374526 22226
rect 374582 22170 404874 22226
rect 404930 22170 404998 22226
rect 405054 22170 405122 22226
rect 405178 22170 405246 22226
rect 405302 22170 435594 22226
rect 435650 22170 435718 22226
rect 435774 22170 435842 22226
rect 435898 22170 435966 22226
rect 436022 22170 466314 22226
rect 466370 22170 466438 22226
rect 466494 22170 466562 22226
rect 466618 22170 466686 22226
rect 466742 22170 497034 22226
rect 497090 22170 497158 22226
rect 497214 22170 497282 22226
rect 497338 22170 497406 22226
rect 497462 22170 527754 22226
rect 527810 22170 527878 22226
rect 527934 22170 528002 22226
rect 528058 22170 528126 22226
rect 528182 22170 558474 22226
rect 558530 22170 558598 22226
rect 558654 22170 558722 22226
rect 558778 22170 558846 22226
rect 558902 22170 589194 22226
rect 589250 22170 589318 22226
rect 589374 22170 589442 22226
rect 589498 22170 589566 22226
rect 589622 22170 596496 22226
rect 596552 22170 596620 22226
rect 596676 22170 596744 22226
rect 596800 22170 596868 22226
rect 596924 22170 597980 22226
rect -1916 22102 597980 22170
rect -1916 22046 -860 22102
rect -804 22046 -736 22102
rect -680 22046 -612 22102
rect -556 22046 -488 22102
rect -432 22046 5514 22102
rect 5570 22046 5638 22102
rect 5694 22046 5762 22102
rect 5818 22046 5886 22102
rect 5942 22046 16518 22102
rect 16574 22046 16642 22102
rect 16698 22046 36234 22102
rect 36290 22046 36358 22102
rect 36414 22046 36482 22102
rect 36538 22046 36606 22102
rect 36662 22046 47238 22102
rect 47294 22046 47362 22102
rect 47418 22046 66954 22102
rect 67010 22046 67078 22102
rect 67134 22046 67202 22102
rect 67258 22046 67326 22102
rect 67382 22046 77958 22102
rect 78014 22046 78082 22102
rect 78138 22046 97674 22102
rect 97730 22046 97798 22102
rect 97854 22046 97922 22102
rect 97978 22046 98046 22102
rect 98102 22046 108678 22102
rect 108734 22046 108802 22102
rect 108858 22046 128394 22102
rect 128450 22046 128518 22102
rect 128574 22046 128642 22102
rect 128698 22046 128766 22102
rect 128822 22046 159114 22102
rect 159170 22046 159238 22102
rect 159294 22046 159362 22102
rect 159418 22046 159486 22102
rect 159542 22046 189834 22102
rect 189890 22046 189958 22102
rect 190014 22046 190082 22102
rect 190138 22046 190206 22102
rect 190262 22046 220554 22102
rect 220610 22046 220678 22102
rect 220734 22046 220802 22102
rect 220858 22046 220926 22102
rect 220982 22046 251274 22102
rect 251330 22046 251398 22102
rect 251454 22046 251522 22102
rect 251578 22046 251646 22102
rect 251702 22046 281994 22102
rect 282050 22046 282118 22102
rect 282174 22046 282242 22102
rect 282298 22046 282366 22102
rect 282422 22046 312714 22102
rect 312770 22046 312838 22102
rect 312894 22046 312962 22102
rect 313018 22046 313086 22102
rect 313142 22046 343434 22102
rect 343490 22046 343558 22102
rect 343614 22046 343682 22102
rect 343738 22046 343806 22102
rect 343862 22046 374154 22102
rect 374210 22046 374278 22102
rect 374334 22046 374402 22102
rect 374458 22046 374526 22102
rect 374582 22046 404874 22102
rect 404930 22046 404998 22102
rect 405054 22046 405122 22102
rect 405178 22046 405246 22102
rect 405302 22046 435594 22102
rect 435650 22046 435718 22102
rect 435774 22046 435842 22102
rect 435898 22046 435966 22102
rect 436022 22046 466314 22102
rect 466370 22046 466438 22102
rect 466494 22046 466562 22102
rect 466618 22046 466686 22102
rect 466742 22046 497034 22102
rect 497090 22046 497158 22102
rect 497214 22046 497282 22102
rect 497338 22046 497406 22102
rect 497462 22046 527754 22102
rect 527810 22046 527878 22102
rect 527934 22046 528002 22102
rect 528058 22046 528126 22102
rect 528182 22046 558474 22102
rect 558530 22046 558598 22102
rect 558654 22046 558722 22102
rect 558778 22046 558846 22102
rect 558902 22046 589194 22102
rect 589250 22046 589318 22102
rect 589374 22046 589442 22102
rect 589498 22046 589566 22102
rect 589622 22046 596496 22102
rect 596552 22046 596620 22102
rect 596676 22046 596744 22102
rect 596800 22046 596868 22102
rect 596924 22046 597980 22102
rect -1916 21978 597980 22046
rect -1916 21922 -860 21978
rect -804 21922 -736 21978
rect -680 21922 -612 21978
rect -556 21922 -488 21978
rect -432 21922 5514 21978
rect 5570 21922 5638 21978
rect 5694 21922 5762 21978
rect 5818 21922 5886 21978
rect 5942 21922 16518 21978
rect 16574 21922 16642 21978
rect 16698 21922 36234 21978
rect 36290 21922 36358 21978
rect 36414 21922 36482 21978
rect 36538 21922 36606 21978
rect 36662 21922 47238 21978
rect 47294 21922 47362 21978
rect 47418 21922 66954 21978
rect 67010 21922 67078 21978
rect 67134 21922 67202 21978
rect 67258 21922 67326 21978
rect 67382 21922 77958 21978
rect 78014 21922 78082 21978
rect 78138 21922 97674 21978
rect 97730 21922 97798 21978
rect 97854 21922 97922 21978
rect 97978 21922 98046 21978
rect 98102 21922 108678 21978
rect 108734 21922 108802 21978
rect 108858 21922 128394 21978
rect 128450 21922 128518 21978
rect 128574 21922 128642 21978
rect 128698 21922 128766 21978
rect 128822 21922 159114 21978
rect 159170 21922 159238 21978
rect 159294 21922 159362 21978
rect 159418 21922 159486 21978
rect 159542 21922 189834 21978
rect 189890 21922 189958 21978
rect 190014 21922 190082 21978
rect 190138 21922 190206 21978
rect 190262 21922 220554 21978
rect 220610 21922 220678 21978
rect 220734 21922 220802 21978
rect 220858 21922 220926 21978
rect 220982 21922 251274 21978
rect 251330 21922 251398 21978
rect 251454 21922 251522 21978
rect 251578 21922 251646 21978
rect 251702 21922 281994 21978
rect 282050 21922 282118 21978
rect 282174 21922 282242 21978
rect 282298 21922 282366 21978
rect 282422 21922 312714 21978
rect 312770 21922 312838 21978
rect 312894 21922 312962 21978
rect 313018 21922 313086 21978
rect 313142 21922 343434 21978
rect 343490 21922 343558 21978
rect 343614 21922 343682 21978
rect 343738 21922 343806 21978
rect 343862 21922 374154 21978
rect 374210 21922 374278 21978
rect 374334 21922 374402 21978
rect 374458 21922 374526 21978
rect 374582 21922 404874 21978
rect 404930 21922 404998 21978
rect 405054 21922 405122 21978
rect 405178 21922 405246 21978
rect 405302 21922 435594 21978
rect 435650 21922 435718 21978
rect 435774 21922 435842 21978
rect 435898 21922 435966 21978
rect 436022 21922 466314 21978
rect 466370 21922 466438 21978
rect 466494 21922 466562 21978
rect 466618 21922 466686 21978
rect 466742 21922 497034 21978
rect 497090 21922 497158 21978
rect 497214 21922 497282 21978
rect 497338 21922 497406 21978
rect 497462 21922 527754 21978
rect 527810 21922 527878 21978
rect 527934 21922 528002 21978
rect 528058 21922 528126 21978
rect 528182 21922 558474 21978
rect 558530 21922 558598 21978
rect 558654 21922 558722 21978
rect 558778 21922 558846 21978
rect 558902 21922 589194 21978
rect 589250 21922 589318 21978
rect 589374 21922 589442 21978
rect 589498 21922 589566 21978
rect 589622 21922 596496 21978
rect 596552 21922 596620 21978
rect 596676 21922 596744 21978
rect 596800 21922 596868 21978
rect 596924 21922 597980 21978
rect -1916 21826 597980 21922
rect 76956 21718 78388 21734
rect 76956 21662 76972 21718
rect 77028 21662 78316 21718
rect 78372 21662 78388 21718
rect 76956 21646 78388 21662
rect 102380 20998 108404 21014
rect 102380 20942 102396 20998
rect 102452 20942 108332 20998
rect 108388 20942 108404 20998
rect 102380 20926 108404 20942
rect 53884 20638 174820 20654
rect 53884 20582 53900 20638
rect 53956 20582 174748 20638
rect 174804 20582 174820 20638
rect 53884 20566 174820 20582
rect 55452 20458 194980 20474
rect 55452 20402 55468 20458
rect 55524 20402 194908 20458
rect 194964 20402 194980 20458
rect 55452 20386 194980 20402
rect 78636 20278 359620 20294
rect 78636 20222 78652 20278
rect 78708 20222 359548 20278
rect 359604 20222 359620 20278
rect 78636 20206 359620 20222
rect 76732 19378 89924 19394
rect 76732 19322 76748 19378
rect 76804 19322 89852 19378
rect 89908 19322 89924 19378
rect 76732 19306 89924 19322
rect 98796 19378 100004 19394
rect 98796 19322 98812 19378
rect 98868 19322 99932 19378
rect 99988 19322 100004 19378
rect 98796 19306 100004 19322
rect 50188 19198 137860 19214
rect 50188 19142 50204 19198
rect 50260 19142 137788 19198
rect 137844 19142 137860 19198
rect 50188 19126 137860 19142
rect 51756 19018 158020 19034
rect 51756 18962 51772 19018
rect 51828 18962 157948 19018
rect 158004 18962 158020 19018
rect 51756 18946 158020 18962
rect 56684 18838 191620 18854
rect 56684 18782 56700 18838
rect 56756 18782 191548 18838
rect 191604 18782 191620 18838
rect 56684 18766 191620 18782
rect 63404 18658 245604 18674
rect 63404 18602 63420 18658
rect 63476 18602 245532 18658
rect 245588 18602 245604 18658
rect 63404 18586 245604 18602
rect 50972 17578 149620 17594
rect 50972 17522 50988 17578
rect 51044 17522 149548 17578
rect 149604 17522 149620 17578
rect 50972 17506 149620 17522
rect 55228 17398 183220 17414
rect 55228 17342 55244 17398
rect 55300 17342 183148 17398
rect 183204 17342 183220 17398
rect 55228 17326 183220 17342
rect 73148 17218 336100 17234
rect 73148 17162 73164 17218
rect 73220 17162 336028 17218
rect 336084 17162 336100 17218
rect 73148 17146 336100 17162
rect 89836 17038 410020 17054
rect 89836 16982 89852 17038
rect 89908 16982 409948 17038
rect 410004 16982 410020 17038
rect 89836 16966 410020 16982
rect 42460 16858 87572 16874
rect 42460 16802 42476 16858
rect 42532 16802 87500 16858
rect 87556 16802 87572 16858
rect 42460 16786 87572 16802
rect 93756 16858 504100 16874
rect 93756 16802 93772 16858
rect 93828 16802 504028 16858
rect 504084 16802 504100 16858
rect 93756 16786 504100 16802
rect 50524 15958 146260 15974
rect 50524 15902 50540 15958
rect 50596 15902 146188 15958
rect 146244 15902 146260 15958
rect 50524 15886 146260 15902
rect 56908 15778 201812 15794
rect 56908 15722 56924 15778
rect 56980 15722 201740 15778
rect 201796 15722 201812 15778
rect 56908 15706 201812 15722
rect 64188 15598 262180 15614
rect 64188 15542 64204 15598
rect 64260 15542 262108 15598
rect 262164 15542 262180 15598
rect 64188 15526 262180 15542
rect 78916 15346 95972 15434
rect 78916 15254 79004 15346
rect 44700 15238 79004 15254
rect 44700 15182 44716 15238
rect 44772 15182 79004 15238
rect 44700 15166 79004 15182
rect 93644 15238 94964 15254
rect 93644 15182 93660 15238
rect 93716 15182 94892 15238
rect 94948 15182 94964 15238
rect 93644 15166 94964 15182
rect 95884 15238 95972 15346
rect 95884 15182 95900 15238
rect 95956 15182 95972 15238
rect 95884 15166 95972 15182
rect 96108 15418 478900 15434
rect 96108 15362 478828 15418
rect 478884 15362 478900 15418
rect 96108 15346 478900 15362
rect 96108 15074 96196 15346
rect 97116 15238 531204 15254
rect 97116 15182 97132 15238
rect 97188 15182 531132 15238
rect 531188 15182 531204 15238
rect 97116 15166 531204 15182
rect 95324 15058 96196 15074
rect 95324 15002 95340 15058
rect 95396 15002 96196 15058
rect 95324 14986 96196 15002
rect 46828 14518 46916 14534
rect 46828 14462 46844 14518
rect 46900 14462 46916 14518
rect 46828 14174 46916 14462
rect 50076 14338 131364 14354
rect 50076 14282 50092 14338
rect 50148 14282 131292 14338
rect 131348 14282 131364 14338
rect 50076 14266 131364 14282
rect 46828 14158 47028 14174
rect 46828 14102 46956 14158
rect 47012 14102 47028 14158
rect 46828 14086 47028 14102
rect 52316 14158 161380 14174
rect 52316 14102 52332 14158
rect 52388 14102 161308 14158
rect 161364 14102 161380 14158
rect 52316 14086 161380 14102
rect 55340 13978 179860 13994
rect 55340 13922 55356 13978
rect 55412 13922 179788 13978
rect 179844 13922 179860 13978
rect 55340 13906 179860 13922
rect 63292 13798 250420 13814
rect 63292 13742 63308 13798
rect 63364 13742 250348 13798
rect 250404 13742 250420 13798
rect 63292 13726 250420 13742
rect 89052 13618 474084 13634
rect 89052 13562 89068 13618
rect 89124 13562 474012 13618
rect 474068 13562 474084 13618
rect 89052 13546 474084 13562
rect 56348 13438 66068 13454
rect 56348 13382 56364 13438
rect 56420 13382 65996 13438
rect 66052 13382 66068 13438
rect 56348 13366 66068 13382
rect 71580 13438 76484 13454
rect 71580 13382 71596 13438
rect 71652 13382 76412 13438
rect 76468 13382 76484 13438
rect 71580 13366 76484 13382
rect 49852 12538 139540 12554
rect 49852 12482 49868 12538
rect 49924 12482 139468 12538
rect 139524 12482 139540 12538
rect 49852 12466 139540 12482
rect 83228 12358 393220 12374
rect 83228 12302 83244 12358
rect 83300 12302 393148 12358
rect 393204 12302 393220 12358
rect 83228 12286 393220 12302
rect 79980 12178 394900 12194
rect 79980 12122 79996 12178
rect 80052 12122 394828 12178
rect 394884 12122 394900 12178
rect 79980 12106 394900 12122
rect 45596 11998 104260 12014
rect 45596 11942 45612 11998
rect 45668 11942 104188 11998
rect 104244 11942 104260 11998
rect 45596 11926 104260 11942
rect 111004 11998 438580 12014
rect 111004 11942 111020 11998
rect 111076 11942 438508 11998
rect 438564 11942 438580 11998
rect 111004 11926 438580 11942
rect 87820 11818 93956 11834
rect 87820 11762 87836 11818
rect 87892 11762 93884 11818
rect 93940 11762 93956 11818
rect 87820 11746 93956 11762
rect 103388 11818 495700 11834
rect 103388 11762 103404 11818
rect 103460 11762 495628 11818
rect 495684 11762 495700 11818
rect 103388 11746 495700 11762
rect 90956 11098 111092 11114
rect 90956 11042 90972 11098
rect 91028 11042 111020 11098
rect 111076 11042 111092 11098
rect 90956 11026 111092 11042
rect 57244 10918 203716 10934
rect 57244 10862 57260 10918
rect 57316 10862 203644 10918
rect 203700 10862 203716 10918
rect 57244 10846 203716 10862
rect 93084 10738 508356 10754
rect 93084 10682 93100 10738
rect 93156 10682 508284 10738
rect 508340 10682 508356 10738
rect 93084 10666 508356 10682
rect -1916 10350 597980 10446
rect -1916 10294 -1820 10350
rect -1764 10294 -1696 10350
rect -1640 10294 -1572 10350
rect -1516 10294 -1448 10350
rect -1392 10294 9234 10350
rect 9290 10294 9358 10350
rect 9414 10294 9482 10350
rect 9538 10294 9606 10350
rect 9662 10294 31878 10350
rect 31934 10294 32002 10350
rect 32058 10294 39954 10350
rect 40010 10294 40078 10350
rect 40134 10294 40202 10350
rect 40258 10294 40326 10350
rect 40382 10294 62598 10350
rect 62654 10294 62722 10350
rect 62778 10294 70674 10350
rect 70730 10294 70798 10350
rect 70854 10294 70922 10350
rect 70978 10294 71046 10350
rect 71102 10294 93318 10350
rect 93374 10294 93442 10350
rect 93498 10294 101394 10350
rect 101450 10294 101518 10350
rect 101574 10294 101642 10350
rect 101698 10294 101766 10350
rect 101822 10294 132114 10350
rect 132170 10294 132238 10350
rect 132294 10294 132362 10350
rect 132418 10294 132486 10350
rect 132542 10294 162834 10350
rect 162890 10294 162958 10350
rect 163014 10294 163082 10350
rect 163138 10294 163206 10350
rect 163262 10294 193554 10350
rect 193610 10294 193678 10350
rect 193734 10294 193802 10350
rect 193858 10294 193926 10350
rect 193982 10294 224274 10350
rect 224330 10294 224398 10350
rect 224454 10294 224522 10350
rect 224578 10294 224646 10350
rect 224702 10294 254994 10350
rect 255050 10294 255118 10350
rect 255174 10294 255242 10350
rect 255298 10294 255366 10350
rect 255422 10294 285714 10350
rect 285770 10294 285838 10350
rect 285894 10294 285962 10350
rect 286018 10294 286086 10350
rect 286142 10294 316434 10350
rect 316490 10294 316558 10350
rect 316614 10294 316682 10350
rect 316738 10294 316806 10350
rect 316862 10294 347154 10350
rect 347210 10294 347278 10350
rect 347334 10294 347402 10350
rect 347458 10294 347526 10350
rect 347582 10294 377874 10350
rect 377930 10294 377998 10350
rect 378054 10294 378122 10350
rect 378178 10294 378246 10350
rect 378302 10294 408594 10350
rect 408650 10294 408718 10350
rect 408774 10294 408842 10350
rect 408898 10294 408966 10350
rect 409022 10294 439314 10350
rect 439370 10294 439438 10350
rect 439494 10294 439562 10350
rect 439618 10294 439686 10350
rect 439742 10294 470034 10350
rect 470090 10294 470158 10350
rect 470214 10294 470282 10350
rect 470338 10294 470406 10350
rect 470462 10294 500754 10350
rect 500810 10294 500878 10350
rect 500934 10294 501002 10350
rect 501058 10294 501126 10350
rect 501182 10294 531474 10350
rect 531530 10294 531598 10350
rect 531654 10294 531722 10350
rect 531778 10294 531846 10350
rect 531902 10294 562194 10350
rect 562250 10294 562318 10350
rect 562374 10294 562442 10350
rect 562498 10294 562566 10350
rect 562622 10294 592914 10350
rect 592970 10294 593038 10350
rect 593094 10294 593162 10350
rect 593218 10294 593286 10350
rect 593342 10294 597456 10350
rect 597512 10294 597580 10350
rect 597636 10294 597704 10350
rect 597760 10294 597828 10350
rect 597884 10294 597980 10350
rect -1916 10226 597980 10294
rect -1916 10170 -1820 10226
rect -1764 10170 -1696 10226
rect -1640 10170 -1572 10226
rect -1516 10170 -1448 10226
rect -1392 10170 9234 10226
rect 9290 10170 9358 10226
rect 9414 10170 9482 10226
rect 9538 10170 9606 10226
rect 9662 10170 31878 10226
rect 31934 10170 32002 10226
rect 32058 10170 39954 10226
rect 40010 10170 40078 10226
rect 40134 10170 40202 10226
rect 40258 10170 40326 10226
rect 40382 10170 62598 10226
rect 62654 10170 62722 10226
rect 62778 10170 70674 10226
rect 70730 10170 70798 10226
rect 70854 10170 70922 10226
rect 70978 10170 71046 10226
rect 71102 10170 93318 10226
rect 93374 10170 93442 10226
rect 93498 10170 101394 10226
rect 101450 10170 101518 10226
rect 101574 10170 101642 10226
rect 101698 10170 101766 10226
rect 101822 10170 132114 10226
rect 132170 10170 132238 10226
rect 132294 10170 132362 10226
rect 132418 10170 132486 10226
rect 132542 10170 162834 10226
rect 162890 10170 162958 10226
rect 163014 10170 163082 10226
rect 163138 10170 163206 10226
rect 163262 10170 193554 10226
rect 193610 10170 193678 10226
rect 193734 10170 193802 10226
rect 193858 10170 193926 10226
rect 193982 10170 224274 10226
rect 224330 10170 224398 10226
rect 224454 10170 224522 10226
rect 224578 10170 224646 10226
rect 224702 10170 254994 10226
rect 255050 10170 255118 10226
rect 255174 10170 255242 10226
rect 255298 10170 255366 10226
rect 255422 10170 285714 10226
rect 285770 10170 285838 10226
rect 285894 10170 285962 10226
rect 286018 10170 286086 10226
rect 286142 10170 316434 10226
rect 316490 10170 316558 10226
rect 316614 10170 316682 10226
rect 316738 10170 316806 10226
rect 316862 10170 347154 10226
rect 347210 10170 347278 10226
rect 347334 10170 347402 10226
rect 347458 10170 347526 10226
rect 347582 10170 377874 10226
rect 377930 10170 377998 10226
rect 378054 10170 378122 10226
rect 378178 10170 378246 10226
rect 378302 10170 408594 10226
rect 408650 10170 408718 10226
rect 408774 10170 408842 10226
rect 408898 10170 408966 10226
rect 409022 10170 439314 10226
rect 439370 10170 439438 10226
rect 439494 10170 439562 10226
rect 439618 10170 439686 10226
rect 439742 10170 470034 10226
rect 470090 10170 470158 10226
rect 470214 10170 470282 10226
rect 470338 10170 470406 10226
rect 470462 10170 500754 10226
rect 500810 10170 500878 10226
rect 500934 10170 501002 10226
rect 501058 10170 501126 10226
rect 501182 10170 531474 10226
rect 531530 10170 531598 10226
rect 531654 10170 531722 10226
rect 531778 10170 531846 10226
rect 531902 10170 562194 10226
rect 562250 10170 562318 10226
rect 562374 10170 562442 10226
rect 562498 10170 562566 10226
rect 562622 10170 592914 10226
rect 592970 10170 593038 10226
rect 593094 10170 593162 10226
rect 593218 10170 593286 10226
rect 593342 10170 597456 10226
rect 597512 10170 597580 10226
rect 597636 10170 597704 10226
rect 597760 10170 597828 10226
rect 597884 10170 597980 10226
rect -1916 10102 597980 10170
rect -1916 10046 -1820 10102
rect -1764 10046 -1696 10102
rect -1640 10046 -1572 10102
rect -1516 10046 -1448 10102
rect -1392 10046 9234 10102
rect 9290 10046 9358 10102
rect 9414 10046 9482 10102
rect 9538 10046 9606 10102
rect 9662 10046 31878 10102
rect 31934 10046 32002 10102
rect 32058 10046 39954 10102
rect 40010 10046 40078 10102
rect 40134 10046 40202 10102
rect 40258 10046 40326 10102
rect 40382 10046 62598 10102
rect 62654 10046 62722 10102
rect 62778 10046 70674 10102
rect 70730 10046 70798 10102
rect 70854 10046 70922 10102
rect 70978 10046 71046 10102
rect 71102 10046 93318 10102
rect 93374 10046 93442 10102
rect 93498 10046 101394 10102
rect 101450 10046 101518 10102
rect 101574 10046 101642 10102
rect 101698 10046 101766 10102
rect 101822 10046 132114 10102
rect 132170 10046 132238 10102
rect 132294 10046 132362 10102
rect 132418 10046 132486 10102
rect 132542 10046 162834 10102
rect 162890 10046 162958 10102
rect 163014 10046 163082 10102
rect 163138 10046 163206 10102
rect 163262 10046 193554 10102
rect 193610 10046 193678 10102
rect 193734 10046 193802 10102
rect 193858 10046 193926 10102
rect 193982 10046 224274 10102
rect 224330 10046 224398 10102
rect 224454 10046 224522 10102
rect 224578 10046 224646 10102
rect 224702 10046 254994 10102
rect 255050 10046 255118 10102
rect 255174 10046 255242 10102
rect 255298 10046 255366 10102
rect 255422 10046 285714 10102
rect 285770 10046 285838 10102
rect 285894 10046 285962 10102
rect 286018 10046 286086 10102
rect 286142 10046 316434 10102
rect 316490 10046 316558 10102
rect 316614 10046 316682 10102
rect 316738 10046 316806 10102
rect 316862 10046 347154 10102
rect 347210 10046 347278 10102
rect 347334 10046 347402 10102
rect 347458 10046 347526 10102
rect 347582 10046 377874 10102
rect 377930 10046 377998 10102
rect 378054 10046 378122 10102
rect 378178 10046 378246 10102
rect 378302 10046 408594 10102
rect 408650 10046 408718 10102
rect 408774 10046 408842 10102
rect 408898 10046 408966 10102
rect 409022 10046 439314 10102
rect 439370 10046 439438 10102
rect 439494 10046 439562 10102
rect 439618 10046 439686 10102
rect 439742 10046 470034 10102
rect 470090 10046 470158 10102
rect 470214 10046 470282 10102
rect 470338 10046 470406 10102
rect 470462 10046 500754 10102
rect 500810 10046 500878 10102
rect 500934 10046 501002 10102
rect 501058 10046 501126 10102
rect 501182 10046 531474 10102
rect 531530 10046 531598 10102
rect 531654 10046 531722 10102
rect 531778 10046 531846 10102
rect 531902 10046 562194 10102
rect 562250 10046 562318 10102
rect 562374 10046 562442 10102
rect 562498 10046 562566 10102
rect 562622 10046 592914 10102
rect 592970 10046 593038 10102
rect 593094 10046 593162 10102
rect 593218 10046 593286 10102
rect 593342 10046 597456 10102
rect 597512 10046 597580 10102
rect 597636 10046 597704 10102
rect 597760 10046 597828 10102
rect 597884 10046 597980 10102
rect -1916 9978 597980 10046
rect -1916 9922 -1820 9978
rect -1764 9922 -1696 9978
rect -1640 9922 -1572 9978
rect -1516 9922 -1448 9978
rect -1392 9922 9234 9978
rect 9290 9922 9358 9978
rect 9414 9922 9482 9978
rect 9538 9922 9606 9978
rect 9662 9922 31878 9978
rect 31934 9922 32002 9978
rect 32058 9922 39954 9978
rect 40010 9922 40078 9978
rect 40134 9922 40202 9978
rect 40258 9922 40326 9978
rect 40382 9922 62598 9978
rect 62654 9922 62722 9978
rect 62778 9922 70674 9978
rect 70730 9922 70798 9978
rect 70854 9922 70922 9978
rect 70978 9922 71046 9978
rect 71102 9922 93318 9978
rect 93374 9922 93442 9978
rect 93498 9922 101394 9978
rect 101450 9922 101518 9978
rect 101574 9922 101642 9978
rect 101698 9922 101766 9978
rect 101822 9922 132114 9978
rect 132170 9922 132238 9978
rect 132294 9922 132362 9978
rect 132418 9922 132486 9978
rect 132542 9922 162834 9978
rect 162890 9922 162958 9978
rect 163014 9922 163082 9978
rect 163138 9922 163206 9978
rect 163262 9922 193554 9978
rect 193610 9922 193678 9978
rect 193734 9922 193802 9978
rect 193858 9922 193926 9978
rect 193982 9922 224274 9978
rect 224330 9922 224398 9978
rect 224454 9922 224522 9978
rect 224578 9922 224646 9978
rect 224702 9922 254994 9978
rect 255050 9922 255118 9978
rect 255174 9922 255242 9978
rect 255298 9922 255366 9978
rect 255422 9922 285714 9978
rect 285770 9922 285838 9978
rect 285894 9922 285962 9978
rect 286018 9922 286086 9978
rect 286142 9922 316434 9978
rect 316490 9922 316558 9978
rect 316614 9922 316682 9978
rect 316738 9922 316806 9978
rect 316862 9922 347154 9978
rect 347210 9922 347278 9978
rect 347334 9922 347402 9978
rect 347458 9922 347526 9978
rect 347582 9922 377874 9978
rect 377930 9922 377998 9978
rect 378054 9922 378122 9978
rect 378178 9922 378246 9978
rect 378302 9922 408594 9978
rect 408650 9922 408718 9978
rect 408774 9922 408842 9978
rect 408898 9922 408966 9978
rect 409022 9922 439314 9978
rect 439370 9922 439438 9978
rect 439494 9922 439562 9978
rect 439618 9922 439686 9978
rect 439742 9922 470034 9978
rect 470090 9922 470158 9978
rect 470214 9922 470282 9978
rect 470338 9922 470406 9978
rect 470462 9922 500754 9978
rect 500810 9922 500878 9978
rect 500934 9922 501002 9978
rect 501058 9922 501126 9978
rect 501182 9922 531474 9978
rect 531530 9922 531598 9978
rect 531654 9922 531722 9978
rect 531778 9922 531846 9978
rect 531902 9922 562194 9978
rect 562250 9922 562318 9978
rect 562374 9922 562442 9978
rect 562498 9922 562566 9978
rect 562622 9922 592914 9978
rect 592970 9922 593038 9978
rect 593094 9922 593162 9978
rect 593218 9922 593286 9978
rect 593342 9922 597456 9978
rect 597512 9922 597580 9978
rect 597636 9922 597704 9978
rect 597760 9922 597828 9978
rect 597884 9922 597980 9978
rect -1916 9826 597980 9922
rect 77292 9118 163732 9134
rect 77292 9062 77308 9118
rect 77364 9062 163660 9118
rect 163716 9062 163732 9118
rect 77292 9046 163732 9062
rect 53212 8938 169444 8954
rect 53212 8882 53228 8938
rect 53284 8882 169372 8938
rect 169428 8882 169444 8938
rect 53212 8866 169444 8882
rect 92412 8758 422676 8774
rect 92412 8702 92428 8758
rect 92484 8702 422604 8758
rect 422660 8702 422676 8758
rect 92412 8686 422676 8702
rect 43132 8578 83652 8594
rect 43132 8522 43148 8578
rect 43204 8522 83580 8578
rect 83636 8522 83652 8578
rect 43132 8506 83652 8522
rect 90732 8578 457060 8594
rect 90732 8522 90748 8578
rect 90804 8522 456988 8578
rect 457044 8522 457060 8578
rect 90732 8506 457060 8522
rect 44924 7858 99108 7874
rect 44924 7802 44940 7858
rect 44996 7802 99036 7858
rect 99092 7802 99108 7858
rect 44924 7786 99108 7802
rect 53660 7678 59796 7694
rect 53660 7622 53676 7678
rect 53732 7622 59724 7678
rect 59780 7622 59796 7678
rect 53660 7606 59796 7622
rect 94876 7498 108404 7514
rect 94876 7442 94892 7498
rect 94948 7442 108332 7498
rect 108388 7442 108404 7498
rect 94876 7426 108404 7442
rect 57916 7318 209428 7334
rect 57916 7262 57932 7318
rect 57988 7262 209356 7318
rect 209412 7262 209428 7318
rect 57916 7246 209428 7262
rect 63740 7138 257140 7154
rect 63740 7082 63756 7138
rect 63812 7082 257068 7138
rect 257124 7082 257140 7138
rect 63740 7066 257140 7082
rect 95324 6958 103476 6974
rect 95324 6902 95340 6958
rect 95396 6902 103404 6958
rect 103460 6902 103476 6958
rect 95324 6886 103476 6902
rect 108316 6958 468372 6974
rect 108316 6902 108332 6958
rect 108388 6902 468300 6958
rect 468356 6902 468372 6958
rect 108316 6886 468372 6902
rect 57020 6778 63044 6794
rect 57020 6722 57036 6778
rect 57092 6722 62972 6778
rect 63028 6722 63044 6778
rect 57020 6706 63044 6722
rect 81884 6778 85724 6794
rect 81884 6722 81900 6778
rect 81956 6722 85724 6778
rect 81884 6706 85724 6722
rect 99580 6778 563572 6794
rect 99580 6722 99596 6778
rect 99652 6722 563500 6778
rect 563556 6722 563572 6778
rect 99580 6706 563572 6722
rect 65196 6598 68420 6614
rect 65196 6542 65212 6598
rect 65268 6542 68348 6598
rect 68404 6542 68420 6598
rect 65196 6526 68420 6542
rect 85636 5894 85724 6706
rect 87372 6058 100116 6074
rect 87372 6002 87388 6058
rect 87444 6002 100044 6058
rect 100100 6002 100116 6058
rect 87372 5986 100116 6002
rect 85636 5878 409348 5894
rect 85636 5822 409276 5878
rect 409332 5822 409348 5878
rect 85636 5806 409348 5822
rect 64860 5698 268452 5714
rect 64860 5642 64876 5698
rect 64932 5642 268380 5698
rect 268436 5642 268452 5698
rect 64860 5626 268452 5642
rect 40892 5518 64836 5534
rect 40892 5462 40908 5518
rect 40964 5462 64764 5518
rect 64820 5462 64836 5518
rect 40892 5446 64836 5462
rect 82892 5518 92500 5534
rect 82892 5462 82908 5518
rect 82964 5462 92428 5518
rect 92484 5462 92500 5518
rect 82892 5446 92500 5462
rect 96332 5518 308436 5534
rect 96332 5462 96348 5518
rect 96404 5462 308364 5518
rect 308420 5462 308436 5518
rect 96332 5446 308436 5462
rect 53772 5338 78052 5354
rect 53772 5282 53788 5338
rect 53844 5282 77980 5338
rect 78036 5282 78052 5338
rect 53772 5266 78052 5282
rect 85636 5338 93284 5354
rect 85636 5282 93212 5338
rect 93268 5282 93284 5338
rect 85636 5266 93284 5282
rect 120972 5338 415060 5354
rect 120972 5282 120988 5338
rect 121044 5282 414988 5338
rect 415044 5282 415060 5338
rect 120972 5266 415060 5282
rect 85636 5174 85724 5266
rect 44252 5158 85724 5174
rect 44252 5102 44268 5158
rect 44324 5102 85724 5158
rect 44252 5086 85724 5102
rect 93868 5158 462660 5174
rect 93868 5102 93884 5158
rect 93940 5102 462588 5158
rect 462644 5102 462660 5158
rect 93868 5086 462660 5102
rect 93084 4618 103364 4634
rect 93084 4562 93100 4618
rect 93156 4562 103292 4618
rect 103348 4562 103364 4618
rect 93084 4546 103364 4562
rect -1916 4350 597980 4446
rect -1916 4294 -860 4350
rect -804 4294 -736 4350
rect -680 4294 -612 4350
rect -556 4294 -488 4350
rect -432 4294 5514 4350
rect 5570 4294 5638 4350
rect 5694 4294 5762 4350
rect 5818 4294 5886 4350
rect 5942 4294 36234 4350
rect 36290 4294 36358 4350
rect 36414 4294 36482 4350
rect 36538 4294 36606 4350
rect 36662 4294 66954 4350
rect 67010 4294 67078 4350
rect 67134 4294 67202 4350
rect 67258 4294 67326 4350
rect 67382 4294 97674 4350
rect 97730 4294 97798 4350
rect 97854 4294 97922 4350
rect 97978 4294 98046 4350
rect 98102 4294 128394 4350
rect 128450 4294 128518 4350
rect 128574 4294 128642 4350
rect 128698 4294 128766 4350
rect 128822 4294 159114 4350
rect 159170 4294 159238 4350
rect 159294 4294 159362 4350
rect 159418 4294 159486 4350
rect 159542 4294 189834 4350
rect 189890 4294 189958 4350
rect 190014 4294 190082 4350
rect 190138 4294 190206 4350
rect 190262 4294 220554 4350
rect 220610 4294 220678 4350
rect 220734 4294 220802 4350
rect 220858 4294 220926 4350
rect 220982 4294 251274 4350
rect 251330 4294 251398 4350
rect 251454 4294 251522 4350
rect 251578 4294 251646 4350
rect 251702 4294 281994 4350
rect 282050 4294 282118 4350
rect 282174 4294 282242 4350
rect 282298 4294 282366 4350
rect 282422 4294 312714 4350
rect 312770 4294 312838 4350
rect 312894 4294 312962 4350
rect 313018 4294 313086 4350
rect 313142 4294 343434 4350
rect 343490 4294 343558 4350
rect 343614 4294 343682 4350
rect 343738 4294 343806 4350
rect 343862 4294 374154 4350
rect 374210 4294 374278 4350
rect 374334 4294 374402 4350
rect 374458 4294 374526 4350
rect 374582 4294 404874 4350
rect 404930 4294 404998 4350
rect 405054 4294 405122 4350
rect 405178 4294 405246 4350
rect 405302 4294 435594 4350
rect 435650 4294 435718 4350
rect 435774 4294 435842 4350
rect 435898 4294 435966 4350
rect 436022 4294 466314 4350
rect 466370 4294 466438 4350
rect 466494 4294 466562 4350
rect 466618 4294 466686 4350
rect 466742 4294 497034 4350
rect 497090 4294 497158 4350
rect 497214 4294 497282 4350
rect 497338 4294 497406 4350
rect 497462 4294 527754 4350
rect 527810 4294 527878 4350
rect 527934 4294 528002 4350
rect 528058 4294 528126 4350
rect 528182 4294 558474 4350
rect 558530 4294 558598 4350
rect 558654 4294 558722 4350
rect 558778 4294 558846 4350
rect 558902 4294 589194 4350
rect 589250 4294 589318 4350
rect 589374 4294 589442 4350
rect 589498 4294 589566 4350
rect 589622 4294 596496 4350
rect 596552 4294 596620 4350
rect 596676 4294 596744 4350
rect 596800 4294 596868 4350
rect 596924 4294 597980 4350
rect -1916 4226 597980 4294
rect -1916 4170 -860 4226
rect -804 4170 -736 4226
rect -680 4170 -612 4226
rect -556 4170 -488 4226
rect -432 4170 5514 4226
rect 5570 4170 5638 4226
rect 5694 4170 5762 4226
rect 5818 4170 5886 4226
rect 5942 4170 36234 4226
rect 36290 4170 36358 4226
rect 36414 4170 36482 4226
rect 36538 4170 36606 4226
rect 36662 4170 66954 4226
rect 67010 4170 67078 4226
rect 67134 4170 67202 4226
rect 67258 4170 67326 4226
rect 67382 4170 97674 4226
rect 97730 4170 97798 4226
rect 97854 4170 97922 4226
rect 97978 4170 98046 4226
rect 98102 4170 128394 4226
rect 128450 4170 128518 4226
rect 128574 4170 128642 4226
rect 128698 4170 128766 4226
rect 128822 4170 159114 4226
rect 159170 4170 159238 4226
rect 159294 4170 159362 4226
rect 159418 4170 159486 4226
rect 159542 4170 189834 4226
rect 189890 4170 189958 4226
rect 190014 4170 190082 4226
rect 190138 4170 190206 4226
rect 190262 4170 220554 4226
rect 220610 4170 220678 4226
rect 220734 4170 220802 4226
rect 220858 4170 220926 4226
rect 220982 4170 251274 4226
rect 251330 4170 251398 4226
rect 251454 4170 251522 4226
rect 251578 4170 251646 4226
rect 251702 4170 281994 4226
rect 282050 4170 282118 4226
rect 282174 4170 282242 4226
rect 282298 4170 282366 4226
rect 282422 4170 312714 4226
rect 312770 4170 312838 4226
rect 312894 4170 312962 4226
rect 313018 4170 313086 4226
rect 313142 4170 343434 4226
rect 343490 4170 343558 4226
rect 343614 4170 343682 4226
rect 343738 4170 343806 4226
rect 343862 4170 374154 4226
rect 374210 4170 374278 4226
rect 374334 4170 374402 4226
rect 374458 4170 374526 4226
rect 374582 4170 404874 4226
rect 404930 4170 404998 4226
rect 405054 4170 405122 4226
rect 405178 4170 405246 4226
rect 405302 4170 435594 4226
rect 435650 4170 435718 4226
rect 435774 4170 435842 4226
rect 435898 4170 435966 4226
rect 436022 4170 466314 4226
rect 466370 4170 466438 4226
rect 466494 4170 466562 4226
rect 466618 4170 466686 4226
rect 466742 4170 497034 4226
rect 497090 4170 497158 4226
rect 497214 4170 497282 4226
rect 497338 4170 497406 4226
rect 497462 4170 527754 4226
rect 527810 4170 527878 4226
rect 527934 4170 528002 4226
rect 528058 4170 528126 4226
rect 528182 4170 558474 4226
rect 558530 4170 558598 4226
rect 558654 4170 558722 4226
rect 558778 4170 558846 4226
rect 558902 4170 589194 4226
rect 589250 4170 589318 4226
rect 589374 4170 589442 4226
rect 589498 4170 589566 4226
rect 589622 4170 596496 4226
rect 596552 4170 596620 4226
rect 596676 4170 596744 4226
rect 596800 4170 596868 4226
rect 596924 4170 597980 4226
rect -1916 4102 597980 4170
rect -1916 4046 -860 4102
rect -804 4046 -736 4102
rect -680 4046 -612 4102
rect -556 4046 -488 4102
rect -432 4046 5514 4102
rect 5570 4046 5638 4102
rect 5694 4046 5762 4102
rect 5818 4046 5886 4102
rect 5942 4046 36234 4102
rect 36290 4046 36358 4102
rect 36414 4046 36482 4102
rect 36538 4046 36606 4102
rect 36662 4046 66954 4102
rect 67010 4046 67078 4102
rect 67134 4046 67202 4102
rect 67258 4046 67326 4102
rect 67382 4046 97674 4102
rect 97730 4046 97798 4102
rect 97854 4046 97922 4102
rect 97978 4046 98046 4102
rect 98102 4046 128394 4102
rect 128450 4046 128518 4102
rect 128574 4046 128642 4102
rect 128698 4046 128766 4102
rect 128822 4046 159114 4102
rect 159170 4046 159238 4102
rect 159294 4046 159362 4102
rect 159418 4046 159486 4102
rect 159542 4046 189834 4102
rect 189890 4046 189958 4102
rect 190014 4046 190082 4102
rect 190138 4046 190206 4102
rect 190262 4046 220554 4102
rect 220610 4046 220678 4102
rect 220734 4046 220802 4102
rect 220858 4046 220926 4102
rect 220982 4046 251274 4102
rect 251330 4046 251398 4102
rect 251454 4046 251522 4102
rect 251578 4046 251646 4102
rect 251702 4046 281994 4102
rect 282050 4046 282118 4102
rect 282174 4046 282242 4102
rect 282298 4046 282366 4102
rect 282422 4046 312714 4102
rect 312770 4046 312838 4102
rect 312894 4046 312962 4102
rect 313018 4046 313086 4102
rect 313142 4046 343434 4102
rect 343490 4046 343558 4102
rect 343614 4046 343682 4102
rect 343738 4046 343806 4102
rect 343862 4046 374154 4102
rect 374210 4046 374278 4102
rect 374334 4046 374402 4102
rect 374458 4046 374526 4102
rect 374582 4046 404874 4102
rect 404930 4046 404998 4102
rect 405054 4046 405122 4102
rect 405178 4046 405246 4102
rect 405302 4046 435594 4102
rect 435650 4046 435718 4102
rect 435774 4046 435842 4102
rect 435898 4046 435966 4102
rect 436022 4046 466314 4102
rect 466370 4046 466438 4102
rect 466494 4046 466562 4102
rect 466618 4046 466686 4102
rect 466742 4046 497034 4102
rect 497090 4046 497158 4102
rect 497214 4046 497282 4102
rect 497338 4046 497406 4102
rect 497462 4046 527754 4102
rect 527810 4046 527878 4102
rect 527934 4046 528002 4102
rect 528058 4046 528126 4102
rect 528182 4046 558474 4102
rect 558530 4046 558598 4102
rect 558654 4046 558722 4102
rect 558778 4046 558846 4102
rect 558902 4046 589194 4102
rect 589250 4046 589318 4102
rect 589374 4046 589442 4102
rect 589498 4046 589566 4102
rect 589622 4046 596496 4102
rect 596552 4046 596620 4102
rect 596676 4046 596744 4102
rect 596800 4046 596868 4102
rect 596924 4046 597980 4102
rect -1916 3978 597980 4046
rect -1916 3922 -860 3978
rect -804 3922 -736 3978
rect -680 3922 -612 3978
rect -556 3922 -488 3978
rect -432 3922 5514 3978
rect 5570 3922 5638 3978
rect 5694 3922 5762 3978
rect 5818 3922 5886 3978
rect 5942 3922 36234 3978
rect 36290 3922 36358 3978
rect 36414 3922 36482 3978
rect 36538 3922 36606 3978
rect 36662 3922 66954 3978
rect 67010 3922 67078 3978
rect 67134 3922 67202 3978
rect 67258 3922 67326 3978
rect 67382 3922 97674 3978
rect 97730 3922 97798 3978
rect 97854 3922 97922 3978
rect 97978 3922 98046 3978
rect 98102 3922 128394 3978
rect 128450 3922 128518 3978
rect 128574 3922 128642 3978
rect 128698 3922 128766 3978
rect 128822 3922 159114 3978
rect 159170 3922 159238 3978
rect 159294 3922 159362 3978
rect 159418 3922 159486 3978
rect 159542 3922 189834 3978
rect 189890 3922 189958 3978
rect 190014 3922 190082 3978
rect 190138 3922 190206 3978
rect 190262 3922 220554 3978
rect 220610 3922 220678 3978
rect 220734 3922 220802 3978
rect 220858 3922 220926 3978
rect 220982 3922 251274 3978
rect 251330 3922 251398 3978
rect 251454 3922 251522 3978
rect 251578 3922 251646 3978
rect 251702 3922 281994 3978
rect 282050 3922 282118 3978
rect 282174 3922 282242 3978
rect 282298 3922 282366 3978
rect 282422 3922 312714 3978
rect 312770 3922 312838 3978
rect 312894 3922 312962 3978
rect 313018 3922 313086 3978
rect 313142 3922 343434 3978
rect 343490 3922 343558 3978
rect 343614 3922 343682 3978
rect 343738 3922 343806 3978
rect 343862 3922 374154 3978
rect 374210 3922 374278 3978
rect 374334 3922 374402 3978
rect 374458 3922 374526 3978
rect 374582 3922 404874 3978
rect 404930 3922 404998 3978
rect 405054 3922 405122 3978
rect 405178 3922 405246 3978
rect 405302 3922 435594 3978
rect 435650 3922 435718 3978
rect 435774 3922 435842 3978
rect 435898 3922 435966 3978
rect 436022 3922 466314 3978
rect 466370 3922 466438 3978
rect 466494 3922 466562 3978
rect 466618 3922 466686 3978
rect 466742 3922 497034 3978
rect 497090 3922 497158 3978
rect 497214 3922 497282 3978
rect 497338 3922 497406 3978
rect 497462 3922 527754 3978
rect 527810 3922 527878 3978
rect 527934 3922 528002 3978
rect 528058 3922 528126 3978
rect 528182 3922 558474 3978
rect 558530 3922 558598 3978
rect 558654 3922 558722 3978
rect 558778 3922 558846 3978
rect 558902 3922 589194 3978
rect 589250 3922 589318 3978
rect 589374 3922 589442 3978
rect 589498 3922 589566 3978
rect 589622 3922 596496 3978
rect 596552 3922 596620 3978
rect 596676 3922 596744 3978
rect 596800 3922 596868 3978
rect 596924 3922 597980 3978
rect -1916 3826 597980 3922
rect 46604 3718 59012 3734
rect 46604 3662 46620 3718
rect 46676 3662 58940 3718
rect 58996 3662 59012 3718
rect 46604 3646 59012 3662
rect 56124 3538 193300 3554
rect 56124 3482 56140 3538
rect 56196 3482 193228 3538
rect 193284 3482 193300 3538
rect 56124 3466 193300 3482
rect 45820 3358 106612 3374
rect 45820 3302 45836 3358
rect 45892 3302 106540 3358
rect 106596 3302 106612 3358
rect 45820 3286 106612 3302
rect 98908 3178 557860 3194
rect 98908 3122 98924 3178
rect 98980 3122 557788 3178
rect 557844 3122 557860 3178
rect 98908 3106 557860 3122
rect 56572 2998 198004 3014
rect 56572 2942 56588 2998
rect 56644 2942 197932 2998
rect 197988 2942 198004 2998
rect 56572 2926 198004 2942
rect 43804 2818 89476 2834
rect 43804 2762 43820 2818
rect 43876 2762 89404 2818
rect 89460 2762 89476 2818
rect 43804 2746 89476 2762
rect 52092 2458 118036 2474
rect 52092 2402 117964 2458
rect 118020 2402 118036 2458
rect 52092 2386 118036 2402
rect 52092 1574 52180 2386
rect 43580 1558 48148 1574
rect 43580 1502 43596 1558
rect 43652 1502 48076 1558
rect 48132 1502 48148 1558
rect 43580 1486 48148 1502
rect 48620 1558 52180 1574
rect 48620 1502 48636 1558
rect 48692 1502 52180 1558
rect 48620 1486 52180 1502
rect 56236 1558 61588 1574
rect 56236 1502 56252 1558
rect 56308 1502 61516 1558
rect 61572 1502 61588 1558
rect 56236 1486 61588 1502
rect 76284 1558 81636 1574
rect 76284 1502 76300 1558
rect 76356 1502 81564 1558
rect 81620 1502 81636 1558
rect 76284 1486 81636 1502
rect 81772 1558 89924 1574
rect 81772 1502 81788 1558
rect 81844 1502 89852 1558
rect 89908 1502 89924 1558
rect 81772 1486 89924 1502
rect 100476 1558 569620 1574
rect 100476 1502 100492 1558
rect 100548 1502 569548 1558
rect 569604 1502 569620 1558
rect 100476 1486 569620 1502
rect 52764 1378 62484 1394
rect 52764 1322 52780 1378
rect 52836 1322 62412 1378
rect 62468 1322 62484 1378
rect 52764 1306 62484 1322
rect 99132 1378 542628 1394
rect 99132 1322 99148 1378
rect 99204 1322 542556 1378
rect 542612 1322 542628 1378
rect 99132 1306 542628 1322
rect 58028 1198 65844 1214
rect 58028 1142 58044 1198
rect 58100 1142 65772 1198
rect 65828 1142 65844 1198
rect 58028 1126 65844 1142
rect 98460 1198 130244 1214
rect 98460 1142 98476 1198
rect 98532 1142 130172 1198
rect 130228 1142 130244 1198
rect 98460 1126 130244 1142
rect 53436 1018 85780 1034
rect 53436 962 53452 1018
rect 53508 962 85708 1018
rect 85764 962 85780 1018
rect 53436 946 85780 962
rect 58140 118 211332 134
rect 58140 62 58156 118
rect 58212 62 211260 118
rect 211316 62 211332 118
rect 58140 46 211332 62
rect -956 -160 597020 -64
rect -956 -216 -860 -160
rect -804 -216 -736 -160
rect -680 -216 -612 -160
rect -556 -216 -488 -160
rect -432 -216 5514 -160
rect 5570 -216 5638 -160
rect 5694 -216 5762 -160
rect 5818 -216 5886 -160
rect 5942 -216 36234 -160
rect 36290 -216 36358 -160
rect 36414 -216 36482 -160
rect 36538 -216 36606 -160
rect 36662 -216 66954 -160
rect 67010 -216 67078 -160
rect 67134 -216 67202 -160
rect 67258 -216 67326 -160
rect 67382 -216 97674 -160
rect 97730 -216 97798 -160
rect 97854 -216 97922 -160
rect 97978 -216 98046 -160
rect 98102 -216 128394 -160
rect 128450 -216 128518 -160
rect 128574 -216 128642 -160
rect 128698 -216 128766 -160
rect 128822 -216 159114 -160
rect 159170 -216 159238 -160
rect 159294 -216 159362 -160
rect 159418 -216 159486 -160
rect 159542 -216 189834 -160
rect 189890 -216 189958 -160
rect 190014 -216 190082 -160
rect 190138 -216 190206 -160
rect 190262 -216 220554 -160
rect 220610 -216 220678 -160
rect 220734 -216 220802 -160
rect 220858 -216 220926 -160
rect 220982 -216 251274 -160
rect 251330 -216 251398 -160
rect 251454 -216 251522 -160
rect 251578 -216 251646 -160
rect 251702 -216 281994 -160
rect 282050 -216 282118 -160
rect 282174 -216 282242 -160
rect 282298 -216 282366 -160
rect 282422 -216 312714 -160
rect 312770 -216 312838 -160
rect 312894 -216 312962 -160
rect 313018 -216 313086 -160
rect 313142 -216 343434 -160
rect 343490 -216 343558 -160
rect 343614 -216 343682 -160
rect 343738 -216 343806 -160
rect 343862 -216 374154 -160
rect 374210 -216 374278 -160
rect 374334 -216 374402 -160
rect 374458 -216 374526 -160
rect 374582 -216 404874 -160
rect 404930 -216 404998 -160
rect 405054 -216 405122 -160
rect 405178 -216 405246 -160
rect 405302 -216 435594 -160
rect 435650 -216 435718 -160
rect 435774 -216 435842 -160
rect 435898 -216 435966 -160
rect 436022 -216 466314 -160
rect 466370 -216 466438 -160
rect 466494 -216 466562 -160
rect 466618 -216 466686 -160
rect 466742 -216 497034 -160
rect 497090 -216 497158 -160
rect 497214 -216 497282 -160
rect 497338 -216 497406 -160
rect 497462 -216 527754 -160
rect 527810 -216 527878 -160
rect 527934 -216 528002 -160
rect 528058 -216 528126 -160
rect 528182 -216 558474 -160
rect 558530 -216 558598 -160
rect 558654 -216 558722 -160
rect 558778 -216 558846 -160
rect 558902 -216 589194 -160
rect 589250 -216 589318 -160
rect 589374 -216 589442 -160
rect 589498 -216 589566 -160
rect 589622 -216 596496 -160
rect 596552 -216 596620 -160
rect 596676 -216 596744 -160
rect 596800 -216 596868 -160
rect 596924 -216 597020 -160
rect -956 -284 597020 -216
rect -956 -340 -860 -284
rect -804 -340 -736 -284
rect -680 -340 -612 -284
rect -556 -340 -488 -284
rect -432 -340 5514 -284
rect 5570 -340 5638 -284
rect 5694 -340 5762 -284
rect 5818 -340 5886 -284
rect 5942 -340 36234 -284
rect 36290 -340 36358 -284
rect 36414 -340 36482 -284
rect 36538 -340 36606 -284
rect 36662 -340 66954 -284
rect 67010 -340 67078 -284
rect 67134 -340 67202 -284
rect 67258 -340 67326 -284
rect 67382 -340 97674 -284
rect 97730 -340 97798 -284
rect 97854 -340 97922 -284
rect 97978 -340 98046 -284
rect 98102 -340 128394 -284
rect 128450 -340 128518 -284
rect 128574 -340 128642 -284
rect 128698 -340 128766 -284
rect 128822 -340 159114 -284
rect 159170 -340 159238 -284
rect 159294 -340 159362 -284
rect 159418 -340 159486 -284
rect 159542 -340 189834 -284
rect 189890 -340 189958 -284
rect 190014 -340 190082 -284
rect 190138 -340 190206 -284
rect 190262 -340 220554 -284
rect 220610 -340 220678 -284
rect 220734 -340 220802 -284
rect 220858 -340 220926 -284
rect 220982 -340 251274 -284
rect 251330 -340 251398 -284
rect 251454 -340 251522 -284
rect 251578 -340 251646 -284
rect 251702 -340 281994 -284
rect 282050 -340 282118 -284
rect 282174 -340 282242 -284
rect 282298 -340 282366 -284
rect 282422 -340 312714 -284
rect 312770 -340 312838 -284
rect 312894 -340 312962 -284
rect 313018 -340 313086 -284
rect 313142 -340 343434 -284
rect 343490 -340 343558 -284
rect 343614 -340 343682 -284
rect 343738 -340 343806 -284
rect 343862 -340 374154 -284
rect 374210 -340 374278 -284
rect 374334 -340 374402 -284
rect 374458 -340 374526 -284
rect 374582 -340 404874 -284
rect 404930 -340 404998 -284
rect 405054 -340 405122 -284
rect 405178 -340 405246 -284
rect 405302 -340 435594 -284
rect 435650 -340 435718 -284
rect 435774 -340 435842 -284
rect 435898 -340 435966 -284
rect 436022 -340 466314 -284
rect 466370 -340 466438 -284
rect 466494 -340 466562 -284
rect 466618 -340 466686 -284
rect 466742 -340 497034 -284
rect 497090 -340 497158 -284
rect 497214 -340 497282 -284
rect 497338 -340 497406 -284
rect 497462 -340 527754 -284
rect 527810 -340 527878 -284
rect 527934 -340 528002 -284
rect 528058 -340 528126 -284
rect 528182 -340 558474 -284
rect 558530 -340 558598 -284
rect 558654 -340 558722 -284
rect 558778 -340 558846 -284
rect 558902 -340 589194 -284
rect 589250 -340 589318 -284
rect 589374 -340 589442 -284
rect 589498 -340 589566 -284
rect 589622 -340 596496 -284
rect 596552 -340 596620 -284
rect 596676 -340 596744 -284
rect 596800 -340 596868 -284
rect 596924 -340 597020 -284
rect -956 -408 597020 -340
rect -956 -464 -860 -408
rect -804 -464 -736 -408
rect -680 -464 -612 -408
rect -556 -464 -488 -408
rect -432 -464 5514 -408
rect 5570 -464 5638 -408
rect 5694 -464 5762 -408
rect 5818 -464 5886 -408
rect 5942 -464 36234 -408
rect 36290 -464 36358 -408
rect 36414 -464 36482 -408
rect 36538 -464 36606 -408
rect 36662 -464 66954 -408
rect 67010 -464 67078 -408
rect 67134 -464 67202 -408
rect 67258 -464 67326 -408
rect 67382 -464 97674 -408
rect 97730 -464 97798 -408
rect 97854 -464 97922 -408
rect 97978 -464 98046 -408
rect 98102 -464 128394 -408
rect 128450 -464 128518 -408
rect 128574 -464 128642 -408
rect 128698 -464 128766 -408
rect 128822 -464 159114 -408
rect 159170 -464 159238 -408
rect 159294 -464 159362 -408
rect 159418 -464 159486 -408
rect 159542 -464 189834 -408
rect 189890 -464 189958 -408
rect 190014 -464 190082 -408
rect 190138 -464 190206 -408
rect 190262 -464 220554 -408
rect 220610 -464 220678 -408
rect 220734 -464 220802 -408
rect 220858 -464 220926 -408
rect 220982 -464 251274 -408
rect 251330 -464 251398 -408
rect 251454 -464 251522 -408
rect 251578 -464 251646 -408
rect 251702 -464 281994 -408
rect 282050 -464 282118 -408
rect 282174 -464 282242 -408
rect 282298 -464 282366 -408
rect 282422 -464 312714 -408
rect 312770 -464 312838 -408
rect 312894 -464 312962 -408
rect 313018 -464 313086 -408
rect 313142 -464 343434 -408
rect 343490 -464 343558 -408
rect 343614 -464 343682 -408
rect 343738 -464 343806 -408
rect 343862 -464 374154 -408
rect 374210 -464 374278 -408
rect 374334 -464 374402 -408
rect 374458 -464 374526 -408
rect 374582 -464 404874 -408
rect 404930 -464 404998 -408
rect 405054 -464 405122 -408
rect 405178 -464 405246 -408
rect 405302 -464 435594 -408
rect 435650 -464 435718 -408
rect 435774 -464 435842 -408
rect 435898 -464 435966 -408
rect 436022 -464 466314 -408
rect 466370 -464 466438 -408
rect 466494 -464 466562 -408
rect 466618 -464 466686 -408
rect 466742 -464 497034 -408
rect 497090 -464 497158 -408
rect 497214 -464 497282 -408
rect 497338 -464 497406 -408
rect 497462 -464 527754 -408
rect 527810 -464 527878 -408
rect 527934 -464 528002 -408
rect 528058 -464 528126 -408
rect 528182 -464 558474 -408
rect 558530 -464 558598 -408
rect 558654 -464 558722 -408
rect 558778 -464 558846 -408
rect 558902 -464 589194 -408
rect 589250 -464 589318 -408
rect 589374 -464 589442 -408
rect 589498 -464 589566 -408
rect 589622 -464 596496 -408
rect 596552 -464 596620 -408
rect 596676 -464 596744 -408
rect 596800 -464 596868 -408
rect 596924 -464 597020 -408
rect -956 -532 597020 -464
rect -956 -588 -860 -532
rect -804 -588 -736 -532
rect -680 -588 -612 -532
rect -556 -588 -488 -532
rect -432 -588 5514 -532
rect 5570 -588 5638 -532
rect 5694 -588 5762 -532
rect 5818 -588 5886 -532
rect 5942 -588 36234 -532
rect 36290 -588 36358 -532
rect 36414 -588 36482 -532
rect 36538 -588 36606 -532
rect 36662 -588 66954 -532
rect 67010 -588 67078 -532
rect 67134 -588 67202 -532
rect 67258 -588 67326 -532
rect 67382 -588 97674 -532
rect 97730 -588 97798 -532
rect 97854 -588 97922 -532
rect 97978 -588 98046 -532
rect 98102 -588 128394 -532
rect 128450 -588 128518 -532
rect 128574 -588 128642 -532
rect 128698 -588 128766 -532
rect 128822 -588 159114 -532
rect 159170 -588 159238 -532
rect 159294 -588 159362 -532
rect 159418 -588 159486 -532
rect 159542 -588 189834 -532
rect 189890 -588 189958 -532
rect 190014 -588 190082 -532
rect 190138 -588 190206 -532
rect 190262 -588 220554 -532
rect 220610 -588 220678 -532
rect 220734 -588 220802 -532
rect 220858 -588 220926 -532
rect 220982 -588 251274 -532
rect 251330 -588 251398 -532
rect 251454 -588 251522 -532
rect 251578 -588 251646 -532
rect 251702 -588 281994 -532
rect 282050 -588 282118 -532
rect 282174 -588 282242 -532
rect 282298 -588 282366 -532
rect 282422 -588 312714 -532
rect 312770 -588 312838 -532
rect 312894 -588 312962 -532
rect 313018 -588 313086 -532
rect 313142 -588 343434 -532
rect 343490 -588 343558 -532
rect 343614 -588 343682 -532
rect 343738 -588 343806 -532
rect 343862 -588 374154 -532
rect 374210 -588 374278 -532
rect 374334 -588 374402 -532
rect 374458 -588 374526 -532
rect 374582 -588 404874 -532
rect 404930 -588 404998 -532
rect 405054 -588 405122 -532
rect 405178 -588 405246 -532
rect 405302 -588 435594 -532
rect 435650 -588 435718 -532
rect 435774 -588 435842 -532
rect 435898 -588 435966 -532
rect 436022 -588 466314 -532
rect 466370 -588 466438 -532
rect 466494 -588 466562 -532
rect 466618 -588 466686 -532
rect 466742 -588 497034 -532
rect 497090 -588 497158 -532
rect 497214 -588 497282 -532
rect 497338 -588 497406 -532
rect 497462 -588 527754 -532
rect 527810 -588 527878 -532
rect 527934 -588 528002 -532
rect 528058 -588 528126 -532
rect 528182 -588 558474 -532
rect 558530 -588 558598 -532
rect 558654 -588 558722 -532
rect 558778 -588 558846 -532
rect 558902 -588 589194 -532
rect 589250 -588 589318 -532
rect 589374 -588 589442 -532
rect 589498 -588 589566 -532
rect 589622 -588 596496 -532
rect 596552 -588 596620 -532
rect 596676 -588 596744 -532
rect 596800 -588 596868 -532
rect 596924 -588 597020 -532
rect -956 -684 597020 -588
rect -1916 -1120 597980 -1024
rect -1916 -1176 -1820 -1120
rect -1764 -1176 -1696 -1120
rect -1640 -1176 -1572 -1120
rect -1516 -1176 -1448 -1120
rect -1392 -1176 9234 -1120
rect 9290 -1176 9358 -1120
rect 9414 -1176 9482 -1120
rect 9538 -1176 9606 -1120
rect 9662 -1176 39954 -1120
rect 40010 -1176 40078 -1120
rect 40134 -1176 40202 -1120
rect 40258 -1176 40326 -1120
rect 40382 -1176 70674 -1120
rect 70730 -1176 70798 -1120
rect 70854 -1176 70922 -1120
rect 70978 -1176 71046 -1120
rect 71102 -1176 101394 -1120
rect 101450 -1176 101518 -1120
rect 101574 -1176 101642 -1120
rect 101698 -1176 101766 -1120
rect 101822 -1176 132114 -1120
rect 132170 -1176 132238 -1120
rect 132294 -1176 132362 -1120
rect 132418 -1176 132486 -1120
rect 132542 -1176 162834 -1120
rect 162890 -1176 162958 -1120
rect 163014 -1176 163082 -1120
rect 163138 -1176 163206 -1120
rect 163262 -1176 193554 -1120
rect 193610 -1176 193678 -1120
rect 193734 -1176 193802 -1120
rect 193858 -1176 193926 -1120
rect 193982 -1176 224274 -1120
rect 224330 -1176 224398 -1120
rect 224454 -1176 224522 -1120
rect 224578 -1176 224646 -1120
rect 224702 -1176 254994 -1120
rect 255050 -1176 255118 -1120
rect 255174 -1176 255242 -1120
rect 255298 -1176 255366 -1120
rect 255422 -1176 285714 -1120
rect 285770 -1176 285838 -1120
rect 285894 -1176 285962 -1120
rect 286018 -1176 286086 -1120
rect 286142 -1176 316434 -1120
rect 316490 -1176 316558 -1120
rect 316614 -1176 316682 -1120
rect 316738 -1176 316806 -1120
rect 316862 -1176 347154 -1120
rect 347210 -1176 347278 -1120
rect 347334 -1176 347402 -1120
rect 347458 -1176 347526 -1120
rect 347582 -1176 377874 -1120
rect 377930 -1176 377998 -1120
rect 378054 -1176 378122 -1120
rect 378178 -1176 378246 -1120
rect 378302 -1176 408594 -1120
rect 408650 -1176 408718 -1120
rect 408774 -1176 408842 -1120
rect 408898 -1176 408966 -1120
rect 409022 -1176 439314 -1120
rect 439370 -1176 439438 -1120
rect 439494 -1176 439562 -1120
rect 439618 -1176 439686 -1120
rect 439742 -1176 470034 -1120
rect 470090 -1176 470158 -1120
rect 470214 -1176 470282 -1120
rect 470338 -1176 470406 -1120
rect 470462 -1176 500754 -1120
rect 500810 -1176 500878 -1120
rect 500934 -1176 501002 -1120
rect 501058 -1176 501126 -1120
rect 501182 -1176 531474 -1120
rect 531530 -1176 531598 -1120
rect 531654 -1176 531722 -1120
rect 531778 -1176 531846 -1120
rect 531902 -1176 562194 -1120
rect 562250 -1176 562318 -1120
rect 562374 -1176 562442 -1120
rect 562498 -1176 562566 -1120
rect 562622 -1176 592914 -1120
rect 592970 -1176 593038 -1120
rect 593094 -1176 593162 -1120
rect 593218 -1176 593286 -1120
rect 593342 -1176 597456 -1120
rect 597512 -1176 597580 -1120
rect 597636 -1176 597704 -1120
rect 597760 -1176 597828 -1120
rect 597884 -1176 597980 -1120
rect -1916 -1244 597980 -1176
rect -1916 -1300 -1820 -1244
rect -1764 -1300 -1696 -1244
rect -1640 -1300 -1572 -1244
rect -1516 -1300 -1448 -1244
rect -1392 -1300 9234 -1244
rect 9290 -1300 9358 -1244
rect 9414 -1300 9482 -1244
rect 9538 -1300 9606 -1244
rect 9662 -1300 39954 -1244
rect 40010 -1300 40078 -1244
rect 40134 -1300 40202 -1244
rect 40258 -1300 40326 -1244
rect 40382 -1300 70674 -1244
rect 70730 -1300 70798 -1244
rect 70854 -1300 70922 -1244
rect 70978 -1300 71046 -1244
rect 71102 -1300 101394 -1244
rect 101450 -1300 101518 -1244
rect 101574 -1300 101642 -1244
rect 101698 -1300 101766 -1244
rect 101822 -1300 132114 -1244
rect 132170 -1300 132238 -1244
rect 132294 -1300 132362 -1244
rect 132418 -1300 132486 -1244
rect 132542 -1300 162834 -1244
rect 162890 -1300 162958 -1244
rect 163014 -1300 163082 -1244
rect 163138 -1300 163206 -1244
rect 163262 -1300 193554 -1244
rect 193610 -1300 193678 -1244
rect 193734 -1300 193802 -1244
rect 193858 -1300 193926 -1244
rect 193982 -1300 224274 -1244
rect 224330 -1300 224398 -1244
rect 224454 -1300 224522 -1244
rect 224578 -1300 224646 -1244
rect 224702 -1300 254994 -1244
rect 255050 -1300 255118 -1244
rect 255174 -1300 255242 -1244
rect 255298 -1300 255366 -1244
rect 255422 -1300 285714 -1244
rect 285770 -1300 285838 -1244
rect 285894 -1300 285962 -1244
rect 286018 -1300 286086 -1244
rect 286142 -1300 316434 -1244
rect 316490 -1300 316558 -1244
rect 316614 -1300 316682 -1244
rect 316738 -1300 316806 -1244
rect 316862 -1300 347154 -1244
rect 347210 -1300 347278 -1244
rect 347334 -1300 347402 -1244
rect 347458 -1300 347526 -1244
rect 347582 -1300 377874 -1244
rect 377930 -1300 377998 -1244
rect 378054 -1300 378122 -1244
rect 378178 -1300 378246 -1244
rect 378302 -1300 408594 -1244
rect 408650 -1300 408718 -1244
rect 408774 -1300 408842 -1244
rect 408898 -1300 408966 -1244
rect 409022 -1300 439314 -1244
rect 439370 -1300 439438 -1244
rect 439494 -1300 439562 -1244
rect 439618 -1300 439686 -1244
rect 439742 -1300 470034 -1244
rect 470090 -1300 470158 -1244
rect 470214 -1300 470282 -1244
rect 470338 -1300 470406 -1244
rect 470462 -1300 500754 -1244
rect 500810 -1300 500878 -1244
rect 500934 -1300 501002 -1244
rect 501058 -1300 501126 -1244
rect 501182 -1300 531474 -1244
rect 531530 -1300 531598 -1244
rect 531654 -1300 531722 -1244
rect 531778 -1300 531846 -1244
rect 531902 -1300 562194 -1244
rect 562250 -1300 562318 -1244
rect 562374 -1300 562442 -1244
rect 562498 -1300 562566 -1244
rect 562622 -1300 592914 -1244
rect 592970 -1300 593038 -1244
rect 593094 -1300 593162 -1244
rect 593218 -1300 593286 -1244
rect 593342 -1300 597456 -1244
rect 597512 -1300 597580 -1244
rect 597636 -1300 597704 -1244
rect 597760 -1300 597828 -1244
rect 597884 -1300 597980 -1244
rect -1916 -1368 597980 -1300
rect -1916 -1424 -1820 -1368
rect -1764 -1424 -1696 -1368
rect -1640 -1424 -1572 -1368
rect -1516 -1424 -1448 -1368
rect -1392 -1424 9234 -1368
rect 9290 -1424 9358 -1368
rect 9414 -1424 9482 -1368
rect 9538 -1424 9606 -1368
rect 9662 -1424 39954 -1368
rect 40010 -1424 40078 -1368
rect 40134 -1424 40202 -1368
rect 40258 -1424 40326 -1368
rect 40382 -1424 70674 -1368
rect 70730 -1424 70798 -1368
rect 70854 -1424 70922 -1368
rect 70978 -1424 71046 -1368
rect 71102 -1424 101394 -1368
rect 101450 -1424 101518 -1368
rect 101574 -1424 101642 -1368
rect 101698 -1424 101766 -1368
rect 101822 -1424 132114 -1368
rect 132170 -1424 132238 -1368
rect 132294 -1424 132362 -1368
rect 132418 -1424 132486 -1368
rect 132542 -1424 162834 -1368
rect 162890 -1424 162958 -1368
rect 163014 -1424 163082 -1368
rect 163138 -1424 163206 -1368
rect 163262 -1424 193554 -1368
rect 193610 -1424 193678 -1368
rect 193734 -1424 193802 -1368
rect 193858 -1424 193926 -1368
rect 193982 -1424 224274 -1368
rect 224330 -1424 224398 -1368
rect 224454 -1424 224522 -1368
rect 224578 -1424 224646 -1368
rect 224702 -1424 254994 -1368
rect 255050 -1424 255118 -1368
rect 255174 -1424 255242 -1368
rect 255298 -1424 255366 -1368
rect 255422 -1424 285714 -1368
rect 285770 -1424 285838 -1368
rect 285894 -1424 285962 -1368
rect 286018 -1424 286086 -1368
rect 286142 -1424 316434 -1368
rect 316490 -1424 316558 -1368
rect 316614 -1424 316682 -1368
rect 316738 -1424 316806 -1368
rect 316862 -1424 347154 -1368
rect 347210 -1424 347278 -1368
rect 347334 -1424 347402 -1368
rect 347458 -1424 347526 -1368
rect 347582 -1424 377874 -1368
rect 377930 -1424 377998 -1368
rect 378054 -1424 378122 -1368
rect 378178 -1424 378246 -1368
rect 378302 -1424 408594 -1368
rect 408650 -1424 408718 -1368
rect 408774 -1424 408842 -1368
rect 408898 -1424 408966 -1368
rect 409022 -1424 439314 -1368
rect 439370 -1424 439438 -1368
rect 439494 -1424 439562 -1368
rect 439618 -1424 439686 -1368
rect 439742 -1424 470034 -1368
rect 470090 -1424 470158 -1368
rect 470214 -1424 470282 -1368
rect 470338 -1424 470406 -1368
rect 470462 -1424 500754 -1368
rect 500810 -1424 500878 -1368
rect 500934 -1424 501002 -1368
rect 501058 -1424 501126 -1368
rect 501182 -1424 531474 -1368
rect 531530 -1424 531598 -1368
rect 531654 -1424 531722 -1368
rect 531778 -1424 531846 -1368
rect 531902 -1424 562194 -1368
rect 562250 -1424 562318 -1368
rect 562374 -1424 562442 -1368
rect 562498 -1424 562566 -1368
rect 562622 -1424 592914 -1368
rect 592970 -1424 593038 -1368
rect 593094 -1424 593162 -1368
rect 593218 -1424 593286 -1368
rect 593342 -1424 597456 -1368
rect 597512 -1424 597580 -1368
rect 597636 -1424 597704 -1368
rect 597760 -1424 597828 -1368
rect 597884 -1424 597980 -1368
rect -1916 -1492 597980 -1424
rect -1916 -1548 -1820 -1492
rect -1764 -1548 -1696 -1492
rect -1640 -1548 -1572 -1492
rect -1516 -1548 -1448 -1492
rect -1392 -1548 9234 -1492
rect 9290 -1548 9358 -1492
rect 9414 -1548 9482 -1492
rect 9538 -1548 9606 -1492
rect 9662 -1548 39954 -1492
rect 40010 -1548 40078 -1492
rect 40134 -1548 40202 -1492
rect 40258 -1548 40326 -1492
rect 40382 -1548 70674 -1492
rect 70730 -1548 70798 -1492
rect 70854 -1548 70922 -1492
rect 70978 -1548 71046 -1492
rect 71102 -1548 101394 -1492
rect 101450 -1548 101518 -1492
rect 101574 -1548 101642 -1492
rect 101698 -1548 101766 -1492
rect 101822 -1548 132114 -1492
rect 132170 -1548 132238 -1492
rect 132294 -1548 132362 -1492
rect 132418 -1548 132486 -1492
rect 132542 -1548 162834 -1492
rect 162890 -1548 162958 -1492
rect 163014 -1548 163082 -1492
rect 163138 -1548 163206 -1492
rect 163262 -1548 193554 -1492
rect 193610 -1548 193678 -1492
rect 193734 -1548 193802 -1492
rect 193858 -1548 193926 -1492
rect 193982 -1548 224274 -1492
rect 224330 -1548 224398 -1492
rect 224454 -1548 224522 -1492
rect 224578 -1548 224646 -1492
rect 224702 -1548 254994 -1492
rect 255050 -1548 255118 -1492
rect 255174 -1548 255242 -1492
rect 255298 -1548 255366 -1492
rect 255422 -1548 285714 -1492
rect 285770 -1548 285838 -1492
rect 285894 -1548 285962 -1492
rect 286018 -1548 286086 -1492
rect 286142 -1548 316434 -1492
rect 316490 -1548 316558 -1492
rect 316614 -1548 316682 -1492
rect 316738 -1548 316806 -1492
rect 316862 -1548 347154 -1492
rect 347210 -1548 347278 -1492
rect 347334 -1548 347402 -1492
rect 347458 -1548 347526 -1492
rect 347582 -1548 377874 -1492
rect 377930 -1548 377998 -1492
rect 378054 -1548 378122 -1492
rect 378178 -1548 378246 -1492
rect 378302 -1548 408594 -1492
rect 408650 -1548 408718 -1492
rect 408774 -1548 408842 -1492
rect 408898 -1548 408966 -1492
rect 409022 -1548 439314 -1492
rect 439370 -1548 439438 -1492
rect 439494 -1548 439562 -1492
rect 439618 -1548 439686 -1492
rect 439742 -1548 470034 -1492
rect 470090 -1548 470158 -1492
rect 470214 -1548 470282 -1492
rect 470338 -1548 470406 -1492
rect 470462 -1548 500754 -1492
rect 500810 -1548 500878 -1492
rect 500934 -1548 501002 -1492
rect 501058 -1548 501126 -1492
rect 501182 -1548 531474 -1492
rect 531530 -1548 531598 -1492
rect 531654 -1548 531722 -1492
rect 531778 -1548 531846 -1492
rect 531902 -1548 562194 -1492
rect 562250 -1548 562318 -1492
rect 562374 -1548 562442 -1492
rect 562498 -1548 562566 -1492
rect 562622 -1548 592914 -1492
rect 592970 -1548 593038 -1492
rect 593094 -1548 593162 -1492
rect 593218 -1548 593286 -1492
rect 593342 -1548 597456 -1492
rect 597512 -1548 597580 -1492
rect 597636 -1548 597704 -1492
rect 597760 -1548 597828 -1492
rect 597884 -1548 597980 -1492
rect -1916 -1644 597980 -1548
use micro_irritating_maze  micro_irritating_maze
timestamp 0
transform 1 0 12000 0 1 3000
box 0 0 112000 69552
<< labels >>
flabel metal3 s 595560 7112 597000 7336 0 FreeSans 896 0 0 0 io_in[0]
port 0 nsew signal input
flabel metal3 s 595560 403592 597000 403816 0 FreeSans 896 0 0 0 io_in[10]
port 1 nsew signal input
flabel metal3 s 595560 443240 597000 443464 0 FreeSans 896 0 0 0 io_in[11]
port 2 nsew signal input
flabel metal3 s 595560 482888 597000 483112 0 FreeSans 896 0 0 0 io_in[12]
port 3 nsew signal input
flabel metal3 s 595560 522536 597000 522760 0 FreeSans 896 0 0 0 io_in[13]
port 4 nsew signal input
flabel metal3 s 595560 562184 597000 562408 0 FreeSans 896 0 0 0 io_in[14]
port 5 nsew signal input
flabel metal2 s 584696 595560 584920 597000 0 FreeSans 896 90 0 0 io_in[15]
port 6 nsew signal input
flabel metal2 s 518504 595560 518728 597000 0 FreeSans 896 90 0 0 io_in[16]
port 7 nsew signal input
flabel metal2 s 452312 595560 452536 597000 0 FreeSans 896 90 0 0 io_in[17]
port 8 nsew signal input
flabel metal2 s 386120 595560 386344 597000 0 FreeSans 896 90 0 0 io_in[18]
port 9 nsew signal input
flabel metal2 s 319928 595560 320152 597000 0 FreeSans 896 90 0 0 io_in[19]
port 10 nsew signal input
flabel metal3 s 595560 46760 597000 46984 0 FreeSans 896 0 0 0 io_in[1]
port 11 nsew signal input
flabel metal2 s 253736 595560 253960 597000 0 FreeSans 896 90 0 0 io_in[20]
port 12 nsew signal input
flabel metal2 s 187544 595560 187768 597000 0 FreeSans 896 90 0 0 io_in[21]
port 13 nsew signal input
flabel metal2 s 121352 595560 121576 597000 0 FreeSans 896 90 0 0 io_in[22]
port 14 nsew signal input
flabel metal2 s 55160 595560 55384 597000 0 FreeSans 896 90 0 0 io_in[23]
port 15 nsew signal input
flabel metal3 s -960 587160 480 587384 0 FreeSans 896 0 0 0 io_in[24]
port 16 nsew signal input
flabel metal3 s -960 544824 480 545048 0 FreeSans 896 0 0 0 io_in[25]
port 17 nsew signal input
flabel metal3 s -960 502488 480 502712 0 FreeSans 896 0 0 0 io_in[26]
port 18 nsew signal input
flabel metal3 s -960 460152 480 460376 0 FreeSans 896 0 0 0 io_in[27]
port 19 nsew signal input
flabel metal3 s -960 417816 480 418040 0 FreeSans 896 0 0 0 io_in[28]
port 20 nsew signal input
flabel metal3 s -960 375480 480 375704 0 FreeSans 896 0 0 0 io_in[29]
port 21 nsew signal input
flabel metal3 s 595560 86408 597000 86632 0 FreeSans 896 0 0 0 io_in[2]
port 22 nsew signal input
flabel metal3 s -960 333144 480 333368 0 FreeSans 896 0 0 0 io_in[30]
port 23 nsew signal input
flabel metal3 s -960 290808 480 291032 0 FreeSans 896 0 0 0 io_in[31]
port 24 nsew signal input
flabel metal3 s -960 248472 480 248696 0 FreeSans 896 0 0 0 io_in[32]
port 25 nsew signal input
flabel metal3 s -960 206136 480 206360 0 FreeSans 896 0 0 0 io_in[33]
port 26 nsew signal input
flabel metal3 s -960 163800 480 164024 0 FreeSans 896 0 0 0 io_in[34]
port 27 nsew signal input
flabel metal3 s -960 121464 480 121688 0 FreeSans 896 0 0 0 io_in[35]
port 28 nsew signal input
flabel metal3 s -960 79128 480 79352 0 FreeSans 896 0 0 0 io_in[36]
port 29 nsew signal input
flabel metal3 s -960 36792 480 37016 0 FreeSans 896 0 0 0 io_in[37]
port 30 nsew signal input
flabel metal3 s 595560 126056 597000 126280 0 FreeSans 896 0 0 0 io_in[3]
port 31 nsew signal input
flabel metal3 s 595560 165704 597000 165928 0 FreeSans 896 0 0 0 io_in[4]
port 32 nsew signal input
flabel metal3 s 595560 205352 597000 205576 0 FreeSans 896 0 0 0 io_in[5]
port 33 nsew signal input
flabel metal3 s 595560 245000 597000 245224 0 FreeSans 896 0 0 0 io_in[6]
port 34 nsew signal input
flabel metal3 s 595560 284648 597000 284872 0 FreeSans 896 0 0 0 io_in[7]
port 35 nsew signal input
flabel metal3 s 595560 324296 597000 324520 0 FreeSans 896 0 0 0 io_in[8]
port 36 nsew signal input
flabel metal3 s 595560 363944 597000 364168 0 FreeSans 896 0 0 0 io_in[9]
port 37 nsew signal input
flabel metal3 s 595560 33544 597000 33768 0 FreeSans 896 0 0 0 io_oeb[0]
port 38 nsew signal tristate
flabel metal3 s 595560 430024 597000 430248 0 FreeSans 896 0 0 0 io_oeb[10]
port 39 nsew signal tristate
flabel metal3 s 595560 469672 597000 469896 0 FreeSans 896 0 0 0 io_oeb[11]
port 40 nsew signal tristate
flabel metal3 s 595560 509320 597000 509544 0 FreeSans 896 0 0 0 io_oeb[12]
port 41 nsew signal tristate
flabel metal3 s 595560 548968 597000 549192 0 FreeSans 896 0 0 0 io_oeb[13]
port 42 nsew signal tristate
flabel metal3 s 595560 588616 597000 588840 0 FreeSans 896 0 0 0 io_oeb[14]
port 43 nsew signal tristate
flabel metal2 s 540568 595560 540792 597000 0 FreeSans 896 90 0 0 io_oeb[15]
port 44 nsew signal tristate
flabel metal2 s 474376 595560 474600 597000 0 FreeSans 896 90 0 0 io_oeb[16]
port 45 nsew signal tristate
flabel metal2 s 408184 595560 408408 597000 0 FreeSans 896 90 0 0 io_oeb[17]
port 46 nsew signal tristate
flabel metal2 s 341992 595560 342216 597000 0 FreeSans 896 90 0 0 io_oeb[18]
port 47 nsew signal tristate
flabel metal2 s 275800 595560 276024 597000 0 FreeSans 896 90 0 0 io_oeb[19]
port 48 nsew signal tristate
flabel metal3 s 595560 73192 597000 73416 0 FreeSans 896 0 0 0 io_oeb[1]
port 49 nsew signal tristate
flabel metal2 s 209608 595560 209832 597000 0 FreeSans 896 90 0 0 io_oeb[20]
port 50 nsew signal tristate
flabel metal2 s 143416 595560 143640 597000 0 FreeSans 896 90 0 0 io_oeb[21]
port 51 nsew signal tristate
flabel metal2 s 77224 595560 77448 597000 0 FreeSans 896 90 0 0 io_oeb[22]
port 52 nsew signal tristate
flabel metal2 s 11032 595560 11256 597000 0 FreeSans 896 90 0 0 io_oeb[23]
port 53 nsew signal tristate
flabel metal3 s -960 558936 480 559160 0 FreeSans 896 0 0 0 io_oeb[24]
port 54 nsew signal tristate
flabel metal3 s -960 516600 480 516824 0 FreeSans 896 0 0 0 io_oeb[25]
port 55 nsew signal tristate
flabel metal3 s -960 474264 480 474488 0 FreeSans 896 0 0 0 io_oeb[26]
port 56 nsew signal tristate
flabel metal3 s -960 431928 480 432152 0 FreeSans 896 0 0 0 io_oeb[27]
port 57 nsew signal tristate
flabel metal3 s -960 389592 480 389816 0 FreeSans 896 0 0 0 io_oeb[28]
port 58 nsew signal tristate
flabel metal3 s -960 347256 480 347480 0 FreeSans 896 0 0 0 io_oeb[29]
port 59 nsew signal tristate
flabel metal3 s 595560 112840 597000 113064 0 FreeSans 896 0 0 0 io_oeb[2]
port 60 nsew signal tristate
flabel metal3 s -960 304920 480 305144 0 FreeSans 896 0 0 0 io_oeb[30]
port 61 nsew signal tristate
flabel metal3 s -960 262584 480 262808 0 FreeSans 896 0 0 0 io_oeb[31]
port 62 nsew signal tristate
flabel metal3 s -960 220248 480 220472 0 FreeSans 896 0 0 0 io_oeb[32]
port 63 nsew signal tristate
flabel metal3 s -960 177912 480 178136 0 FreeSans 896 0 0 0 io_oeb[33]
port 64 nsew signal tristate
flabel metal3 s -960 135576 480 135800 0 FreeSans 896 0 0 0 io_oeb[34]
port 65 nsew signal tristate
flabel metal3 s -960 93240 480 93464 0 FreeSans 896 0 0 0 io_oeb[35]
port 66 nsew signal tristate
flabel metal3 s -960 50904 480 51128 0 FreeSans 896 0 0 0 io_oeb[36]
port 67 nsew signal tristate
flabel metal3 s -960 8568 480 8792 0 FreeSans 896 0 0 0 io_oeb[37]
port 68 nsew signal tristate
flabel metal3 s 595560 152488 597000 152712 0 FreeSans 896 0 0 0 io_oeb[3]
port 69 nsew signal tristate
flabel metal3 s 595560 192136 597000 192360 0 FreeSans 896 0 0 0 io_oeb[4]
port 70 nsew signal tristate
flabel metal3 s 595560 231784 597000 232008 0 FreeSans 896 0 0 0 io_oeb[5]
port 71 nsew signal tristate
flabel metal3 s 595560 271432 597000 271656 0 FreeSans 896 0 0 0 io_oeb[6]
port 72 nsew signal tristate
flabel metal3 s 595560 311080 597000 311304 0 FreeSans 896 0 0 0 io_oeb[7]
port 73 nsew signal tristate
flabel metal3 s 595560 350728 597000 350952 0 FreeSans 896 0 0 0 io_oeb[8]
port 74 nsew signal tristate
flabel metal3 s 595560 390376 597000 390600 0 FreeSans 896 0 0 0 io_oeb[9]
port 75 nsew signal tristate
flabel metal3 s 595560 20328 597000 20552 0 FreeSans 896 0 0 0 io_out[0]
port 76 nsew signal tristate
flabel metal3 s 595560 416808 597000 417032 0 FreeSans 896 0 0 0 io_out[10]
port 77 nsew signal tristate
flabel metal3 s 595560 456456 597000 456680 0 FreeSans 896 0 0 0 io_out[11]
port 78 nsew signal tristate
flabel metal3 s 595560 496104 597000 496328 0 FreeSans 896 0 0 0 io_out[12]
port 79 nsew signal tristate
flabel metal3 s 595560 535752 597000 535976 0 FreeSans 896 0 0 0 io_out[13]
port 80 nsew signal tristate
flabel metal3 s 595560 575400 597000 575624 0 FreeSans 896 0 0 0 io_out[14]
port 81 nsew signal tristate
flabel metal2 s 562632 595560 562856 597000 0 FreeSans 896 90 0 0 io_out[15]
port 82 nsew signal tristate
flabel metal2 s 496440 595560 496664 597000 0 FreeSans 896 90 0 0 io_out[16]
port 83 nsew signal tristate
flabel metal2 s 430248 595560 430472 597000 0 FreeSans 896 90 0 0 io_out[17]
port 84 nsew signal tristate
flabel metal2 s 364056 595560 364280 597000 0 FreeSans 896 90 0 0 io_out[18]
port 85 nsew signal tristate
flabel metal2 s 297864 595560 298088 597000 0 FreeSans 896 90 0 0 io_out[19]
port 86 nsew signal tristate
flabel metal3 s 595560 59976 597000 60200 0 FreeSans 896 0 0 0 io_out[1]
port 87 nsew signal tristate
flabel metal2 s 231672 595560 231896 597000 0 FreeSans 896 90 0 0 io_out[20]
port 88 nsew signal tristate
flabel metal2 s 165480 595560 165704 597000 0 FreeSans 896 90 0 0 io_out[21]
port 89 nsew signal tristate
flabel metal2 s 99288 595560 99512 597000 0 FreeSans 896 90 0 0 io_out[22]
port 90 nsew signal tristate
flabel metal2 s 33096 595560 33320 597000 0 FreeSans 896 90 0 0 io_out[23]
port 91 nsew signal tristate
flabel metal3 s -960 573048 480 573272 0 FreeSans 896 0 0 0 io_out[24]
port 92 nsew signal tristate
flabel metal3 s -960 530712 480 530936 0 FreeSans 896 0 0 0 io_out[25]
port 93 nsew signal tristate
flabel metal3 s -960 488376 480 488600 0 FreeSans 896 0 0 0 io_out[26]
port 94 nsew signal tristate
flabel metal3 s -960 446040 480 446264 0 FreeSans 896 0 0 0 io_out[27]
port 95 nsew signal tristate
flabel metal3 s -960 403704 480 403928 0 FreeSans 896 0 0 0 io_out[28]
port 96 nsew signal tristate
flabel metal3 s -960 361368 480 361592 0 FreeSans 896 0 0 0 io_out[29]
port 97 nsew signal tristate
flabel metal3 s 595560 99624 597000 99848 0 FreeSans 896 0 0 0 io_out[2]
port 98 nsew signal tristate
flabel metal3 s -960 319032 480 319256 0 FreeSans 896 0 0 0 io_out[30]
port 99 nsew signal tristate
flabel metal3 s -960 276696 480 276920 0 FreeSans 896 0 0 0 io_out[31]
port 100 nsew signal tristate
flabel metal3 s -960 234360 480 234584 0 FreeSans 896 0 0 0 io_out[32]
port 101 nsew signal tristate
flabel metal3 s -960 192024 480 192248 0 FreeSans 896 0 0 0 io_out[33]
port 102 nsew signal tristate
flabel metal3 s -960 149688 480 149912 0 FreeSans 896 0 0 0 io_out[34]
port 103 nsew signal tristate
flabel metal3 s -960 107352 480 107576 0 FreeSans 896 0 0 0 io_out[35]
port 104 nsew signal tristate
flabel metal3 s -960 65016 480 65240 0 FreeSans 896 0 0 0 io_out[36]
port 105 nsew signal tristate
flabel metal3 s -960 22680 480 22904 0 FreeSans 896 0 0 0 io_out[37]
port 106 nsew signal tristate
flabel metal3 s 595560 139272 597000 139496 0 FreeSans 896 0 0 0 io_out[3]
port 107 nsew signal tristate
flabel metal3 s 595560 178920 597000 179144 0 FreeSans 896 0 0 0 io_out[4]
port 108 nsew signal tristate
flabel metal3 s 595560 218568 597000 218792 0 FreeSans 896 0 0 0 io_out[5]
port 109 nsew signal tristate
flabel metal3 s 595560 258216 597000 258440 0 FreeSans 896 0 0 0 io_out[6]
port 110 nsew signal tristate
flabel metal3 s 595560 297864 597000 298088 0 FreeSans 896 0 0 0 io_out[7]
port 111 nsew signal tristate
flabel metal3 s 595560 337512 597000 337736 0 FreeSans 896 0 0 0 io_out[8]
port 112 nsew signal tristate
flabel metal3 s 595560 377160 597000 377384 0 FreeSans 896 0 0 0 io_out[9]
port 113 nsew signal tristate
flabel metal2 s 213192 -960 213416 480 0 FreeSans 896 90 0 0 la_data_in[0]
port 114 nsew signal input
flabel metal2 s 270312 -960 270536 480 0 FreeSans 896 90 0 0 la_data_in[10]
port 115 nsew signal input
flabel metal2 s 276024 -960 276248 480 0 FreeSans 896 90 0 0 la_data_in[11]
port 116 nsew signal input
flabel metal2 s 281736 -960 281960 480 0 FreeSans 896 90 0 0 la_data_in[12]
port 117 nsew signal input
flabel metal2 s 287448 -960 287672 480 0 FreeSans 896 90 0 0 la_data_in[13]
port 118 nsew signal input
flabel metal2 s 293160 -960 293384 480 0 FreeSans 896 90 0 0 la_data_in[14]
port 119 nsew signal input
flabel metal2 s 298872 -960 299096 480 0 FreeSans 896 90 0 0 la_data_in[15]
port 120 nsew signal input
flabel metal2 s 304584 -960 304808 480 0 FreeSans 896 90 0 0 la_data_in[16]
port 121 nsew signal input
flabel metal2 s 310296 -960 310520 480 0 FreeSans 896 90 0 0 la_data_in[17]
port 122 nsew signal input
flabel metal2 s 316008 -960 316232 480 0 FreeSans 896 90 0 0 la_data_in[18]
port 123 nsew signal input
flabel metal2 s 321720 -960 321944 480 0 FreeSans 896 90 0 0 la_data_in[19]
port 124 nsew signal input
flabel metal2 s 218904 -960 219128 480 0 FreeSans 896 90 0 0 la_data_in[1]
port 125 nsew signal input
flabel metal2 s 327432 -960 327656 480 0 FreeSans 896 90 0 0 la_data_in[20]
port 126 nsew signal input
flabel metal2 s 333144 -960 333368 480 0 FreeSans 896 90 0 0 la_data_in[21]
port 127 nsew signal input
flabel metal2 s 338856 -960 339080 480 0 FreeSans 896 90 0 0 la_data_in[22]
port 128 nsew signal input
flabel metal2 s 344568 -960 344792 480 0 FreeSans 896 90 0 0 la_data_in[23]
port 129 nsew signal input
flabel metal2 s 350280 -960 350504 480 0 FreeSans 896 90 0 0 la_data_in[24]
port 130 nsew signal input
flabel metal2 s 355992 -960 356216 480 0 FreeSans 896 90 0 0 la_data_in[25]
port 131 nsew signal input
flabel metal2 s 361704 -960 361928 480 0 FreeSans 896 90 0 0 la_data_in[26]
port 132 nsew signal input
flabel metal2 s 367416 -960 367640 480 0 FreeSans 896 90 0 0 la_data_in[27]
port 133 nsew signal input
flabel metal2 s 373128 -960 373352 480 0 FreeSans 896 90 0 0 la_data_in[28]
port 134 nsew signal input
flabel metal2 s 378840 -960 379064 480 0 FreeSans 896 90 0 0 la_data_in[29]
port 135 nsew signal input
flabel metal2 s 224616 -960 224840 480 0 FreeSans 896 90 0 0 la_data_in[2]
port 136 nsew signal input
flabel metal2 s 384552 -960 384776 480 0 FreeSans 896 90 0 0 la_data_in[30]
port 137 nsew signal input
flabel metal2 s 390264 -960 390488 480 0 FreeSans 896 90 0 0 la_data_in[31]
port 138 nsew signal input
flabel metal2 s 395976 -960 396200 480 0 FreeSans 896 90 0 0 la_data_in[32]
port 139 nsew signal input
flabel metal2 s 401688 -960 401912 480 0 FreeSans 896 90 0 0 la_data_in[33]
port 140 nsew signal input
flabel metal2 s 407400 -960 407624 480 0 FreeSans 896 90 0 0 la_data_in[34]
port 141 nsew signal input
flabel metal2 s 413112 -960 413336 480 0 FreeSans 896 90 0 0 la_data_in[35]
port 142 nsew signal input
flabel metal2 s 418824 -960 419048 480 0 FreeSans 896 90 0 0 la_data_in[36]
port 143 nsew signal input
flabel metal2 s 424536 -960 424760 480 0 FreeSans 896 90 0 0 la_data_in[37]
port 144 nsew signal input
flabel metal2 s 430248 -960 430472 480 0 FreeSans 896 90 0 0 la_data_in[38]
port 145 nsew signal input
flabel metal2 s 435960 -960 436184 480 0 FreeSans 896 90 0 0 la_data_in[39]
port 146 nsew signal input
flabel metal2 s 230328 -960 230552 480 0 FreeSans 896 90 0 0 la_data_in[3]
port 147 nsew signal input
flabel metal2 s 441672 -960 441896 480 0 FreeSans 896 90 0 0 la_data_in[40]
port 148 nsew signal input
flabel metal2 s 447384 -960 447608 480 0 FreeSans 896 90 0 0 la_data_in[41]
port 149 nsew signal input
flabel metal2 s 453096 -960 453320 480 0 FreeSans 896 90 0 0 la_data_in[42]
port 150 nsew signal input
flabel metal2 s 458808 -960 459032 480 0 FreeSans 896 90 0 0 la_data_in[43]
port 151 nsew signal input
flabel metal2 s 464520 -960 464744 480 0 FreeSans 896 90 0 0 la_data_in[44]
port 152 nsew signal input
flabel metal2 s 470232 -960 470456 480 0 FreeSans 896 90 0 0 la_data_in[45]
port 153 nsew signal input
flabel metal2 s 475944 -960 476168 480 0 FreeSans 896 90 0 0 la_data_in[46]
port 154 nsew signal input
flabel metal2 s 481656 -960 481880 480 0 FreeSans 896 90 0 0 la_data_in[47]
port 155 nsew signal input
flabel metal2 s 487368 -960 487592 480 0 FreeSans 896 90 0 0 la_data_in[48]
port 156 nsew signal input
flabel metal2 s 493080 -960 493304 480 0 FreeSans 896 90 0 0 la_data_in[49]
port 157 nsew signal input
flabel metal2 s 236040 -960 236264 480 0 FreeSans 896 90 0 0 la_data_in[4]
port 158 nsew signal input
flabel metal2 s 498792 -960 499016 480 0 FreeSans 896 90 0 0 la_data_in[50]
port 159 nsew signal input
flabel metal2 s 504504 -960 504728 480 0 FreeSans 896 90 0 0 la_data_in[51]
port 160 nsew signal input
flabel metal2 s 510216 -960 510440 480 0 FreeSans 896 90 0 0 la_data_in[52]
port 161 nsew signal input
flabel metal2 s 515928 -960 516152 480 0 FreeSans 896 90 0 0 la_data_in[53]
port 162 nsew signal input
flabel metal2 s 521640 -960 521864 480 0 FreeSans 896 90 0 0 la_data_in[54]
port 163 nsew signal input
flabel metal2 s 527352 -960 527576 480 0 FreeSans 896 90 0 0 la_data_in[55]
port 164 nsew signal input
flabel metal2 s 533064 -960 533288 480 0 FreeSans 896 90 0 0 la_data_in[56]
port 165 nsew signal input
flabel metal2 s 538776 -960 539000 480 0 FreeSans 896 90 0 0 la_data_in[57]
port 166 nsew signal input
flabel metal2 s 544488 -960 544712 480 0 FreeSans 896 90 0 0 la_data_in[58]
port 167 nsew signal input
flabel metal2 s 550200 -960 550424 480 0 FreeSans 896 90 0 0 la_data_in[59]
port 168 nsew signal input
flabel metal2 s 241752 -960 241976 480 0 FreeSans 896 90 0 0 la_data_in[5]
port 169 nsew signal input
flabel metal2 s 555912 -960 556136 480 0 FreeSans 896 90 0 0 la_data_in[60]
port 170 nsew signal input
flabel metal2 s 561624 -960 561848 480 0 FreeSans 896 90 0 0 la_data_in[61]
port 171 nsew signal input
flabel metal2 s 567336 -960 567560 480 0 FreeSans 896 90 0 0 la_data_in[62]
port 172 nsew signal input
flabel metal2 s 573048 -960 573272 480 0 FreeSans 896 90 0 0 la_data_in[63]
port 173 nsew signal input
flabel metal2 s 247464 -960 247688 480 0 FreeSans 896 90 0 0 la_data_in[6]
port 174 nsew signal input
flabel metal2 s 253176 -960 253400 480 0 FreeSans 896 90 0 0 la_data_in[7]
port 175 nsew signal input
flabel metal2 s 258888 -960 259112 480 0 FreeSans 896 90 0 0 la_data_in[8]
port 176 nsew signal input
flabel metal2 s 264600 -960 264824 480 0 FreeSans 896 90 0 0 la_data_in[9]
port 177 nsew signal input
flabel metal2 s 215096 -960 215320 480 0 FreeSans 896 90 0 0 la_data_out[0]
port 178 nsew signal tristate
flabel metal2 s 272216 -960 272440 480 0 FreeSans 896 90 0 0 la_data_out[10]
port 179 nsew signal tristate
flabel metal2 s 277928 -960 278152 480 0 FreeSans 896 90 0 0 la_data_out[11]
port 180 nsew signal tristate
flabel metal2 s 283640 -960 283864 480 0 FreeSans 896 90 0 0 la_data_out[12]
port 181 nsew signal tristate
flabel metal2 s 289352 -960 289576 480 0 FreeSans 896 90 0 0 la_data_out[13]
port 182 nsew signal tristate
flabel metal2 s 295064 -960 295288 480 0 FreeSans 896 90 0 0 la_data_out[14]
port 183 nsew signal tristate
flabel metal2 s 300776 -960 301000 480 0 FreeSans 896 90 0 0 la_data_out[15]
port 184 nsew signal tristate
flabel metal2 s 306488 -960 306712 480 0 FreeSans 896 90 0 0 la_data_out[16]
port 185 nsew signal tristate
flabel metal2 s 312200 -960 312424 480 0 FreeSans 896 90 0 0 la_data_out[17]
port 186 nsew signal tristate
flabel metal2 s 317912 -960 318136 480 0 FreeSans 896 90 0 0 la_data_out[18]
port 187 nsew signal tristate
flabel metal2 s 323624 -960 323848 480 0 FreeSans 896 90 0 0 la_data_out[19]
port 188 nsew signal tristate
flabel metal2 s 220808 -960 221032 480 0 FreeSans 896 90 0 0 la_data_out[1]
port 189 nsew signal tristate
flabel metal2 s 329336 -960 329560 480 0 FreeSans 896 90 0 0 la_data_out[20]
port 190 nsew signal tristate
flabel metal2 s 335048 -960 335272 480 0 FreeSans 896 90 0 0 la_data_out[21]
port 191 nsew signal tristate
flabel metal2 s 340760 -960 340984 480 0 FreeSans 896 90 0 0 la_data_out[22]
port 192 nsew signal tristate
flabel metal2 s 346472 -960 346696 480 0 FreeSans 896 90 0 0 la_data_out[23]
port 193 nsew signal tristate
flabel metal2 s 352184 -960 352408 480 0 FreeSans 896 90 0 0 la_data_out[24]
port 194 nsew signal tristate
flabel metal2 s 357896 -960 358120 480 0 FreeSans 896 90 0 0 la_data_out[25]
port 195 nsew signal tristate
flabel metal2 s 363608 -960 363832 480 0 FreeSans 896 90 0 0 la_data_out[26]
port 196 nsew signal tristate
flabel metal2 s 369320 -960 369544 480 0 FreeSans 896 90 0 0 la_data_out[27]
port 197 nsew signal tristate
flabel metal2 s 375032 -960 375256 480 0 FreeSans 896 90 0 0 la_data_out[28]
port 198 nsew signal tristate
flabel metal2 s 380744 -960 380968 480 0 FreeSans 896 90 0 0 la_data_out[29]
port 199 nsew signal tristate
flabel metal2 s 226520 -960 226744 480 0 FreeSans 896 90 0 0 la_data_out[2]
port 200 nsew signal tristate
flabel metal2 s 386456 -960 386680 480 0 FreeSans 896 90 0 0 la_data_out[30]
port 201 nsew signal tristate
flabel metal2 s 392168 -960 392392 480 0 FreeSans 896 90 0 0 la_data_out[31]
port 202 nsew signal tristate
flabel metal2 s 397880 -960 398104 480 0 FreeSans 896 90 0 0 la_data_out[32]
port 203 nsew signal tristate
flabel metal2 s 403592 -960 403816 480 0 FreeSans 896 90 0 0 la_data_out[33]
port 204 nsew signal tristate
flabel metal2 s 409304 -960 409528 480 0 FreeSans 896 90 0 0 la_data_out[34]
port 205 nsew signal tristate
flabel metal2 s 415016 -960 415240 480 0 FreeSans 896 90 0 0 la_data_out[35]
port 206 nsew signal tristate
flabel metal2 s 420728 -960 420952 480 0 FreeSans 896 90 0 0 la_data_out[36]
port 207 nsew signal tristate
flabel metal2 s 426440 -960 426664 480 0 FreeSans 896 90 0 0 la_data_out[37]
port 208 nsew signal tristate
flabel metal2 s 432152 -960 432376 480 0 FreeSans 896 90 0 0 la_data_out[38]
port 209 nsew signal tristate
flabel metal2 s 437864 -960 438088 480 0 FreeSans 896 90 0 0 la_data_out[39]
port 210 nsew signal tristate
flabel metal2 s 232232 -960 232456 480 0 FreeSans 896 90 0 0 la_data_out[3]
port 211 nsew signal tristate
flabel metal2 s 443576 -960 443800 480 0 FreeSans 896 90 0 0 la_data_out[40]
port 212 nsew signal tristate
flabel metal2 s 449288 -960 449512 480 0 FreeSans 896 90 0 0 la_data_out[41]
port 213 nsew signal tristate
flabel metal2 s 455000 -960 455224 480 0 FreeSans 896 90 0 0 la_data_out[42]
port 214 nsew signal tristate
flabel metal2 s 460712 -960 460936 480 0 FreeSans 896 90 0 0 la_data_out[43]
port 215 nsew signal tristate
flabel metal2 s 466424 -960 466648 480 0 FreeSans 896 90 0 0 la_data_out[44]
port 216 nsew signal tristate
flabel metal2 s 472136 -960 472360 480 0 FreeSans 896 90 0 0 la_data_out[45]
port 217 nsew signal tristate
flabel metal2 s 477848 -960 478072 480 0 FreeSans 896 90 0 0 la_data_out[46]
port 218 nsew signal tristate
flabel metal2 s 483560 -960 483784 480 0 FreeSans 896 90 0 0 la_data_out[47]
port 219 nsew signal tristate
flabel metal2 s 489272 -960 489496 480 0 FreeSans 896 90 0 0 la_data_out[48]
port 220 nsew signal tristate
flabel metal2 s 494984 -960 495208 480 0 FreeSans 896 90 0 0 la_data_out[49]
port 221 nsew signal tristate
flabel metal2 s 237944 -960 238168 480 0 FreeSans 896 90 0 0 la_data_out[4]
port 222 nsew signal tristate
flabel metal2 s 500696 -960 500920 480 0 FreeSans 896 90 0 0 la_data_out[50]
port 223 nsew signal tristate
flabel metal2 s 506408 -960 506632 480 0 FreeSans 896 90 0 0 la_data_out[51]
port 224 nsew signal tristate
flabel metal2 s 512120 -960 512344 480 0 FreeSans 896 90 0 0 la_data_out[52]
port 225 nsew signal tristate
flabel metal2 s 517832 -960 518056 480 0 FreeSans 896 90 0 0 la_data_out[53]
port 226 nsew signal tristate
flabel metal2 s 523544 -960 523768 480 0 FreeSans 896 90 0 0 la_data_out[54]
port 227 nsew signal tristate
flabel metal2 s 529256 -960 529480 480 0 FreeSans 896 90 0 0 la_data_out[55]
port 228 nsew signal tristate
flabel metal2 s 534968 -960 535192 480 0 FreeSans 896 90 0 0 la_data_out[56]
port 229 nsew signal tristate
flabel metal2 s 540680 -960 540904 480 0 FreeSans 896 90 0 0 la_data_out[57]
port 230 nsew signal tristate
flabel metal2 s 546392 -960 546616 480 0 FreeSans 896 90 0 0 la_data_out[58]
port 231 nsew signal tristate
flabel metal2 s 552104 -960 552328 480 0 FreeSans 896 90 0 0 la_data_out[59]
port 232 nsew signal tristate
flabel metal2 s 243656 -960 243880 480 0 FreeSans 896 90 0 0 la_data_out[5]
port 233 nsew signal tristate
flabel metal2 s 557816 -960 558040 480 0 FreeSans 896 90 0 0 la_data_out[60]
port 234 nsew signal tristate
flabel metal2 s 563528 -960 563752 480 0 FreeSans 896 90 0 0 la_data_out[61]
port 235 nsew signal tristate
flabel metal2 s 569240 -960 569464 480 0 FreeSans 896 90 0 0 la_data_out[62]
port 236 nsew signal tristate
flabel metal2 s 574952 -960 575176 480 0 FreeSans 896 90 0 0 la_data_out[63]
port 237 nsew signal tristate
flabel metal2 s 249368 -960 249592 480 0 FreeSans 896 90 0 0 la_data_out[6]
port 238 nsew signal tristate
flabel metal2 s 255080 -960 255304 480 0 FreeSans 896 90 0 0 la_data_out[7]
port 239 nsew signal tristate
flabel metal2 s 260792 -960 261016 480 0 FreeSans 896 90 0 0 la_data_out[8]
port 240 nsew signal tristate
flabel metal2 s 266504 -960 266728 480 0 FreeSans 896 90 0 0 la_data_out[9]
port 241 nsew signal tristate
flabel metal2 s 217000 -960 217224 480 0 FreeSans 896 90 0 0 la_oenb[0]
port 242 nsew signal input
flabel metal2 s 274120 -960 274344 480 0 FreeSans 896 90 0 0 la_oenb[10]
port 243 nsew signal input
flabel metal2 s 279832 -960 280056 480 0 FreeSans 896 90 0 0 la_oenb[11]
port 244 nsew signal input
flabel metal2 s 285544 -960 285768 480 0 FreeSans 896 90 0 0 la_oenb[12]
port 245 nsew signal input
flabel metal2 s 291256 -960 291480 480 0 FreeSans 896 90 0 0 la_oenb[13]
port 246 nsew signal input
flabel metal2 s 296968 -960 297192 480 0 FreeSans 896 90 0 0 la_oenb[14]
port 247 nsew signal input
flabel metal2 s 302680 -960 302904 480 0 FreeSans 896 90 0 0 la_oenb[15]
port 248 nsew signal input
flabel metal2 s 308392 -960 308616 480 0 FreeSans 896 90 0 0 la_oenb[16]
port 249 nsew signal input
flabel metal2 s 314104 -960 314328 480 0 FreeSans 896 90 0 0 la_oenb[17]
port 250 nsew signal input
flabel metal2 s 319816 -960 320040 480 0 FreeSans 896 90 0 0 la_oenb[18]
port 251 nsew signal input
flabel metal2 s 325528 -960 325752 480 0 FreeSans 896 90 0 0 la_oenb[19]
port 252 nsew signal input
flabel metal2 s 222712 -960 222936 480 0 FreeSans 896 90 0 0 la_oenb[1]
port 253 nsew signal input
flabel metal2 s 331240 -960 331464 480 0 FreeSans 896 90 0 0 la_oenb[20]
port 254 nsew signal input
flabel metal2 s 336952 -960 337176 480 0 FreeSans 896 90 0 0 la_oenb[21]
port 255 nsew signal input
flabel metal2 s 342664 -960 342888 480 0 FreeSans 896 90 0 0 la_oenb[22]
port 256 nsew signal input
flabel metal2 s 348376 -960 348600 480 0 FreeSans 896 90 0 0 la_oenb[23]
port 257 nsew signal input
flabel metal2 s 354088 -960 354312 480 0 FreeSans 896 90 0 0 la_oenb[24]
port 258 nsew signal input
flabel metal2 s 359800 -960 360024 480 0 FreeSans 896 90 0 0 la_oenb[25]
port 259 nsew signal input
flabel metal2 s 365512 -960 365736 480 0 FreeSans 896 90 0 0 la_oenb[26]
port 260 nsew signal input
flabel metal2 s 371224 -960 371448 480 0 FreeSans 896 90 0 0 la_oenb[27]
port 261 nsew signal input
flabel metal2 s 376936 -960 377160 480 0 FreeSans 896 90 0 0 la_oenb[28]
port 262 nsew signal input
flabel metal2 s 382648 -960 382872 480 0 FreeSans 896 90 0 0 la_oenb[29]
port 263 nsew signal input
flabel metal2 s 228424 -960 228648 480 0 FreeSans 896 90 0 0 la_oenb[2]
port 264 nsew signal input
flabel metal2 s 388360 -960 388584 480 0 FreeSans 896 90 0 0 la_oenb[30]
port 265 nsew signal input
flabel metal2 s 394072 -960 394296 480 0 FreeSans 896 90 0 0 la_oenb[31]
port 266 nsew signal input
flabel metal2 s 399784 -960 400008 480 0 FreeSans 896 90 0 0 la_oenb[32]
port 267 nsew signal input
flabel metal2 s 405496 -960 405720 480 0 FreeSans 896 90 0 0 la_oenb[33]
port 268 nsew signal input
flabel metal2 s 411208 -960 411432 480 0 FreeSans 896 90 0 0 la_oenb[34]
port 269 nsew signal input
flabel metal2 s 416920 -960 417144 480 0 FreeSans 896 90 0 0 la_oenb[35]
port 270 nsew signal input
flabel metal2 s 422632 -960 422856 480 0 FreeSans 896 90 0 0 la_oenb[36]
port 271 nsew signal input
flabel metal2 s 428344 -960 428568 480 0 FreeSans 896 90 0 0 la_oenb[37]
port 272 nsew signal input
flabel metal2 s 434056 -960 434280 480 0 FreeSans 896 90 0 0 la_oenb[38]
port 273 nsew signal input
flabel metal2 s 439768 -960 439992 480 0 FreeSans 896 90 0 0 la_oenb[39]
port 274 nsew signal input
flabel metal2 s 234136 -960 234360 480 0 FreeSans 896 90 0 0 la_oenb[3]
port 275 nsew signal input
flabel metal2 s 445480 -960 445704 480 0 FreeSans 896 90 0 0 la_oenb[40]
port 276 nsew signal input
flabel metal2 s 451192 -960 451416 480 0 FreeSans 896 90 0 0 la_oenb[41]
port 277 nsew signal input
flabel metal2 s 456904 -960 457128 480 0 FreeSans 896 90 0 0 la_oenb[42]
port 278 nsew signal input
flabel metal2 s 462616 -960 462840 480 0 FreeSans 896 90 0 0 la_oenb[43]
port 279 nsew signal input
flabel metal2 s 468328 -960 468552 480 0 FreeSans 896 90 0 0 la_oenb[44]
port 280 nsew signal input
flabel metal2 s 474040 -960 474264 480 0 FreeSans 896 90 0 0 la_oenb[45]
port 281 nsew signal input
flabel metal2 s 479752 -960 479976 480 0 FreeSans 896 90 0 0 la_oenb[46]
port 282 nsew signal input
flabel metal2 s 485464 -960 485688 480 0 FreeSans 896 90 0 0 la_oenb[47]
port 283 nsew signal input
flabel metal2 s 491176 -960 491400 480 0 FreeSans 896 90 0 0 la_oenb[48]
port 284 nsew signal input
flabel metal2 s 496888 -960 497112 480 0 FreeSans 896 90 0 0 la_oenb[49]
port 285 nsew signal input
flabel metal2 s 239848 -960 240072 480 0 FreeSans 896 90 0 0 la_oenb[4]
port 286 nsew signal input
flabel metal2 s 502600 -960 502824 480 0 FreeSans 896 90 0 0 la_oenb[50]
port 287 nsew signal input
flabel metal2 s 508312 -960 508536 480 0 FreeSans 896 90 0 0 la_oenb[51]
port 288 nsew signal input
flabel metal2 s 514024 -960 514248 480 0 FreeSans 896 90 0 0 la_oenb[52]
port 289 nsew signal input
flabel metal2 s 519736 -960 519960 480 0 FreeSans 896 90 0 0 la_oenb[53]
port 290 nsew signal input
flabel metal2 s 525448 -960 525672 480 0 FreeSans 896 90 0 0 la_oenb[54]
port 291 nsew signal input
flabel metal2 s 531160 -960 531384 480 0 FreeSans 896 90 0 0 la_oenb[55]
port 292 nsew signal input
flabel metal2 s 536872 -960 537096 480 0 FreeSans 896 90 0 0 la_oenb[56]
port 293 nsew signal input
flabel metal2 s 542584 -960 542808 480 0 FreeSans 896 90 0 0 la_oenb[57]
port 294 nsew signal input
flabel metal2 s 548296 -960 548520 480 0 FreeSans 896 90 0 0 la_oenb[58]
port 295 nsew signal input
flabel metal2 s 554008 -960 554232 480 0 FreeSans 896 90 0 0 la_oenb[59]
port 296 nsew signal input
flabel metal2 s 245560 -960 245784 480 0 FreeSans 896 90 0 0 la_oenb[5]
port 297 nsew signal input
flabel metal2 s 559720 -960 559944 480 0 FreeSans 896 90 0 0 la_oenb[60]
port 298 nsew signal input
flabel metal2 s 565432 -960 565656 480 0 FreeSans 896 90 0 0 la_oenb[61]
port 299 nsew signal input
flabel metal2 s 571144 -960 571368 480 0 FreeSans 896 90 0 0 la_oenb[62]
port 300 nsew signal input
flabel metal2 s 576856 -960 577080 480 0 FreeSans 896 90 0 0 la_oenb[63]
port 301 nsew signal input
flabel metal2 s 251272 -960 251496 480 0 FreeSans 896 90 0 0 la_oenb[6]
port 302 nsew signal input
flabel metal2 s 256984 -960 257208 480 0 FreeSans 896 90 0 0 la_oenb[7]
port 303 nsew signal input
flabel metal2 s 262696 -960 262920 480 0 FreeSans 896 90 0 0 la_oenb[8]
port 304 nsew signal input
flabel metal2 s 268408 -960 268632 480 0 FreeSans 896 90 0 0 la_oenb[9]
port 305 nsew signal input
flabel metal2 s 578760 -960 578984 480 0 FreeSans 896 90 0 0 user_clock2
port 306 nsew signal input
flabel metal2 s 580664 -960 580888 480 0 FreeSans 896 90 0 0 user_irq[0]
port 307 nsew signal tristate
flabel metal2 s 582568 -960 582792 480 0 FreeSans 896 90 0 0 user_irq[1]
port 308 nsew signal tristate
flabel metal2 s 584472 -960 584696 480 0 FreeSans 896 90 0 0 user_irq[2]
port 309 nsew signal tristate
flabel metal4 s -956 -684 -336 597308 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -956 -684 597020 -64 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -956 596688 597020 597308 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 596400 -684 597020 597308 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 5418 -1644 6038 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 36138 -1644 36758 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 66858 -1644 67478 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 97578 -1644 98198 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 128298 -1644 128918 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 159018 -1644 159638 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 189738 -1644 190358 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 220458 -1644 221078 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 251178 -1644 251798 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 281898 -1644 282518 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 312618 -1644 313238 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 343338 -1644 343958 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 374058 -1644 374678 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 404778 -1644 405398 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 435498 -1644 436118 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 466218 -1644 466838 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 496938 -1644 497558 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 527658 -1644 528278 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 558378 -1644 558998 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 589098 -1644 589718 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 3826 597980 4446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 21826 597980 22446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 39826 597980 40446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 57826 597980 58446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 75826 597980 76446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 93826 597980 94446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 111826 597980 112446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 129826 597980 130446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 147826 597980 148446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 165826 597980 166446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 183826 597980 184446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 201826 597980 202446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 219826 597980 220446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 237826 597980 238446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 255826 597980 256446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 273826 597980 274446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 291826 597980 292446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 309826 597980 310446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 327826 597980 328446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 345826 597980 346446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 363826 597980 364446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 381826 597980 382446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 399826 597980 400446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 417826 597980 418446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 435826 597980 436446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 453826 597980 454446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 471826 597980 472446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 489826 597980 490446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 507826 597980 508446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 525826 597980 526446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 543826 597980 544446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 561826 597980 562446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 579826 597980 580446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s -1916 -1644 -1296 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 -1644 597980 -1024 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 597648 597980 598268 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 597360 -1644 597980 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 9138 -1644 9758 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 39858 -1644 40478 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 70578 -1644 71198 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 101298 -1644 101918 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 132018 -1644 132638 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 162738 -1644 163358 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 193458 -1644 194078 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 224178 -1644 224798 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 254898 -1644 255518 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 285618 -1644 286238 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 316338 -1644 316958 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 347058 -1644 347678 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 377778 -1644 378398 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 408498 -1644 409118 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 439218 -1644 439838 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 469938 -1644 470558 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 500658 -1644 501278 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 531378 -1644 531998 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 562098 -1644 562718 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 592818 -1644 593438 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 9826 597980 10446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 27826 597980 28446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 45826 597980 46446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 63826 597980 64446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 81826 597980 82446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 99826 597980 100446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 117826 597980 118446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 135826 597980 136446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 153826 597980 154446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 171826 597980 172446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 189826 597980 190446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 207826 597980 208446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 225826 597980 226446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 243826 597980 244446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 261826 597980 262446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 279826 597980 280446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 297826 597980 298446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 315826 597980 316446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 333826 597980 334446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 351826 597980 352446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 369826 597980 370446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 387826 597980 388446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 405826 597980 406446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 423826 597980 424446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 441826 597980 442446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 459826 597980 460446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 477826 597980 478446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 495826 597980 496446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 513826 597980 514446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 531826 597980 532446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 549826 597980 550446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 567826 597980 568446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 585826 597980 586446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal2 s 11368 -960 11592 480 0 FreeSans 896 90 0 0 wb_clk_i
port 312 nsew signal input
flabel metal2 s 13272 -960 13496 480 0 FreeSans 896 90 0 0 wb_rst_i
port 313 nsew signal input
flabel metal2 s 15176 -960 15400 480 0 FreeSans 896 90 0 0 wbs_ack_o
port 314 nsew signal tristate
flabel metal2 s 22792 -960 23016 480 0 FreeSans 896 90 0 0 wbs_adr_i[0]
port 315 nsew signal input
flabel metal2 s 87528 -960 87752 480 0 FreeSans 896 90 0 0 wbs_adr_i[10]
port 316 nsew signal input
flabel metal2 s 93240 -960 93464 480 0 FreeSans 896 90 0 0 wbs_adr_i[11]
port 317 nsew signal input
flabel metal2 s 98952 -960 99176 480 0 FreeSans 896 90 0 0 wbs_adr_i[12]
port 318 nsew signal input
flabel metal2 s 104664 -960 104888 480 0 FreeSans 896 90 0 0 wbs_adr_i[13]
port 319 nsew signal input
flabel metal2 s 110376 -960 110600 480 0 FreeSans 896 90 0 0 wbs_adr_i[14]
port 320 nsew signal input
flabel metal2 s 116088 -960 116312 480 0 FreeSans 896 90 0 0 wbs_adr_i[15]
port 321 nsew signal input
flabel metal2 s 121800 -960 122024 480 0 FreeSans 896 90 0 0 wbs_adr_i[16]
port 322 nsew signal input
flabel metal2 s 127512 -960 127736 480 0 FreeSans 896 90 0 0 wbs_adr_i[17]
port 323 nsew signal input
flabel metal2 s 133224 -960 133448 480 0 FreeSans 896 90 0 0 wbs_adr_i[18]
port 324 nsew signal input
flabel metal2 s 138936 -960 139160 480 0 FreeSans 896 90 0 0 wbs_adr_i[19]
port 325 nsew signal input
flabel metal2 s 30408 -960 30632 480 0 FreeSans 896 90 0 0 wbs_adr_i[1]
port 326 nsew signal input
flabel metal2 s 144648 -960 144872 480 0 FreeSans 896 90 0 0 wbs_adr_i[20]
port 327 nsew signal input
flabel metal2 s 150360 -960 150584 480 0 FreeSans 896 90 0 0 wbs_adr_i[21]
port 328 nsew signal input
flabel metal2 s 156072 -960 156296 480 0 FreeSans 896 90 0 0 wbs_adr_i[22]
port 329 nsew signal input
flabel metal2 s 161784 -960 162008 480 0 FreeSans 896 90 0 0 wbs_adr_i[23]
port 330 nsew signal input
flabel metal2 s 167496 -960 167720 480 0 FreeSans 896 90 0 0 wbs_adr_i[24]
port 331 nsew signal input
flabel metal2 s 173208 -960 173432 480 0 FreeSans 896 90 0 0 wbs_adr_i[25]
port 332 nsew signal input
flabel metal2 s 178920 -960 179144 480 0 FreeSans 896 90 0 0 wbs_adr_i[26]
port 333 nsew signal input
flabel metal2 s 184632 -960 184856 480 0 FreeSans 896 90 0 0 wbs_adr_i[27]
port 334 nsew signal input
flabel metal2 s 190344 -960 190568 480 0 FreeSans 896 90 0 0 wbs_adr_i[28]
port 335 nsew signal input
flabel metal2 s 196056 -960 196280 480 0 FreeSans 896 90 0 0 wbs_adr_i[29]
port 336 nsew signal input
flabel metal2 s 38024 -960 38248 480 0 FreeSans 896 90 0 0 wbs_adr_i[2]
port 337 nsew signal input
flabel metal2 s 201768 -960 201992 480 0 FreeSans 896 90 0 0 wbs_adr_i[30]
port 338 nsew signal input
flabel metal2 s 207480 -960 207704 480 0 FreeSans 896 90 0 0 wbs_adr_i[31]
port 339 nsew signal input
flabel metal2 s 45640 -960 45864 480 0 FreeSans 896 90 0 0 wbs_adr_i[3]
port 340 nsew signal input
flabel metal2 s 53256 -960 53480 480 0 FreeSans 896 90 0 0 wbs_adr_i[4]
port 341 nsew signal input
flabel metal2 s 58968 -960 59192 480 0 FreeSans 896 90 0 0 wbs_adr_i[5]
port 342 nsew signal input
flabel metal2 s 64680 -960 64904 480 0 FreeSans 896 90 0 0 wbs_adr_i[6]
port 343 nsew signal input
flabel metal2 s 70392 -960 70616 480 0 FreeSans 896 90 0 0 wbs_adr_i[7]
port 344 nsew signal input
flabel metal2 s 76104 -960 76328 480 0 FreeSans 896 90 0 0 wbs_adr_i[8]
port 345 nsew signal input
flabel metal2 s 81816 -960 82040 480 0 FreeSans 896 90 0 0 wbs_adr_i[9]
port 346 nsew signal input
flabel metal2 s 17080 -960 17304 480 0 FreeSans 896 90 0 0 wbs_cyc_i
port 347 nsew signal input
flabel metal2 s 24696 -960 24920 480 0 FreeSans 896 90 0 0 wbs_dat_i[0]
port 348 nsew signal input
flabel metal2 s 89432 -960 89656 480 0 FreeSans 896 90 0 0 wbs_dat_i[10]
port 349 nsew signal input
flabel metal2 s 95144 -960 95368 480 0 FreeSans 896 90 0 0 wbs_dat_i[11]
port 350 nsew signal input
flabel metal2 s 100856 -960 101080 480 0 FreeSans 896 90 0 0 wbs_dat_i[12]
port 351 nsew signal input
flabel metal2 s 106568 -960 106792 480 0 FreeSans 896 90 0 0 wbs_dat_i[13]
port 352 nsew signal input
flabel metal2 s 112280 -960 112504 480 0 FreeSans 896 90 0 0 wbs_dat_i[14]
port 353 nsew signal input
flabel metal2 s 117992 -960 118216 480 0 FreeSans 896 90 0 0 wbs_dat_i[15]
port 354 nsew signal input
flabel metal2 s 123704 -960 123928 480 0 FreeSans 896 90 0 0 wbs_dat_i[16]
port 355 nsew signal input
flabel metal2 s 129416 -960 129640 480 0 FreeSans 896 90 0 0 wbs_dat_i[17]
port 356 nsew signal input
flabel metal2 s 135128 -960 135352 480 0 FreeSans 896 90 0 0 wbs_dat_i[18]
port 357 nsew signal input
flabel metal2 s 140840 -960 141064 480 0 FreeSans 896 90 0 0 wbs_dat_i[19]
port 358 nsew signal input
flabel metal2 s 32312 -960 32536 480 0 FreeSans 896 90 0 0 wbs_dat_i[1]
port 359 nsew signal input
flabel metal2 s 146552 -960 146776 480 0 FreeSans 896 90 0 0 wbs_dat_i[20]
port 360 nsew signal input
flabel metal2 s 152264 -960 152488 480 0 FreeSans 896 90 0 0 wbs_dat_i[21]
port 361 nsew signal input
flabel metal2 s 157976 -960 158200 480 0 FreeSans 896 90 0 0 wbs_dat_i[22]
port 362 nsew signal input
flabel metal2 s 163688 -960 163912 480 0 FreeSans 896 90 0 0 wbs_dat_i[23]
port 363 nsew signal input
flabel metal2 s 169400 -960 169624 480 0 FreeSans 896 90 0 0 wbs_dat_i[24]
port 364 nsew signal input
flabel metal2 s 175112 -960 175336 480 0 FreeSans 896 90 0 0 wbs_dat_i[25]
port 365 nsew signal input
flabel metal2 s 180824 -960 181048 480 0 FreeSans 896 90 0 0 wbs_dat_i[26]
port 366 nsew signal input
flabel metal2 s 186536 -960 186760 480 0 FreeSans 896 90 0 0 wbs_dat_i[27]
port 367 nsew signal input
flabel metal2 s 192248 -960 192472 480 0 FreeSans 896 90 0 0 wbs_dat_i[28]
port 368 nsew signal input
flabel metal2 s 197960 -960 198184 480 0 FreeSans 896 90 0 0 wbs_dat_i[29]
port 369 nsew signal input
flabel metal2 s 39928 -960 40152 480 0 FreeSans 896 90 0 0 wbs_dat_i[2]
port 370 nsew signal input
flabel metal2 s 203672 -960 203896 480 0 FreeSans 896 90 0 0 wbs_dat_i[30]
port 371 nsew signal input
flabel metal2 s 209384 -960 209608 480 0 FreeSans 896 90 0 0 wbs_dat_i[31]
port 372 nsew signal input
flabel metal2 s 47544 -960 47768 480 0 FreeSans 896 90 0 0 wbs_dat_i[3]
port 373 nsew signal input
flabel metal2 s 55160 -960 55384 480 0 FreeSans 896 90 0 0 wbs_dat_i[4]
port 374 nsew signal input
flabel metal2 s 60872 -960 61096 480 0 FreeSans 896 90 0 0 wbs_dat_i[5]
port 375 nsew signal input
flabel metal2 s 66584 -960 66808 480 0 FreeSans 896 90 0 0 wbs_dat_i[6]
port 376 nsew signal input
flabel metal2 s 72296 -960 72520 480 0 FreeSans 896 90 0 0 wbs_dat_i[7]
port 377 nsew signal input
flabel metal2 s 78008 -960 78232 480 0 FreeSans 896 90 0 0 wbs_dat_i[8]
port 378 nsew signal input
flabel metal2 s 83720 -960 83944 480 0 FreeSans 896 90 0 0 wbs_dat_i[9]
port 379 nsew signal input
flabel metal2 s 26600 -960 26824 480 0 FreeSans 896 90 0 0 wbs_dat_o[0]
port 380 nsew signal tristate
flabel metal2 s 91336 -960 91560 480 0 FreeSans 896 90 0 0 wbs_dat_o[10]
port 381 nsew signal tristate
flabel metal2 s 97048 -960 97272 480 0 FreeSans 896 90 0 0 wbs_dat_o[11]
port 382 nsew signal tristate
flabel metal2 s 102760 -960 102984 480 0 FreeSans 896 90 0 0 wbs_dat_o[12]
port 383 nsew signal tristate
flabel metal2 s 108472 -960 108696 480 0 FreeSans 896 90 0 0 wbs_dat_o[13]
port 384 nsew signal tristate
flabel metal2 s 114184 -960 114408 480 0 FreeSans 896 90 0 0 wbs_dat_o[14]
port 385 nsew signal tristate
flabel metal2 s 119896 -960 120120 480 0 FreeSans 896 90 0 0 wbs_dat_o[15]
port 386 nsew signal tristate
flabel metal2 s 125608 -960 125832 480 0 FreeSans 896 90 0 0 wbs_dat_o[16]
port 387 nsew signal tristate
flabel metal2 s 131320 -960 131544 480 0 FreeSans 896 90 0 0 wbs_dat_o[17]
port 388 nsew signal tristate
flabel metal2 s 137032 -960 137256 480 0 FreeSans 896 90 0 0 wbs_dat_o[18]
port 389 nsew signal tristate
flabel metal2 s 142744 -960 142968 480 0 FreeSans 896 90 0 0 wbs_dat_o[19]
port 390 nsew signal tristate
flabel metal2 s 34216 -960 34440 480 0 FreeSans 896 90 0 0 wbs_dat_o[1]
port 391 nsew signal tristate
flabel metal2 s 148456 -960 148680 480 0 FreeSans 896 90 0 0 wbs_dat_o[20]
port 392 nsew signal tristate
flabel metal2 s 154168 -960 154392 480 0 FreeSans 896 90 0 0 wbs_dat_o[21]
port 393 nsew signal tristate
flabel metal2 s 159880 -960 160104 480 0 FreeSans 896 90 0 0 wbs_dat_o[22]
port 394 nsew signal tristate
flabel metal2 s 165592 -960 165816 480 0 FreeSans 896 90 0 0 wbs_dat_o[23]
port 395 nsew signal tristate
flabel metal2 s 171304 -960 171528 480 0 FreeSans 896 90 0 0 wbs_dat_o[24]
port 396 nsew signal tristate
flabel metal2 s 177016 -960 177240 480 0 FreeSans 896 90 0 0 wbs_dat_o[25]
port 397 nsew signal tristate
flabel metal2 s 182728 -960 182952 480 0 FreeSans 896 90 0 0 wbs_dat_o[26]
port 398 nsew signal tristate
flabel metal2 s 188440 -960 188664 480 0 FreeSans 896 90 0 0 wbs_dat_o[27]
port 399 nsew signal tristate
flabel metal2 s 194152 -960 194376 480 0 FreeSans 896 90 0 0 wbs_dat_o[28]
port 400 nsew signal tristate
flabel metal2 s 199864 -960 200088 480 0 FreeSans 896 90 0 0 wbs_dat_o[29]
port 401 nsew signal tristate
flabel metal2 s 41832 -960 42056 480 0 FreeSans 896 90 0 0 wbs_dat_o[2]
port 402 nsew signal tristate
flabel metal2 s 205576 -960 205800 480 0 FreeSans 896 90 0 0 wbs_dat_o[30]
port 403 nsew signal tristate
flabel metal2 s 211288 -960 211512 480 0 FreeSans 896 90 0 0 wbs_dat_o[31]
port 404 nsew signal tristate
flabel metal2 s 49448 -960 49672 480 0 FreeSans 896 90 0 0 wbs_dat_o[3]
port 405 nsew signal tristate
flabel metal2 s 57064 -960 57288 480 0 FreeSans 896 90 0 0 wbs_dat_o[4]
port 406 nsew signal tristate
flabel metal2 s 62776 -960 63000 480 0 FreeSans 896 90 0 0 wbs_dat_o[5]
port 407 nsew signal tristate
flabel metal2 s 68488 -960 68712 480 0 FreeSans 896 90 0 0 wbs_dat_o[6]
port 408 nsew signal tristate
flabel metal2 s 74200 -960 74424 480 0 FreeSans 896 90 0 0 wbs_dat_o[7]
port 409 nsew signal tristate
flabel metal2 s 79912 -960 80136 480 0 FreeSans 896 90 0 0 wbs_dat_o[8]
port 410 nsew signal tristate
flabel metal2 s 85624 -960 85848 480 0 FreeSans 896 90 0 0 wbs_dat_o[9]
port 411 nsew signal tristate
flabel metal2 s 28504 -960 28728 480 0 FreeSans 896 90 0 0 wbs_sel_i[0]
port 412 nsew signal input
flabel metal2 s 36120 -960 36344 480 0 FreeSans 896 90 0 0 wbs_sel_i[1]
port 413 nsew signal input
flabel metal2 s 43736 -960 43960 480 0 FreeSans 896 90 0 0 wbs_sel_i[2]
port 414 nsew signal input
flabel metal2 s 51352 -960 51576 480 0 FreeSans 896 90 0 0 wbs_sel_i[3]
port 415 nsew signal input
flabel metal2 s 18984 -960 19208 480 0 FreeSans 896 90 0 0 wbs_stb_i
port 416 nsew signal input
flabel metal2 s 20888 -960 21112 480 0 FreeSans 896 90 0 0 wbs_we_i
port 417 nsew signal input
rlabel via4 108830 58322 108830 58322 0 vdd
rlabel via4 101794 64322 101794 64322 0 vss
rlabel metal3 125454 5544 125454 5544 0 io_in[0]
rlabel metal4 8232 234472 8232 234472 0 io_in[10]
rlabel metal3 12488 63014 12488 63014 0 io_in[11]
rlabel metal4 8344 271432 8344 271432 0 io_in[12]
rlabel metal3 593082 522536 593082 522536 0 io_in[13]
rlabel metal3 593194 562184 593194 562184 0 io_in[14]
rlabel metal2 584696 593082 584696 593082 0 io_in[15]
rlabel metal2 8008 67032 8008 67032 0 io_in[16]
rlabel metal2 452312 341922 452312 341922 0 io_in[17]
rlabel metal2 8232 66864 8232 66864 0 io_in[18]
rlabel metal2 8344 66360 8344 66360 0 io_in[19]
rlabel metal3 593082 46760 593082 46760 0 io_in[1]
rlabel metal2 1624 311136 1624 311136 0 io_in[20]
rlabel metal3 187040 590184 187040 590184 0 io_in[21]
rlabel metal3 121184 590184 121184 590184 0 io_in[22]
rlabel metal2 55160 334362 55160 334362 0 io_in[23]
rlabel metal3 1918 587160 1918 587160 0 io_in[24]
rlabel metal3 280 544712 280 544712 0 io_in[25]
rlabel metal3 1470 502488 1470 502488 0 io_in[26]
rlabel metal3 3990 460152 3990 460152 0 io_in[27]
rlabel metal3 392 417704 392 417704 0 io_in[28]
rlabel metal3 1526 375480 1526 375480 0 io_in[29]
rlabel metal3 125678 23016 125678 23016 0 io_in[2]
rlabel metal3 518 333144 518 333144 0 io_in[30]
rlabel metal3 4046 290808 4046 290808 0 io_in[31]
rlabel metal3 126518 31752 126518 31752 0 io_in[3]
rlabel metal4 590184 164752 590184 164752 0 io_in[4]
rlabel metal3 129598 49224 129598 49224 0 io_in[5]
rlabel metal3 593474 245000 593474 245000 0 io_in[6]
rlabel metal3 384762 284648 384762 284648 0 io_in[7]
rlabel metal4 47880 202888 47880 202888 0 io_in[8]
rlabel metal3 591402 363944 591402 363944 0 io_in[9]
rlabel metal3 125510 11368 125510 11368 0 io_oeb[0]
rlabel metal3 303674 430136 303674 430136 0 io_oeb[10]
rlabel metal2 22680 271544 22680 271544 0 io_oeb[11]
rlabel metal3 12600 58478 12600 58478 0 io_oeb[12]
rlabel metal4 24360 302969 24360 302969 0 io_oeb[13]
rlabel metal4 26040 321623 26040 321623 0 io_oeb[14]
rlabel metal2 540568 346122 540568 346122 0 io_oeb[15]
rlabel metal2 474376 346962 474376 346962 0 io_oeb[16]
rlabel metal4 27720 320111 27720 320111 0 io_oeb[17]
rlabel metal4 6552 60943 6552 60943 0 io_oeb[18]
rlabel metal3 143920 101640 143920 101640 0 io_oeb[19]
rlabel metal3 128856 30296 128856 30296 0 io_oeb[1]
rlabel metal2 1512 61600 1512 61600 0 io_oeb[20]
rlabel metal2 3304 60312 3304 60312 0 io_oeb[21]
rlabel metal2 8120 53088 8120 53088 0 io_oeb[22]
rlabel metal3 11522 28616 11522 28616 0 io_oeb[23]
rlabel metal3 11466 25928 11466 25928 0 io_oeb[24]
rlabel metal4 11984 26550 11984 26550 0 io_oeb[25]
rlabel metal3 336 474152 336 474152 0 io_oeb[26]
rlabel metal3 2310 431928 2310 431928 0 io_oeb[27]
rlabel metal3 2366 389592 2366 389592 0 io_oeb[28]
rlabel metal3 1582 347256 1582 347256 0 io_oeb[29]
rlabel metal4 138600 70840 138600 70840 0 io_oeb[2]
rlabel metal3 2422 304920 2422 304920 0 io_oeb[30]
rlabel metal3 2534 262584 2534 262584 0 io_oeb[31]
rlabel metal4 140280 95032 140280 95032 0 io_oeb[3]
rlabel metal4 141960 120008 141960 120008 0 io_oeb[4]
rlabel metal4 148680 143472 148680 143472 0 io_oeb[5]
rlabel metal4 145320 167608 145320 167608 0 io_oeb[6]
rlabel metal3 125398 72520 125398 72520 0 io_oeb[7]
rlabel metal4 12712 68983 12712 68983 0 io_oeb[8]
rlabel metal4 29400 228713 29400 228713 0 io_oeb[9]
rlabel metal3 591402 20552 591402 20552 0 io_out[0]
rlabel metal4 76440 241119 76440 241119 0 io_out[10]
rlabel metal4 21000 259233 21000 259233 0 io_out[11]
rlabel metal4 590184 495432 590184 495432 0 io_out[12]
rlabel metal3 22176 73304 22176 73304 0 io_out[13]
rlabel via4 12712 53717 12712 53717 0 io_out[14]
rlabel metal4 22680 317025 22680 317025 0 io_out[15]
rlabel metal2 496440 587202 496440 587202 0 io_out[16]
rlabel metal2 430248 349482 430248 349482 0 io_out[17]
rlabel metal2 4872 63056 4872 63056 0 io_out[18]
rlabel metal4 6664 59237 6664 59237 0 io_out[19]
rlabel metal3 125398 17192 125398 17192 0 io_out[1]
rlabel metal2 4984 61264 4984 61264 0 io_out[20]
rlabel metal3 165088 590184 165088 590184 0 io_out[21]
rlabel metal2 99288 592914 99288 592914 0 io_out[22]
rlabel metal2 6664 51352 6664 51352 0 io_out[23]
rlabel metal4 12040 29372 12040 29372 0 io_out[24]
rlabel metal3 10514 24136 10514 24136 0 io_out[25]
rlabel metal3 10458 21448 10458 21448 0 io_out[26]
rlabel metal3 2534 446040 2534 446040 0 io_out[27]
rlabel metal3 11088 72968 11088 72968 0 io_out[28]
rlabel metal3 5488 275576 5488 275576 0 io_out[29]
rlabel metal4 590184 98952 590184 98952 0 io_out[2]
rlabel metal3 10304 73976 10304 73976 0 io_out[30]
rlabel metal3 2478 276696 2478 276696 0 io_out[31]
rlabel metal3 361466 139272 361466 139272 0 io_out[3]
rlabel metal3 125566 43400 125566 43400 0 io_out[4]
rlabel metal3 125510 52136 125510 52136 0 io_out[5]
rlabel metal3 361298 258216 361298 258216 0 io_out[6]
rlabel metal4 590184 297192 590184 297192 0 io_out[7]
rlabel metal4 21112 206136 21112 206136 0 io_out[8]
rlabel metal2 46200 226800 46200 226800 0 io_out[9]
rlabel metal2 213192 36918 213192 36918 0 la_data_in[0]
rlabel metal3 167832 74648 167832 74648 0 la_data_in[10]
rlabel metal2 65800 2282 65800 2282 0 la_data_in[11]
rlabel metal2 281736 37478 281736 37478 0 la_data_in[12]
rlabel metal2 287448 36694 287448 36694 0 la_data_in[13]
rlabel metal3 180488 74424 180488 74424 0 la_data_in[14]
rlabel metal3 183848 72744 183848 72744 0 la_data_in[15]
rlabel metal2 304584 37366 304584 37366 0 la_data_in[16]
rlabel metal2 310296 39326 310296 39326 0 la_data_in[17]
rlabel metal3 193200 80696 193200 80696 0 la_data_in[18]
rlabel metal3 196728 78120 196728 78120 0 la_data_in[19]
rlabel metal2 218904 38430 218904 38430 0 la_data_in[1]
rlabel metal5 74312 25110 74312 25110 0 la_data_in[20]
rlabel metal2 333144 38262 333144 38262 0 la_data_in[21]
rlabel metal3 73976 3192 73976 3192 0 la_data_in[22]
rlabel metal3 209216 75992 209216 75992 0 la_data_in[23]
rlabel metal2 350280 39102 350280 39102 0 la_data_in[24]
rlabel metal3 75152 3192 75152 3192 0 la_data_in[25]
rlabel metal3 218792 79576 218792 79576 0 la_data_in[26]
rlabel metal3 222264 74088 222264 74088 0 la_data_in[27]
rlabel metal5 77672 21690 77672 21690 0 la_data_in[28]
rlabel metal2 378840 39830 378840 39830 0 la_data_in[29]
rlabel metal4 53704 31950 53704 31950 0 la_data_in[2]
rlabel metal3 383824 4200 383824 4200 0 la_data_in[30]
rlabel metal3 234864 77672 234864 77672 0 la_data_in[31]
rlabel metal3 395416 4200 395416 4200 0 la_data_in[32]
rlabel metal2 401688 38094 401688 38094 0 la_data_in[33]
rlabel metal3 407008 4200 407008 4200 0 la_data_in[34]
rlabel metal4 81928 20160 81928 20160 0 la_data_in[35]
rlabel metal3 250712 74872 250712 74872 0 la_data_in[36]
rlabel metal2 424536 38990 424536 38990 0 la_data_in[37]
rlabel metal2 430248 40166 430248 40166 0 la_data_in[38]
rlabel metal3 435568 4200 435568 4200 0 la_data_in[39]
rlabel metal3 145376 76328 145376 76328 0 la_data_in[3]
rlabel metal3 263648 77448 263648 77448 0 la_data_in[40]
rlabel metal3 447160 4200 447160 4200 0 la_data_in[41]
rlabel metal3 452536 4200 452536 4200 0 la_data_in[42]
rlabel metal2 458808 2310 458808 2310 0 la_data_in[43]
rlabel metal3 276248 76552 276248 76552 0 la_data_in[44]
rlabel metal3 469504 4200 469504 4200 0 la_data_in[45]
rlabel metal3 475720 4200 475720 4200 0 la_data_in[46]
rlabel metal3 481096 4200 481096 4200 0 la_data_in[47]
rlabel metal2 487368 2310 487368 2310 0 la_data_in[48]
rlabel metal3 492688 4200 492688 4200 0 la_data_in[49]
rlabel metal3 235648 4200 235648 4200 0 la_data_in[4]
rlabel metal3 498232 4200 498232 4200 0 la_data_in[50]
rlabel metal3 93240 3192 93240 3192 0 la_data_in[51]
rlabel metal3 509656 4200 509656 4200 0 la_data_in[52]
rlabel metal3 93464 3304 93464 3304 0 la_data_in[53]
rlabel metal3 95144 3304 95144 3304 0 la_data_in[54]
rlabel metal3 526624 4200 526624 4200 0 la_data_in[55]
rlabel metal3 532840 4200 532840 4200 0 la_data_in[56]
rlabel metal3 538216 4200 538216 4200 0 la_data_in[57]
rlabel metal2 544488 2310 544488 2310 0 la_data_in[58]
rlabel metal3 98392 3416 98392 3416 0 la_data_in[59]
rlabel metal2 241752 37590 241752 37590 0 la_data_in[5]
rlabel metal3 98672 3752 98672 3752 0 la_data_in[60]
rlabel metal3 561400 4200 561400 4200 0 la_data_in[61]
rlabel metal3 100296 3416 100296 3416 0 la_data_in[62]
rlabel metal3 100688 3752 100688 3752 0 la_data_in[63]
rlabel metal4 52808 38783 52808 38783 0 la_data_in[6]
rlabel metal3 252616 4200 252616 4200 0 la_data_in[7]
rlabel metal2 258888 2310 258888 2310 0 la_data_in[8]
rlabel metal3 264208 4200 264208 4200 0 la_data_in[9]
rlabel metal2 215096 2310 215096 2310 0 la_data_out[0]
rlabel metal3 168840 79800 168840 79800 0 la_data_out[10]
rlabel metal3 167160 72856 167160 72856 0 la_data_out[11]
rlabel metal3 283136 4200 283136 4200 0 la_data_out[12]
rlabel metal3 68040 3192 68040 3192 0 la_data_out[13]
rlabel metal3 67368 3080 67368 3080 0 la_data_out[14]
rlabel metal2 300776 2310 300776 2310 0 la_data_out[15]
rlabel metal3 306152 4200 306152 4200 0 la_data_out[16]
rlabel metal2 70056 2338 70056 2338 0 la_data_out[17]
rlabel metal5 78512 51570 78512 51570 0 la_data_out[18]
rlabel metal2 71400 2898 71400 2898 0 la_data_out[19]
rlabel metal3 220472 4200 220472 4200 0 la_data_out[1]
rlabel metal3 70952 3192 70952 3192 0 la_data_out[20]
rlabel metal2 335048 37310 335048 37310 0 la_data_out[21]
rlabel metal3 340088 4200 340088 4200 0 la_data_out[22]
rlabel metal2 74088 2170 74088 2170 0 la_data_out[23]
rlabel metal3 351680 4200 351680 4200 0 la_data_out[24]
rlabel metal2 357896 38150 357896 38150 0 la_data_out[25]
rlabel metal3 363272 4200 363272 4200 0 la_data_out[26]
rlabel metal3 77616 3192 77616 3192 0 la_data_out[27]
rlabel metal2 375032 2310 375032 2310 0 la_data_out[28]
rlabel metal3 380240 4200 380240 4200 0 la_data_out[29]
rlabel metal3 59248 3304 59248 3304 0 la_data_out[2]
rlabel metal2 78792 1666 78792 1666 0 la_data_out[30]
rlabel metal3 80584 3304 80584 3304 0 la_data_out[31]
rlabel metal3 397208 4200 397208 4200 0 la_data_out[32]
rlabel metal3 403424 4200 403424 4200 0 la_data_out[33]
rlabel metal4 409304 4633 409304 4633 0 la_data_out[34]
rlabel metal4 121016 4755 121016 4755 0 la_data_out[35]
rlabel metal3 420392 4200 420392 4200 0 la_data_out[36]
rlabel metal3 425768 4200 425768 4200 0 la_data_out[37]
rlabel metal3 431984 4200 431984 4200 0 la_data_out[38]
rlabel metal3 437360 4200 437360 4200 0 la_data_out[39]
rlabel metal3 232064 4200 232064 4200 0 la_data_out[3]
rlabel metal2 443576 2310 443576 2310 0 la_data_out[40]
rlabel metal3 448952 4200 448952 4200 0 la_data_out[41]
rlabel metal3 454328 4200 454328 4200 0 la_data_out[42]
rlabel metal3 460544 4200 460544 4200 0 la_data_out[43]
rlabel metal3 465920 4200 465920 4200 0 la_data_out[44]
rlabel metal2 472136 2310 472136 2310 0 la_data_out[45]
rlabel metal3 477512 4200 477512 4200 0 la_data_out[46]
rlabel metal3 482888 4200 482888 4200 0 la_data_out[47]
rlabel metal3 489104 4200 489104 4200 0 la_data_out[48]
rlabel metal3 91896 3304 91896 3304 0 la_data_out[49]
rlabel metal3 237440 4200 237440 4200 0 la_data_out[4]
rlabel metal2 500920 2310 500920 2310 0 la_data_out[50]
rlabel metal3 506072 4200 506072 4200 0 la_data_out[51]
rlabel metal5 94304 15210 94304 15210 0 la_data_out[52]
rlabel metal3 517664 4200 517664 4200 0 la_data_out[53]
rlabel metal3 523040 4200 523040 4200 0 la_data_out[54]
rlabel metal3 95032 3192 95032 3192 0 la_data_out[55]
rlabel metal3 534632 4200 534632 4200 0 la_data_out[56]
rlabel metal3 540008 4200 540008 4200 0 la_data_out[57]
rlabel metal3 98224 3304 98224 3304 0 la_data_out[58]
rlabel metal3 101416 3192 101416 3192 0 la_data_out[59]
rlabel metal3 61880 3752 61880 3752 0 la_data_out[5]
rlabel via4 98952 3171 98952 3171 0 la_data_out[60]
rlabel metal4 99624 5251 99624 5251 0 la_data_out[61]
rlabel metal3 100240 3752 100240 3752 0 la_data_out[62]
rlabel metal3 101696 3752 101696 3752 0 la_data_out[63]
rlabel metal3 63112 3192 63112 3192 0 la_data_out[6]
rlabel metal4 78456 58050 78456 58050 0 la_data_out[7]
rlabel metal3 260624 4200 260624 4200 0 la_data_out[8]
rlabel metal3 266000 4200 266000 4200 0 la_data_out[9]
rlabel metal2 217000 2310 217000 2310 0 la_oenb[0]
rlabel metal4 73192 42930 73192 42930 0 la_oenb[10]
rlabel metal3 279384 4200 279384 4200 0 la_oenb[11]
rlabel metal2 285768 2310 285768 2310 0 la_oenb[12]
rlabel metal3 290976 4200 290976 4200 0 la_oenb[13]
rlabel metal3 68320 3080 68320 3080 0 la_oenb[14]
rlabel metal2 302680 2310 302680 2310 0 la_oenb[15]
rlabel metal2 78904 2016 78904 2016 0 la_oenb[16]
rlabel metal2 314216 2310 314216 2310 0 la_oenb[17]
rlabel metal2 70952 2114 70952 2114 0 la_oenb[18]
rlabel metal3 324912 4200 324912 4200 0 la_oenb[19]
rlabel metal3 222264 4200 222264 4200 0 la_oenb[1]
rlabel metal2 331240 2310 331240 2310 0 la_oenb[20]
rlabel metal3 336504 4200 336504 4200 0 la_oenb[21]
rlabel metal4 104104 28350 104104 28350 0 la_oenb[22]
rlabel metal3 75600 3080 75600 3080 0 la_oenb[23]
rlabel metal3 353472 4200 353472 4200 0 la_oenb[24]
rlabel metal2 75656 2786 75656 2786 0 la_oenb[25]
rlabel metal4 76328 1577 76328 1577 0 la_oenb[26]
rlabel metal2 371336 2310 371336 2310 0 la_oenb[27]
rlabel metal3 376656 4200 376656 4200 0 la_oenb[28]
rlabel metal2 78344 2226 78344 2226 0 la_oenb[29]
rlabel metal2 228536 2310 228536 2310 0 la_oenb[2]
rlabel metal2 79016 2898 79016 2898 0 la_oenb[30]
rlabel metal2 79688 2338 79688 2338 0 la_oenb[31]
rlabel metal2 95704 1960 95704 1960 0 la_oenb[32]
rlabel metal2 405496 1078 405496 1078 0 la_oenb[33]
rlabel metal2 81704 2170 81704 2170 0 la_oenb[34]
rlabel metal4 100072 24030 100072 24030 0 la_oenb[35]
rlabel metal2 422632 2310 422632 2310 0 la_oenb[36]
rlabel metal2 428456 2310 428456 2310 0 la_oenb[37]
rlabel metal3 99064 78680 99064 78680 0 la_oenb[38]
rlabel metal2 85064 2058 85064 2058 0 la_oenb[39]
rlabel metal3 233856 4200 233856 4200 0 la_oenb[3]
rlabel metal2 445480 1470 445480 1470 0 la_oenb[40]
rlabel metal3 450744 4200 450744 4200 0 la_oenb[41]
rlabel metal3 88872 1568 88872 1568 0 la_oenb[42]
rlabel metal2 87752 2114 87752 2114 0 la_oenb[43]
rlabel metal4 468328 5229 468328 5229 0 la_oenb[44]
rlabel metal2 474040 2310 474040 2310 0 la_oenb[45]
rlabel metal2 89768 2282 89768 2282 0 la_oenb[46]
rlabel metal2 95592 2856 95592 2856 0 la_oenb[47]
rlabel metal3 95592 2856 95592 2856 0 la_oenb[48]
rlabel metal2 91784 2338 91784 2338 0 la_oenb[49]
rlabel metal3 239232 4200 239232 4200 0 la_oenb[4]
rlabel metal2 92456 1946 92456 1946 0 la_oenb[50]
rlabel metal2 508312 2310 508312 2310 0 la_oenb[51]
rlabel metal2 93800 2058 93800 2058 0 la_oenb[52]
rlabel metal2 94472 2114 94472 2114 0 la_oenb[53]
rlabel metal3 96264 1344 96264 1344 0 la_oenb[54]
rlabel metal3 96488 3304 96488 3304 0 la_oenb[55]
rlabel metal2 96488 2226 96488 2226 0 la_oenb[56]
rlabel metal2 97384 1120 97384 1120 0 la_oenb[57]
rlabel metal2 97832 2282 97832 2282 0 la_oenb[58]
rlabel metal4 98504 1397 98504 1397 0 la_oenb[59]
rlabel metal3 62832 3080 62832 3080 0 la_oenb[5]
rlabel metal4 99176 1487 99176 1487 0 la_oenb[60]
rlabel metal3 564984 4200 564984 4200 0 la_oenb[61]
rlabel metal4 100520 1577 100520 1577 0 la_oenb[62]
rlabel metal2 101654 3416 101654 3416 0 la_oenb[63]
rlabel metal3 250824 4200 250824 4200 0 la_oenb[6]
rlabel metal4 257096 5319 257096 5319 0 la_oenb[7]
rlabel metal3 262416 4200 262416 4200 0 la_oenb[8]
rlabel metal4 268408 4543 268408 4543 0 la_oenb[9]
rlabel metal2 11592 1918 11592 1918 0 wb_clk_i
rlabel metal2 13384 742 13384 742 0 wb_rst_i
rlabel metal2 15400 1750 15400 1750 0 wbs_ack_o
rlabel metal2 23016 462 23016 462 0 wbs_adr_i[0]
rlabel metal3 43064 3304 43064 3304 0 wbs_adr_i[10]
rlabel metal4 44296 4441 44296 4441 0 wbs_adr_i[11]
rlabel metal4 44968 5791 44968 5791 0 wbs_adr_i[12]
rlabel metal4 45640 7861 45640 7861 0 wbs_adr_i[13]
rlabel metal3 46424 3752 46424 3752 0 wbs_adr_i[14]
rlabel metal3 46872 3528 46872 3528 0 wbs_adr_i[15]
rlabel metal3 121464 3528 121464 3528 0 wbs_adr_i[16]
rlabel metal3 48272 3752 48272 3752 0 wbs_adr_i[17]
rlabel metal4 49000 24151 49000 24151 0 wbs_adr_i[18]
rlabel metal3 49952 3528 49952 3528 0 wbs_adr_i[19]
rlabel metal2 30632 630 30632 630 0 wbs_adr_i[1]
rlabel metal2 144648 2310 144648 2310 0 wbs_adr_i[20]
rlabel metal4 51016 10651 51016 10651 0 wbs_adr_i[21]
rlabel metal3 51856 3528 51856 3528 0 wbs_adr_i[22]
rlabel metal3 161560 4200 161560 4200 0 wbs_adr_i[23]
rlabel metal3 53816 3416 53816 3416 0 wbs_adr_i[24]
rlabel metal3 53592 3752 53592 3752 0 wbs_adr_i[25]
rlabel metal4 54376 18121 54376 18121 0 wbs_adr_i[26]
rlabel metal3 55160 3752 55160 3752 0 wbs_adr_i[27]
rlabel metal2 190456 2310 190456 2310 0 wbs_adr_i[28]
rlabel metal3 195496 4200 195496 4200 0 wbs_adr_i[29]
rlabel metal2 38024 1022 38024 1022 0 wbs_adr_i[2]
rlabel metal3 57008 3752 57008 3752 0 wbs_adr_i[30]
rlabel metal4 94920 63000 94920 63000 0 wbs_adr_i[31]
rlabel metal2 45640 686 45640 686 0 wbs_adr_i[3]
rlabel metal4 53144 3192 53144 3192 0 wbs_adr_i[4]
rlabel metal3 44408 1456 44408 1456 0 wbs_adr_i[5]
rlabel metal4 40936 4621 40936 4621 0 wbs_adr_i[6]
rlabel metal2 70392 1302 70392 1302 0 wbs_adr_i[7]
rlabel metal3 76216 2856 76216 2856 0 wbs_adr_i[8]
rlabel metal2 42952 2730 42952 2730 0 wbs_adr_i[9]
rlabel metal2 17416 336 17416 336 0 wbs_cyc_i
rlabel metal2 24920 518 24920 518 0 wbs_dat_i[0]
rlabel metal4 43848 2935 43848 2935 0 wbs_dat_i[10]
rlabel metal4 49896 1848 49896 1848 0 wbs_dat_i[11]
rlabel metal2 45192 1778 45192 1778 0 wbs_dat_i[12]
rlabel via4 45864 3317 45864 3317 0 wbs_dat_i[13]
rlabel metal3 46760 3416 46760 3416 0 wbs_dat_i[14]
rlabel metal5 52136 1980 52136 1980 0 wbs_dat_i[15]
rlabel metal3 48160 3528 48160 3528 0 wbs_dat_i[16]
rlabel metal4 48552 43120 48552 43120 0 wbs_dat_i[17]
rlabel metal4 73976 49500 73976 49500 0 wbs_dat_i[18]
rlabel metal3 140168 4200 140168 4200 0 wbs_dat_i[19]
rlabel metal2 32536 1974 32536 1974 0 wbs_dat_i[1]
rlabel metal3 146384 4200 146384 4200 0 wbs_dat_i[20]
rlabel metal4 51240 20731 51240 20731 0 wbs_dat_i[21]
rlabel metal3 51856 3752 51856 3752 0 wbs_dat_i[22]
rlabel metal2 52584 2170 52584 2170 0 wbs_dat_i[23]
rlabel metal2 169400 2310 169400 2310 0 wbs_dat_i[24]
rlabel metal4 53928 12181 53928 12181 0 wbs_dat_i[25]
rlabel metal3 54992 3528 54992 3528 0 wbs_dat_i[26]
rlabel metal2 55272 2282 55272 2282 0 wbs_dat_i[27]
rlabel metal3 191912 4200 191912 4200 0 wbs_dat_i[28]
rlabel metal4 56616 3025 56616 3025 0 wbs_dat_i[29]
rlabel metal2 39928 966 39928 966 0 wbs_dat_i[2]
rlabel metal2 203672 2310 203672 2310 0 wbs_dat_i[30]
rlabel metal4 209384 5465 209384 5465 0 wbs_dat_i[31]
rlabel metal4 46312 2856 46312 2856 0 wbs_dat_i[3]
rlabel metal2 55104 840 55104 840 0 wbs_dat_i[4]
rlabel metal2 40488 2842 40488 2842 0 wbs_dat_i[5]
rlabel metal2 41160 2898 41160 2898 0 wbs_dat_i[6]
rlabel metal2 72408 1638 72408 1638 0 wbs_dat_i[7]
rlabel metal4 53816 2851 53816 2851 0 wbs_dat_i[8]
rlabel metal3 83720 2856 83720 2856 0 wbs_dat_i[9]
rlabel metal2 26824 686 26824 686 0 wbs_dat_o[0]
rlabel metal3 54264 1456 54264 1456 0 wbs_dat_o[10]
rlabel metal3 96488 2744 96488 2744 0 wbs_dat_o[11]
rlabel metal2 45416 2114 45416 2114 0 wbs_dat_o[12]
rlabel metal3 46256 3528 46256 3528 0 wbs_dat_o[13]
rlabel metal3 46816 3752 46816 3752 0 wbs_dat_o[14]
rlabel metal3 47880 3416 47880 3416 0 wbs_dat_o[15]
rlabel metal4 48104 1577 48104 1577 0 wbs_dat_o[16]
rlabel metal3 49448 3416 49448 3416 0 wbs_dat_o[17]
rlabel metal3 55272 896 55272 896 0 wbs_dat_o[18]
rlabel metal3 51352 3304 51352 3304 0 wbs_dat_o[19]
rlabel metal2 34440 966 34440 966 0 wbs_dat_o[1]
rlabel metal2 50792 2226 50792 2226 0 wbs_dat_o[20]
rlabel metal3 51688 3416 51688 3416 0 wbs_dat_o[21]
rlabel metal2 52136 1890 52136 1890 0 wbs_dat_o[22]
rlabel metal3 53200 3528 53200 3528 0 wbs_dat_o[23]
rlabel metal4 53480 1307 53480 1307 0 wbs_dat_o[24]
rlabel metal4 54152 3920 54152 3920 0 wbs_dat_o[25]
rlabel metal3 55132 3304 55132 3304 0 wbs_dat_o[26]
rlabel metal2 188440 686 188440 686 0 wbs_dat_o[27]
rlabel metal4 193256 3463 193256 3463 0 wbs_dat_o[28]
rlabel metal3 61880 336 61880 336 0 wbs_dat_o[29]
rlabel metal2 41832 462 41832 462 0 wbs_dat_o[2]
rlabel metal3 57568 3304 57568 3304 0 wbs_dat_o[30]
rlabel metal4 211288 353 211288 353 0 wbs_dat_o[31]
rlabel metal2 49448 854 49448 854 0 wbs_dat_o[3]
rlabel metal3 40376 3752 40376 3752 0 wbs_dat_o[4]
rlabel metal4 60536 2744 60536 2744 0 wbs_dat_o[5]
rlabel metal3 68376 2744 68376 2744 0 wbs_dat_o[6]
rlabel metal2 74200 1638 74200 1638 0 wbs_dat_o[7]
rlabel metal3 79912 2856 79912 2856 0 wbs_dat_o[8]
rlabel metal2 43400 2058 43400 2058 0 wbs_dat_o[9]
rlabel metal2 28728 574 28728 574 0 wbs_sel_i[0]
rlabel metal2 36344 462 36344 462 0 wbs_sel_i[1]
rlabel metal2 43736 910 43736 910 0 wbs_sel_i[2]
rlabel metal2 51240 280 51240 280 0 wbs_sel_i[3]
rlabel metal2 19320 392 19320 392 0 wbs_stb_i
rlabel metal2 21112 462 21112 462 0 wbs_we_i
<< properties >>
string FIXED_BBOX 0 0 596040 596040
<< end >>
